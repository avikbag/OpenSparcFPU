
module dffrl_async_SIZE1_0 ( din, clk, rst_l, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  wire   N4, n1;

  DFFARX1_RVT \q_reg[0]  ( .D(N4), .CLK(clk), .RSTB(rst_l), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
endmodule


module dffr_SIZE1_0 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dff_SIZE1_0 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE5_0 ( din, clk, se, si, so, \q[4] , \q[3] , \q[2] , \q[1]_BAR , 
        \q[0]_BAR  );
  input [4:0] din;
  input [4:0] si;
  output [4:0] so;
  input clk, se;
  output \q[4] , \q[3] , \q[2] , \q[1]_BAR , \q[0]_BAR ;
  wire   N3, N4, N5, N6, N7, n1;
  wire   [4:0] q;

  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .QN(\q[1]_BAR ) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .QN(\q[0]_BAR ) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_0 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_0 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_6 ( din, rst, en, clk, se, si, so, \q[3]_BAR , \q[2] , 
        \q[1] , \q[0]  );
  input [3:0] din;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  output \q[3]_BAR , \q[2] , \q[1] , \q[0] ;
  wire   N10, N11, N12, N13, net24426, n2, n3, n5, n6;
  wire   [3:0] q;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_6 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .QN(\q[3]_BAR ) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n3) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n5) );
  AND2X1_RVT U4 ( .A1(en), .A2(n5), .Y(n2) );
  AND2X1_RVT U5 ( .A1(n2), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n2), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n2), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n2), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n5), .A2(n3), .Y(n6) );
endmodule


module dff_SIZE4_0 ( din, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, n1;

  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
endmodule


module dff_SIZE4_3 ( din, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, n1;

  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
endmodule


module dff_SIZE4_2 ( din, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, n1;

  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
endmodule


module dff_SIZE1_31 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE4_1 ( din, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, n1;

  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
endmodule


module dffre_SIZE1_0 ( rst, en, clk, q, se, si, so, \din[0]_BAR  );
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se, \din[0]_BAR ;
  wire   \din[0] , n4;
  assign \din[0]  = \din[0]_BAR ;

  DFFX1_RVT \q_reg[0]  ( .D(n4), .CLK(clk), .Q(q[0]) );
  NOR3X0_RVT U2 ( .A1(rst), .A2(se), .A3(\din[0] ), .Y(n4) );
endmodule


module dff_SIZE8_0 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;

  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
endmodule


module dff_SIZE8_5 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;

  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
endmodule


module dff_SIZE16 ( din, clk, q, se, si, so );
  input [15:0] din;
  output [15:0] q;
  input [15:0] si;
  output [15:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, n1;

  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_0 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_0 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_18 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_18 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_17 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_17 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_16 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_16 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_15 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_15 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_14 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_14 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_13 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_13 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_12 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_12 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_11 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_11 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_10 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_10 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_9 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_9 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_8 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_8 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_7 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_7 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_6 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_6 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_5 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_5 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_4 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_4 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffre_SIZE1_14 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffre_SIZE1_13 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffre_SIZE1_12 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffre_SIZE1_11 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module fpu_in_ctl ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, fp_op_in, 
        fp_op_in_7in, a1stg_step, m1stg_step, d1stg_step, add_pipe_active, 
        mul_pipe_active, div_pipe_active, sehold, arst_l, grst_l, rclk, 
        fp_data_rdy, fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_we, 
        inq_wraddr, inq_read_en, inq_rdaddr, inq_bp, inq_bp_inv, inq_fwrd, 
        inq_fwrd_inv, inq_add, inq_mul, inq_div, se, si, so );
  input [123:118] pcx_fpio_data_px2;
  input [3:2] fp_op_in;
  output [3:0] inq_wraddr;
  output [3:0] inq_rdaddr;
  input pcx_fpio_data_rdy_px2, fp_op_in_7in, a1stg_step, m1stg_step,
         d1stg_step, add_pipe_active, mul_pipe_active, div_pipe_active, sehold,
         arst_l, grst_l, rclk, se, si;
  output fp_data_rdy, fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_we,
         inq_read_en, inq_bp, inq_bp_inv, inq_fwrd, inq_fwrd_inv, inq_add,
         inq_mul, inq_div, so;
  wire   in_ctl_rst_l, fp_vld_in, inq_wrptr_step, inq_div_rd, valid_packet,
         valid_packet_dly, fp_add_in, fp_mul_in, inq_pipe0_we, inq_pipe1_we,
         inq_pipe2_we, inq_pipe3_we, inq_pipe4_we, inq_pipe5_we, inq_pipe6_we,
         inq_pipe7_we, inq_pipe8_we, inq_pipe9_we, inq_pipe10_we,
         inq_pipe11_we, inq_pipe12_we, inq_pipe13_we, inq_pipe14_we,
         inq_pipe15_we, d1stg_step_dly, inq_diva_dly, inq_adda_dly,
         inq_mula_dly, n108, n109, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97;
  wire   [4:0] fp_type_in;
  wire   [3:0] inq_wrptr;
  wire   [3:0] inq_wrptr_plus1;
  wire   [3:0] inq_div_wrptr;
  wire   [3:0] inq_div_wrptr_plus1;
  wire   [3:0] inq_wraddr_del;
  wire   [3:0] inq_rdptr;
  wire   [3:0] inq_rdptr_in;
  wire   [3:0] inq_div_rdptr;
  wire   [3:0] inq_div_rdptr_in;
  wire   [3:0] inq_rdaddr_del;
  wire   [7:0] inq_rdptr_dec;
  wire   [7:0] inq_rdptr_dec_in;
  wire   [7:0] inq_div_rdptr_dec;
  wire   [7:0] inq_div_rdptr_dec_in;
  wire   [15:0] inq_rdaddr_del_dec_in;
  wire   [15:0] inq_rdaddr_del_dec;
  wire   [2:0] inq_pipe0;
  wire   [2:0] inq_pipe1;
  wire   [2:0] inq_pipe2;
  wire   [2:0] inq_pipe3;
  wire   [2:0] inq_pipe4;
  wire   [2:0] inq_pipe5;
  wire   [2:0] inq_pipe6;
  wire   [2:0] inq_pipe7;
  wire   [2:0] inq_pipe8;
  wire   [2:0] inq_pipe9;
  wire   [2:0] inq_pipe10;
  wire   [2:0] inq_pipe11;
  wire   [2:0] inq_pipe12;
  wire   [2:0] inq_pipe13;
  wire   [2:0] inq_pipe14;
  wire   [2:0] inq_pipe15;
  assign so = 1'b0;

  dffrl_async_SIZE1_0 dffrl_in_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(in_ctl_rst_l), .se(se), .si(1'b0) );
  dffr_SIZE1_0 i_fp_data_rdy ( .din(pcx_fpio_data_rdy_px2), .clk(rclk), .rst(
        n97), .q(fp_data_rdy), .se(se), .si(1'b0) );
  dff_SIZE1_0 i_fp_vld_in ( .din(pcx_fpio_data_px2[123]), .clk(rclk), .q(
        fp_vld_in), .se(se), .si(1'b0) );
  dff_SIZE5_0 i_fp_type_in ( .din(pcx_fpio_data_px2[122:118]), .clk(rclk), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\q[4] (fp_type_in[4]), 
        .\q[3] (fp_type_in[3]), .\q[2] (fp_type_in[2]), .\q[1]_BAR (
        fp_type_in[1]), .\q[0]_BAR (fp_type_in[0]) );
  dffre_SIZE4_0 i_inq_wrptr ( .din({inq_wrptr_plus1[3:1], n108}), .rst(n97), 
        .en(inq_wrptr_step), .clk(rclk), .q(inq_wrptr), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_6 i_inq_div_wrptr ( .din({inq_div_wrptr_plus1[3:1], n109}), 
        .rst(n97), .en(inq_wraddr[3]), .clk(rclk), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0}), .\q[3]_BAR (inq_div_wrptr[3]), .\q[2] (inq_div_wrptr[2]), 
        .\q[1] (inq_div_wrptr[1]), .\q[0] (inq_div_wrptr[0]) );
  dff_SIZE4_0 i_inq_wraddr_del ( .din(inq_wraddr), .clk(rclk), .q(
        inq_wraddr_del), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE4_3 i_inq_rdptr ( .din(inq_rdptr_in), .clk(rclk), .q(inq_rdptr), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE4_2 i_inq_div_rdptr ( .din(inq_div_rdptr_in), .clk(rclk), .q(
        inq_div_rdptr), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE1_31 i_inq_div_rd ( .din(inq_rdaddr[3]), .clk(rclk), .q(inq_div_rd), 
        .se(se), .si(1'b0) );
  dff_SIZE4_1 i_inq_rdaddr_del ( .din(inq_rdaddr), .clk(rclk), .q(
        inq_rdaddr_del), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_0 i_valid_packet_dly ( .rst(n97), .en(1'b1), .clk(rclk), .q(
        valid_packet_dly), .se(se), .si(1'b0), .\din[0]_BAR (n25) );
  dff_SIZE8_0 i_inq_rdptr_dec ( .din(inq_rdptr_dec_in), .clk(rclk), .q(
        inq_rdptr_dec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dff_SIZE8_5 i_inq_div_rdptr_dec ( .din(inq_div_rdptr_dec_in), .clk(rclk), 
        .q(inq_div_rdptr_dec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE16 i_inq_rdaddr_del_dec ( .din(inq_rdaddr_del_dec_in), .clk(rclk), 
        .q(inq_rdaddr_del_dec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_0 i_inq_pipe0 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe0_we), .clk(rclk), .q(inq_pipe0), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_18 i_inq_pipe1 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe1_we), .clk(rclk), .q(inq_pipe1), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_17 i_inq_pipe2 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe2_we), .clk(rclk), .q(inq_pipe2), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_16 i_inq_pipe3 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe3_we), .clk(rclk), .q(inq_pipe3), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_15 i_inq_pipe4 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe4_we), .clk(rclk), .q(inq_pipe4), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_14 i_inq_pipe5 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe5_we), .clk(rclk), .q(inq_pipe5), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_13 i_inq_pipe6 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe6_we), .clk(rclk), .q(inq_pipe6), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_12 i_inq_pipe7 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe7_we), .clk(rclk), .q(inq_pipe7), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_11 i_inq_pipe8 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe8_we), .clk(rclk), .q(inq_pipe8), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_10 i_inq_pipe9 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe9_we), .clk(rclk), .q(inq_pipe9), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_9 i_inq_pipe10 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe10_we), .clk(rclk), .q(inq_pipe10), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_8 i_inq_pipe11 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe11_we), .clk(rclk), .q(inq_pipe11), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_7 i_inq_pipe12 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe12_we), .clk(rclk), .q(inq_pipe12), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_6 i_inq_pipe13 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe13_we), .clk(rclk), .q(inq_pipe13), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_5 i_inq_pipe14 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe14_we), .clk(rclk), .q(inq_pipe14), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_4 i_inq_pipe15 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(n97), .en(inq_pipe15_we), .clk(rclk), .q(inq_pipe15), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_14 i_inq_adda_dly ( .din(inq_add), .rst(n97), .en(1'b1), .clk(
        rclk), .q(inq_adda_dly), .se(se), .si(1'b0) );
  dffre_SIZE1_13 i_inq_mula_dly ( .din(inq_mul), .rst(n97), .en(1'b1), .clk(
        rclk), .q(inq_mula_dly), .se(se), .si(1'b0) );
  dffre_SIZE1_12 i_inq_diva_dly ( .din(inq_div), .rst(n97), .en(1'b1), .clk(
        rclk), .q(inq_diva_dly), .se(se), .si(1'b0) );
  dffre_SIZE1_11 i_d1stg_step_dly ( .din(d1stg_step), .rst(n97), .en(1'b1), 
        .clk(rclk), .q(d1stg_step_dly), .se(se), .si(1'b0) );
  INVX0_RVT U2 ( .A(n67), .Y(n69) );
  INVX0_RVT U3 ( .A(n70), .Y(n72) );
  INVX0_RVT U4 ( .A(n62), .Y(n66) );
  INVX0_RVT U5 ( .A(n73), .Y(n40) );
  INVX0_RVT U6 ( .A(n46), .Y(n41) );
  INVX0_RVT U7 ( .A(inq_div), .Y(n24) );
  INVX0_RVT U8 ( .A(n23), .Y(n65) );
  INVX0_RVT U9 ( .A(inq_div_rdptr[3]), .Y(n71) );
  INVX0_RVT U10 ( .A(fp_op_in[3]), .Y(n26) );
  INVX0_RVT U11 ( .A(fp_op_in[2]), .Y(n3) );
  INVX1_RVT U12 ( .A(fp_data_rdy), .Y(n1) );
  NOR4X1_RVT U13 ( .A1(fp_type_in[2]), .A2(fp_type_in[1]), .A3(fp_type_in[4]), 
        .A4(n1), .Y(n2) );
  NAND3X0_RVT U14 ( .A1(fp_vld_in), .A2(fp_type_in[3]), .A3(n2), .Y(n25) );
  NOR3X0_RVT U15 ( .A1(fp_type_in[0]), .A2(fp_op_in_7in), .A3(n25), .Y(n28) );
  NAND3X0_RVT U16 ( .A1(fp_op_in[3]), .A2(n28), .A3(fp_op_in[2]), .Y(n63) );
  INVX1_RVT U17 ( .A(n63), .Y(inq_wraddr[3]) );
  AND3X1_RVT U18 ( .A1(n28), .A2(fp_op_in[3]), .A3(n3), .Y(fp_mul_in) );
  INVX1_RVT U19 ( .A(inq_div_wrptr[0]), .Y(n109) );
  INVX1_RVT U20 ( .A(inq_div_rdptr[0]), .Y(n74) );
  INVX1_RVT U21 ( .A(inq_div_wrptr[2]), .Y(n85) );
  INVX1_RVT U22 ( .A(inq_div_rdptr[2]), .Y(n42) );
  INVX1_RVT U23 ( .A(inq_div_wrptr[1]), .Y(n86) );
  AOI22X1_RVT U24 ( .A1(n86), .A2(inq_div_rdptr[1]), .A3(inq_div_wrptr[3]), 
        .A4(inq_div_rdptr[3]), .Y(n4) );
  OA221X1_RVT U25 ( .A1(n86), .A2(inq_div_rdptr[1]), .A3(inq_div_wrptr[3]), 
        .A4(inq_div_rdptr[3]), .A5(n4), .Y(n5) );
  OA221X1_RVT U26 ( .A1(inq_div_rdptr[2]), .A2(n85), .A3(n42), .A4(
        inq_div_wrptr[2]), .A5(n5), .Y(n6) );
  OA221X1_RVT U27 ( .A1(inq_div_rdptr[0]), .A2(n109), .A3(n74), .A4(
        inq_div_wrptr[0]), .A5(n6), .Y(n23) );
  NAND3X0_RVT U28 ( .A1(n23), .A2(d1stg_step), .A3(inq_wraddr[3]), .Y(n10) );
  NOR2X0_RVT U29 ( .A1(inq_diva_dly), .A2(n10), .Y(n22) );
  INVX1_RVT U30 ( .A(inq_rdptr[2]), .Y(n60) );
  INVX1_RVT U31 ( .A(inq_wrptr[2]), .Y(n84) );
  INVX1_RVT U32 ( .A(inq_wrptr[0]), .Y(n108) );
  INVX1_RVT U33 ( .A(inq_rdptr[0]), .Y(n75) );
  INVX1_RVT U34 ( .A(inq_rdptr[3]), .Y(n68) );
  INVX1_RVT U35 ( .A(inq_wrptr[1]), .Y(n88) );
  OAI22X1_RVT U36 ( .A1(inq_wrptr[3]), .A2(n68), .A3(n88), .A4(inq_rdptr[1]), 
        .Y(n7) );
  AO221X1_RVT U37 ( .A1(n68), .A2(inq_wrptr[3]), .A3(n88), .A4(inq_rdptr[1]), 
        .A5(n7), .Y(n8) );
  AO221X1_RVT U38 ( .A1(inq_rdptr[0]), .A2(n108), .A3(n75), .A4(inq_wrptr[0]), 
        .A5(n8), .Y(n9) );
  AO221X1_RVT U39 ( .A1(inq_wrptr[2]), .A2(n60), .A3(n84), .A4(inq_rdptr[2]), 
        .A5(n9), .Y(n64) );
  OA21X1_RVT U40 ( .A1(inq_div_rd), .A2(n64), .A3(n10), .Y(n59) );
  AO22X1_RVT U41 ( .A1(inq_rdaddr_del_dec[1]), .A2(inq_pipe1[2]), .A3(
        inq_rdaddr_del_dec[0]), .A4(inq_pipe0[2]), .Y(n14) );
  AO22X1_RVT U42 ( .A1(inq_rdaddr_del_dec[3]), .A2(inq_pipe3[2]), .A3(
        inq_rdaddr_del_dec[2]), .A4(inq_pipe2[2]), .Y(n13) );
  AO22X1_RVT U43 ( .A1(inq_rdaddr_del_dec[5]), .A2(inq_pipe5[2]), .A3(
        inq_rdaddr_del_dec[4]), .A4(inq_pipe4[2]), .Y(n12) );
  AO22X1_RVT U44 ( .A1(inq_rdaddr_del_dec[7]), .A2(inq_pipe7[2]), .A3(
        inq_rdaddr_del_dec[6]), .A4(inq_pipe6[2]), .Y(n11) );
  NOR4X1_RVT U45 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .Y(n20) );
  AO22X1_RVT U46 ( .A1(inq_rdaddr_del_dec[9]), .A2(inq_pipe9[2]), .A3(
        inq_rdaddr_del_dec[8]), .A4(inq_pipe8[2]), .Y(n18) );
  AO22X1_RVT U47 ( .A1(inq_rdaddr_del_dec[11]), .A2(inq_pipe11[2]), .A3(
        inq_rdaddr_del_dec[10]), .A4(inq_pipe10[2]), .Y(n17) );
  AO22X1_RVT U48 ( .A1(inq_rdaddr_del_dec[13]), .A2(inq_pipe13[2]), .A3(
        inq_rdaddr_del_dec[12]), .A4(inq_pipe12[2]), .Y(n16) );
  AO22X1_RVT U49 ( .A1(inq_rdaddr_del_dec[15]), .A2(inq_pipe15[2]), .A3(
        inq_rdaddr_del_dec[14]), .A4(inq_pipe14[2]), .Y(n15) );
  NOR4X1_RVT U50 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .Y(n19) );
  NAND2X0_RVT U51 ( .A1(n20), .A2(n19), .Y(n21) );
  AO22X1_RVT U52 ( .A1(d1stg_step_dly), .A2(n22), .A3(n59), .A4(n21), .Y(
        inq_div) );
  NAND3X0_RVT U53 ( .A1(d1stg_step), .A2(n24), .A3(n65), .Y(n83) );
  INVX1_RVT U54 ( .A(n83), .Y(inq_rdaddr[3]) );
  INVX1_RVT U55 ( .A(n25), .Y(valid_packet) );
  AND3X1_RVT U56 ( .A1(valid_packet), .A2(fp_type_in[0]), .A3(fp_op_in_7in), 
        .Y(n27) );
  AO21X1_RVT U57 ( .A1(n28), .A2(n26), .A3(n27), .Y(fp_add_in) );
  OR2X1_RVT U58 ( .A1(n28), .A2(n27), .Y(inq_we) );
  AND2X1_RVT U59 ( .A1(n63), .A2(inq_we), .Y(inq_wrptr_step) );
  INVX1_RVT U60 ( .A(in_ctl_rst_l), .Y(n97) );
  AO22X1_RVT U61 ( .A1(inq_rdaddr_del_dec[11]), .A2(inq_pipe11[0]), .A3(
        inq_rdaddr_del_dec[10]), .A4(inq_pipe10[0]), .Y(n32) );
  AO22X1_RVT U62 ( .A1(inq_rdaddr_del_dec[9]), .A2(inq_pipe9[0]), .A3(
        inq_rdaddr_del_dec[8]), .A4(inq_pipe8[0]), .Y(n31) );
  AO22X1_RVT U63 ( .A1(inq_rdaddr_del_dec[15]), .A2(inq_pipe15[0]), .A3(
        inq_rdaddr_del_dec[14]), .A4(inq_pipe14[0]), .Y(n30) );
  AO22X1_RVT U64 ( .A1(inq_rdaddr_del_dec[13]), .A2(inq_pipe13[0]), .A3(
        inq_rdaddr_del_dec[12]), .A4(inq_pipe12[0]), .Y(n29) );
  NOR4X1_RVT U65 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .Y(n38) );
  AO22X1_RVT U66 ( .A1(inq_rdaddr_del_dec[1]), .A2(inq_pipe1[0]), .A3(
        inq_rdaddr_del_dec[0]), .A4(inq_pipe0[0]), .Y(n36) );
  AO22X1_RVT U67 ( .A1(inq_rdaddr_del_dec[3]), .A2(inq_pipe3[0]), .A3(
        inq_rdaddr_del_dec[2]), .A4(inq_pipe2[0]), .Y(n35) );
  AO22X1_RVT U68 ( .A1(inq_rdaddr_del_dec[5]), .A2(inq_pipe5[0]), .A3(
        inq_rdaddr_del_dec[4]), .A4(inq_pipe4[0]), .Y(n34) );
  AO22X1_RVT U69 ( .A1(inq_rdaddr_del_dec[7]), .A2(inq_pipe7[0]), .A3(
        inq_rdaddr_del_dec[6]), .A4(inq_pipe6[0]), .Y(n33) );
  NOR4X1_RVT U70 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .Y(n37) );
  NAND2X0_RVT U71 ( .A1(n38), .A2(n37), .Y(n39) );
  INVX1_RVT U72 ( .A(n59), .Y(n57) );
  AO22X1_RVT U73 ( .A1(n59), .A2(n39), .A3(n57), .A4(fp_add_in), .Y(inq_add)
         );
  NAND2X0_RVT U74 ( .A1(d1stg_step), .A2(inq_div), .Y(n73) );
  AO221X1_RVT U75 ( .A1(n40), .A2(inq_div_rdptr_dec[7]), .A3(n73), .A4(
        inq_div_rdptr_dec[0]), .A5(n97), .Y(inq_div_rdptr_dec_in[0]) );
  NAND4X0_RVT U76 ( .A1(inq_div_rdptr[0]), .A2(inq_div_rdptr[1]), .A3(
        d1stg_step), .A4(inq_div), .Y(n46) );
  NAND2X0_RVT U77 ( .A1(inq_div_rdptr[2]), .A2(n41), .Y(n70) );
  AND2X1_RVT U78 ( .A1(n70), .A2(in_ctl_rst_l), .Y(n44) );
  NAND2X0_RVT U79 ( .A1(n42), .A2(n46), .Y(n43) );
  AND2X1_RVT U80 ( .A1(n44), .A2(n43), .Y(inq_div_rdptr_in[2]) );
  INVX1_RVT U81 ( .A(sehold), .Y(n95) );
  NAND3X0_RVT U82 ( .A1(valid_packet), .A2(n57), .A3(n95), .Y(inq_fwrd_inv) );
  AND3X1_RVT U84 ( .A1(d1stg_step), .A2(in_ctl_rst_l), .A3(inq_div), .Y(n77)
         );
  AO22X1_RVT U85 ( .A1(in_ctl_rst_l), .A2(inq_div_rdptr[1]), .A3(
        inq_div_rdptr[0]), .A4(n77), .Y(n45) );
  AND2X1_RVT U86 ( .A1(n46), .A2(n45), .Y(inq_div_rdptr_in[1]) );
  AO22X1_RVT U87 ( .A1(inq_rdaddr_del_dec[11]), .A2(inq_pipe11[1]), .A3(
        inq_rdaddr_del_dec[10]), .A4(inq_pipe10[1]), .Y(n50) );
  AO22X1_RVT U88 ( .A1(inq_rdaddr_del_dec[9]), .A2(inq_pipe9[1]), .A3(
        inq_rdaddr_del_dec[8]), .A4(inq_pipe8[1]), .Y(n49) );
  AO22X1_RVT U89 ( .A1(inq_rdaddr_del_dec[15]), .A2(inq_pipe15[1]), .A3(
        inq_rdaddr_del_dec[14]), .A4(inq_pipe14[1]), .Y(n48) );
  AO22X1_RVT U90 ( .A1(inq_rdaddr_del_dec[13]), .A2(inq_pipe13[1]), .A3(
        inq_rdaddr_del_dec[12]), .A4(inq_pipe12[1]), .Y(n47) );
  NOR4X1_RVT U91 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .Y(n56) );
  AO22X1_RVT U92 ( .A1(inq_rdaddr_del_dec[1]), .A2(inq_pipe1[1]), .A3(
        inq_rdaddr_del_dec[0]), .A4(inq_pipe0[1]), .Y(n54) );
  AO22X1_RVT U93 ( .A1(inq_rdaddr_del_dec[3]), .A2(inq_pipe3[1]), .A3(
        inq_rdaddr_del_dec[2]), .A4(inq_pipe2[1]), .Y(n53) );
  AO22X1_RVT U94 ( .A1(inq_rdaddr_del_dec[5]), .A2(inq_pipe5[1]), .A3(
        inq_rdaddr_del_dec[4]), .A4(inq_pipe4[1]), .Y(n52) );
  AO22X1_RVT U95 ( .A1(inq_rdaddr_del_dec[7]), .A2(inq_pipe7[1]), .A3(
        inq_rdaddr_del_dec[6]), .A4(inq_pipe6[1]), .Y(n51) );
  NOR4X1_RVT U96 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .Y(n55) );
  NAND2X0_RVT U97 ( .A1(n56), .A2(n55), .Y(n58) );
  AO22X1_RVT U98 ( .A1(n59), .A2(n58), .A3(n57), .A4(fp_mul_in), .Y(inq_mul)
         );
  AO22X1_RVT U99 ( .A1(inq_add), .A2(a1stg_step), .A3(inq_mul), .A4(m1stg_step), .Y(n81) );
  NAND3X0_RVT U100 ( .A1(inq_rdptr[0]), .A2(inq_rdptr[1]), .A3(n81), .Y(n62)
         );
  OA221X1_RVT U101 ( .A1(inq_rdptr[2]), .A2(n66), .A3(n60), .A4(n62), .A5(
        in_ctl_rst_l), .Y(inq_rdptr_in[2]) );
  AND2X1_RVT U102 ( .A1(in_ctl_rst_l), .A2(n81), .Y(n80) );
  AO22X1_RVT U103 ( .A1(in_ctl_rst_l), .A2(inq_rdptr[1]), .A3(inq_rdptr[0]), 
        .A4(n80), .Y(n61) );
  AND2X1_RVT U104 ( .A1(n62), .A2(n61), .Y(inq_rdptr_in[1]) );
  AO22X1_RVT U105 ( .A1(inq_wraddr[3]), .A2(inq_div_wrptr[2]), .A3(n63), .A4(
        inq_wrptr[2]), .Y(inq_wraddr[2]) );
  AO22X1_RVT U106 ( .A1(inq_wraddr[3]), .A2(inq_div_wrptr[1]), .A3(n63), .A4(
        inq_wrptr[1]), .Y(inq_wraddr[1]) );
  AO22X1_RVT U107 ( .A1(inq_wraddr[3]), .A2(inq_div_wrptr[0]), .A3(n63), .A4(
        inq_wrptr[0]), .Y(inq_wraddr[0]) );
  OR2X1_RVT U108 ( .A1(n65), .A2(n64), .Y(inq_read_en) );
  NAND2X0_RVT U109 ( .A1(inq_rdptr[2]), .A2(n66), .Y(n67) );
  OA221X1_RVT U110 ( .A1(inq_rdptr[3]), .A2(n69), .A3(n68), .A4(n67), .A5(
        in_ctl_rst_l), .Y(inq_rdptr_in[3]) );
  OA221X1_RVT U111 ( .A1(inq_div_rdptr[3]), .A2(n72), .A3(n71), .A4(n70), .A5(
        in_ctl_rst_l), .Y(inq_div_rdptr_in[3]) );
  AND2X1_RVT U112 ( .A1(in_ctl_rst_l), .A2(n73), .Y(n76) );
  AO22X1_RVT U113 ( .A1(inq_div_rdptr[0]), .A2(n76), .A3(n74), .A4(n77), .Y(
        inq_div_rdptr_in[0]) );
  AND2X1_RVT U114 ( .A1(in_ctl_rst_l), .A2(inq_rdaddr[3]), .Y(n78) );
  AO22X1_RVT U115 ( .A1(inq_div_rdptr[2]), .A2(n78), .A3(inq_rdptr_in[2]), 
        .A4(n83), .Y(inq_rdaddr[2]) );
  AO22X1_RVT U116 ( .A1(inq_div_rdptr[1]), .A2(n78), .A3(inq_rdptr_in[1]), 
        .A4(n83), .Y(inq_rdaddr[1]) );
  INVX1_RVT U117 ( .A(n81), .Y(n82) );
  AND2X1_RVT U118 ( .A1(in_ctl_rst_l), .A2(n82), .Y(n79) );
  AO22X1_RVT U119 ( .A1(inq_rdptr[0]), .A2(n79), .A3(n75), .A4(n80), .Y(
        inq_rdptr_in[0]) );
  AO22X1_RVT U120 ( .A1(inq_div_rdptr[0]), .A2(n78), .A3(n83), .A4(
        inq_rdptr_in[0]), .Y(inq_rdaddr[0]) );
  AO22X1_RVT U121 ( .A1(n77), .A2(inq_div_rdptr_dec[6]), .A3(n76), .A4(
        inq_div_rdptr_dec[7]), .Y(inq_div_rdptr_dec_in[7]) );
  AO22X1_RVT U122 ( .A1(n77), .A2(inq_div_rdptr_dec[5]), .A3(n76), .A4(
        inq_div_rdptr_dec[6]), .Y(inq_div_rdptr_dec_in[6]) );
  AO22X1_RVT U123 ( .A1(n77), .A2(inq_div_rdptr_dec[4]), .A3(n76), .A4(
        inq_div_rdptr_dec[5]), .Y(inq_div_rdptr_dec_in[5]) );
  AO22X1_RVT U124 ( .A1(n77), .A2(inq_div_rdptr_dec[3]), .A3(n76), .A4(
        inq_div_rdptr_dec[4]), .Y(inq_div_rdptr_dec_in[4]) );
  AO22X1_RVT U125 ( .A1(n77), .A2(inq_div_rdptr_dec[2]), .A3(n76), .A4(
        inq_div_rdptr_dec[3]), .Y(inq_div_rdptr_dec_in[3]) );
  AO22X1_RVT U126 ( .A1(n77), .A2(inq_div_rdptr_dec[1]), .A3(n76), .A4(
        inq_div_rdptr_dec[2]), .Y(inq_div_rdptr_dec_in[2]) );
  AO22X1_RVT U127 ( .A1(n77), .A2(inq_div_rdptr_dec[0]), .A3(n76), .A4(
        inq_div_rdptr_dec[1]), .Y(inq_div_rdptr_dec_in[1]) );
  AND2X1_RVT U128 ( .A1(n78), .A2(inq_div_rdptr_dec[7]), .Y(
        inq_rdaddr_del_dec_in[15]) );
  AND2X1_RVT U129 ( .A1(n78), .A2(inq_div_rdptr_dec[6]), .Y(
        inq_rdaddr_del_dec_in[14]) );
  AND2X1_RVT U130 ( .A1(n78), .A2(inq_div_rdptr_dec[5]), .Y(
        inq_rdaddr_del_dec_in[13]) );
  AND2X1_RVT U131 ( .A1(n78), .A2(inq_div_rdptr_dec[4]), .Y(
        inq_rdaddr_del_dec_in[12]) );
  AND2X1_RVT U132 ( .A1(n78), .A2(inq_div_rdptr_dec[3]), .Y(
        inq_rdaddr_del_dec_in[11]) );
  AND2X1_RVT U133 ( .A1(n78), .A2(inq_div_rdptr_dec[2]), .Y(
        inq_rdaddr_del_dec_in[10]) );
  AND2X1_RVT U134 ( .A1(n78), .A2(inq_div_rdptr_dec[1]), .Y(
        inq_rdaddr_del_dec_in[9]) );
  OA21X1_RVT U135 ( .A1(inq_div_rdptr_dec[0]), .A2(n97), .A3(inq_rdaddr[3]), 
        .Y(inq_rdaddr_del_dec_in[8]) );
  AO22X1_RVT U136 ( .A1(n80), .A2(inq_rdptr_dec[6]), .A3(n79), .A4(
        inq_rdptr_dec[7]), .Y(inq_rdptr_dec_in[7]) );
  AND2X1_RVT U137 ( .A1(n83), .A2(inq_rdptr_dec_in[7]), .Y(
        inq_rdaddr_del_dec_in[7]) );
  AO22X1_RVT U138 ( .A1(n80), .A2(inq_rdptr_dec[5]), .A3(n79), .A4(
        inq_rdptr_dec[6]), .Y(inq_rdptr_dec_in[6]) );
  AND2X1_RVT U139 ( .A1(n83), .A2(inq_rdptr_dec_in[6]), .Y(
        inq_rdaddr_del_dec_in[6]) );
  AO22X1_RVT U140 ( .A1(n80), .A2(inq_rdptr_dec[4]), .A3(n79), .A4(
        inq_rdptr_dec[5]), .Y(inq_rdptr_dec_in[5]) );
  AND2X1_RVT U141 ( .A1(n83), .A2(inq_rdptr_dec_in[5]), .Y(
        inq_rdaddr_del_dec_in[5]) );
  AO22X1_RVT U142 ( .A1(n80), .A2(inq_rdptr_dec[3]), .A3(n79), .A4(
        inq_rdptr_dec[4]), .Y(inq_rdptr_dec_in[4]) );
  AND2X1_RVT U143 ( .A1(n83), .A2(inq_rdptr_dec_in[4]), .Y(
        inq_rdaddr_del_dec_in[4]) );
  AO22X1_RVT U144 ( .A1(n80), .A2(inq_rdptr_dec[2]), .A3(n79), .A4(
        inq_rdptr_dec[3]), .Y(inq_rdptr_dec_in[3]) );
  AND2X1_RVT U145 ( .A1(n83), .A2(inq_rdptr_dec_in[3]), .Y(
        inq_rdaddr_del_dec_in[3]) );
  AO22X1_RVT U146 ( .A1(n80), .A2(inq_rdptr_dec[1]), .A3(n79), .A4(
        inq_rdptr_dec[2]), .Y(inq_rdptr_dec_in[2]) );
  AND2X1_RVT U147 ( .A1(n83), .A2(inq_rdptr_dec_in[2]), .Y(
        inq_rdaddr_del_dec_in[2]) );
  AO22X1_RVT U148 ( .A1(n80), .A2(inq_rdptr_dec[0]), .A3(n79), .A4(
        inq_rdptr_dec[1]), .Y(inq_rdptr_dec_in[1]) );
  AND2X1_RVT U149 ( .A1(n83), .A2(inq_rdptr_dec_in[1]), .Y(
        inq_rdaddr_del_dec_in[1]) );
  AO221X1_RVT U150 ( .A1(n82), .A2(inq_rdptr_dec[0]), .A3(n81), .A4(
        inq_rdptr_dec[7]), .A5(n97), .Y(inq_rdptr_dec_in[0]) );
  AND2X1_RVT U151 ( .A1(n83), .A2(inq_rdptr_dec_in[0]), .Y(
        inq_rdaddr_del_dec_in[0]) );
  AND4X1_RVT U152 ( .A1(inq_wrptr_step), .A2(n84), .A3(n88), .A4(n108), .Y(
        inq_pipe0_we) );
  AND4X1_RVT U153 ( .A1(inq_wrptr[0]), .A2(inq_wrptr_step), .A3(n84), .A4(n88), 
        .Y(inq_pipe1_we) );
  AND4X1_RVT U154 ( .A1(inq_wrptr[1]), .A2(inq_wrptr_step), .A3(n84), .A4(n108), .Y(inq_pipe2_we) );
  AND4X1_RVT U155 ( .A1(inq_wrptr[1]), .A2(inq_wrptr[0]), .A3(inq_wrptr_step), 
        .A4(n84), .Y(inq_pipe3_we) );
  AND4X1_RVT U156 ( .A1(inq_wrptr[2]), .A2(inq_wrptr_step), .A3(n108), .A4(n88), .Y(inq_pipe4_we) );
  AND4X1_RVT U157 ( .A1(inq_wrptr[2]), .A2(inq_wrptr[0]), .A3(inq_wrptr_step), 
        .A4(n88), .Y(inq_pipe5_we) );
  AND4X1_RVT U158 ( .A1(inq_wrptr[1]), .A2(inq_wrptr[2]), .A3(inq_wrptr_step), 
        .A4(n108), .Y(inq_pipe6_we) );
  AND4X1_RVT U159 ( .A1(inq_wrptr[2]), .A2(inq_wrptr[1]), .A3(inq_wrptr[0]), 
        .A4(inq_wrptr_step), .Y(inq_pipe7_we) );
  AND4X1_RVT U160 ( .A1(inq_wraddr[3]), .A2(n86), .A3(n109), .A4(n85), .Y(
        inq_pipe8_we) );
  AND4X1_RVT U161 ( .A1(inq_div_wrptr[0]), .A2(inq_wraddr[3]), .A3(n86), .A4(
        n85), .Y(inq_pipe9_we) );
  AND4X1_RVT U162 ( .A1(inq_div_wrptr[1]), .A2(inq_wraddr[3]), .A3(n85), .A4(
        n109), .Y(inq_pipe10_we) );
  AND4X1_RVT U163 ( .A1(inq_div_wrptr[0]), .A2(inq_div_wrptr[1]), .A3(
        inq_wraddr[3]), .A4(n85), .Y(inq_pipe11_we) );
  AND4X1_RVT U164 ( .A1(inq_div_wrptr[2]), .A2(inq_wraddr[3]), .A3(n86), .A4(
        n109), .Y(inq_pipe12_we) );
  AND4X1_RVT U165 ( .A1(inq_div_wrptr[0]), .A2(inq_div_wrptr[2]), .A3(
        inq_wraddr[3]), .A4(n86), .Y(inq_pipe13_we) );
  AND4X1_RVT U166 ( .A1(inq_div_wrptr[1]), .A2(inq_div_wrptr[2]), .A3(
        inq_wraddr[3]), .A4(n109), .Y(inq_pipe14_we) );
  AND4X1_RVT U167 ( .A1(inq_div_wrptr[1]), .A2(inq_div_wrptr[0]), .A3(
        inq_div_wrptr[2]), .A4(inq_wraddr[3]), .Y(inq_pipe15_we) );
  AO22X1_RVT U168 ( .A1(inq_div_wrptr[1]), .A2(n109), .A3(n86), .A4(
        inq_div_wrptr[0]), .Y(inq_div_wrptr_plus1[1]) );
  NAND3X0_RVT U169 ( .A1(inq_div_wrptr[1]), .A2(inq_div_wrptr[0]), .A3(
        inq_div_wrptr[2]), .Y(n87) );
  OA221X1_RVT U170 ( .A1(inq_div_wrptr[2]), .A2(inq_div_wrptr[0]), .A3(
        inq_div_wrptr[2]), .A4(inq_div_wrptr[1]), .A5(n87), .Y(
        inq_div_wrptr_plus1[2]) );
  HADDX1_RVT U171 ( .A0(inq_div_wrptr[3]), .B0(n87), .SO(
        inq_div_wrptr_plus1[3]) );
  AO22X1_RVT U172 ( .A1(inq_wrptr[1]), .A2(n108), .A3(n88), .A4(inq_wrptr[0]), 
        .Y(inq_wrptr_plus1[1]) );
  NAND3X0_RVT U173 ( .A1(inq_wrptr[2]), .A2(inq_wrptr[1]), .A3(inq_wrptr[0]), 
        .Y(n89) );
  OA221X1_RVT U174 ( .A1(inq_wrptr[2]), .A2(inq_wrptr[1]), .A3(inq_wrptr[2]), 
        .A4(inq_wrptr[0]), .A5(n89), .Y(inq_wrptr_plus1[2]) );
  INVX1_RVT U175 ( .A(n89), .Y(n90) );
  HADDX1_RVT U176 ( .A0(inq_wrptr[3]), .B0(n90), .SO(inq_wrptr_plus1[3]) );
  HADDX1_RVT U177 ( .A0(inq_wraddr_del[2]), .B0(inq_rdaddr_del[2]), .SO(n93)
         );
  HADDX1_RVT U178 ( .A0(inq_rdaddr_del[1]), .B0(inq_wraddr_del[1]), .SO(n92)
         );
  HADDX1_RVT U179 ( .A0(inq_wraddr_del[0]), .B0(inq_rdaddr_del[0]), .SO(n91)
         );
  NOR3X0_RVT U180 ( .A1(n93), .A2(n92), .A3(n91), .Y(n96) );
  XNOR2X1_RVT U181 ( .A1(inq_wraddr_del[3]), .A2(inq_rdaddr_del[3]), .Y(n94)
         );
  NAND4X0_RVT U182 ( .A1(valid_packet_dly), .A2(n96), .A3(n95), .A4(n94), .Y(
        inq_bp_inv) );
  NOR4X1_RVT U184 ( .A1(inq_diva_dly), .A2(div_pipe_active), .A3(n97), .A4(
        inq_div), .Y(fdiv_clken_l) );
  NOR4X1_RVT U185 ( .A1(mul_pipe_active), .A2(inq_mul), .A3(inq_mula_dly), 
        .A4(n97), .Y(fmul_clken_l) );
  NOR4X1_RVT U186 ( .A1(add_pipe_active), .A2(inq_add), .A3(inq_adda_dly), 
        .A4(n97), .Y(fadd_clken_l) );
endmodule


module clken_buf_0 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   rclk;
  assign clk = rclk;

endmodule


module dff_SIZE5_2 ( din, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, n1;

  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
endmodule


module dff_SIZE8_4 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;

  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
endmodule


module dff_SIZE2_0 ( din, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input clk, se;
  wire   N3, N4, n1;

  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
endmodule


module dff_SIZE2_2 ( din, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input clk, se;
  wire   N3, N4, n1;

  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
endmodule


module dff_SIZE64_0 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n3), .Y(N57) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n4), .Y(N58) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n2), .Y(N60) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n3), .Y(N61) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n4), .Y(N62) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n2), .Y(N64) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n3), .Y(N65) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n4), .Y(N66) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE69 ( din, en, clk, q, se, si, so );
  input [68:0] din;
  output [68:0] q;
  input [68:0] si;
  output [68:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, net24683,
         n3, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE69 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24683), .TE(1'b0) );
  DFFX1_RVT \q_reg[68]  ( .D(N72), .CLK(net24683), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N71), .CLK(net24683), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N70), .CLK(net24683), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N69), .CLK(net24683), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N68), .CLK(net24683), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24683), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24683), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24683), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24683), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24683), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24683), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24683), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24683), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24683), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24683), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24683), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24683), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24683), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24683), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24683), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24683), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24683), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24683), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24683), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24683), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24683), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24683), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24683), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24683), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24683), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24683), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24683), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24683), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24683), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24683), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24683), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24683), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24683), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24683), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24683), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24683), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24683), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24683), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24683), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24683), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24683), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24683), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24683), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24683), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24683), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24683), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24683), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24683), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24683), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24683), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24683), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24683), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24683), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24683), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24683), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24683), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24683), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24683), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24683), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24683), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24683), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24683), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24683), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24683), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n6) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n6), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n6), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n6), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n6), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n6), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n6), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n6), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n6), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n6), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n6), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n6), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n6), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n1), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n2), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n4), .Y(N66) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n5), .Y(N67) );
  AND2X1_RVT U71 ( .A1(din[64]), .A2(n6), .Y(N68) );
  AND2X1_RVT U72 ( .A1(din[65]), .A2(n1), .Y(N69) );
  AND2X1_RVT U73 ( .A1(din[66]), .A2(n2), .Y(N70) );
  AND2X1_RVT U74 ( .A1(din[67]), .A2(n4), .Y(N71) );
  AND2X1_RVT U75 ( .A1(din[68]), .A2(n5), .Y(N72) );
  OR2X1_RVT U77 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module dff_SIZE155 ( din, clk, q, se, si, so );
  input [154:0] din;
  output [154:0] q;
  input [154:0] si;
  output [154:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, n1;

  DFFX1_RVT \q_reg[154]  ( .D(N157), .CLK(clk), .Q(q[154]) );
  DFFX1_RVT \q_reg[153]  ( .D(N156), .CLK(clk), .Q(q[153]) );
  DFFX1_RVT \q_reg[152]  ( .D(N155), .CLK(clk), .Q(q[152]) );
  DFFX1_RVT \q_reg[151]  ( .D(N154), .CLK(clk), .Q(q[151]) );
  DFFX1_RVT \q_reg[150]  ( .D(N153), .CLK(clk), .Q(q[150]) );
  DFFX1_RVT \q_reg[149]  ( .D(N152), .CLK(clk), .Q(q[149]) );
  DFFX1_RVT \q_reg[148]  ( .D(N151), .CLK(clk), .Q(q[148]) );
  DFFX1_RVT \q_reg[147]  ( .D(N150), .CLK(clk), .Q(q[147]) );
  DFFX1_RVT \q_reg[146]  ( .D(N149), .CLK(clk), .Q(q[146]) );
  DFFX1_RVT \q_reg[145]  ( .D(N148), .CLK(clk), .Q(q[145]) );
  DFFX1_RVT \q_reg[144]  ( .D(N147), .CLK(clk), .Q(q[144]) );
  DFFX1_RVT \q_reg[143]  ( .D(N146), .CLK(clk), .Q(q[143]) );
  DFFX1_RVT \q_reg[142]  ( .D(N145), .CLK(clk), .Q(q[142]) );
  DFFX1_RVT \q_reg[141]  ( .D(N144), .CLK(clk), .Q(q[141]) );
  DFFX1_RVT \q_reg[140]  ( .D(N143), .CLK(clk), .Q(q[140]) );
  DFFX1_RVT \q_reg[139]  ( .D(N142), .CLK(clk), .Q(q[139]) );
  DFFX1_RVT \q_reg[138]  ( .D(N141), .CLK(clk), .Q(q[138]) );
  DFFX1_RVT \q_reg[137]  ( .D(N140), .CLK(clk), .Q(q[137]) );
  DFFX1_RVT \q_reg[136]  ( .D(N139), .CLK(clk), .Q(q[136]) );
  DFFX1_RVT \q_reg[135]  ( .D(N138), .CLK(clk), .Q(q[135]) );
  DFFX1_RVT \q_reg[134]  ( .D(N137), .CLK(clk), .Q(q[134]) );
  DFFX1_RVT \q_reg[133]  ( .D(N136), .CLK(clk), .Q(q[133]) );
  DFFX1_RVT \q_reg[132]  ( .D(N135), .CLK(clk), .Q(q[132]) );
  DFFX1_RVT \q_reg[131]  ( .D(N134), .CLK(clk), .Q(q[131]) );
  DFFX1_RVT \q_reg[130]  ( .D(N133), .CLK(clk), .Q(q[130]) );
  DFFX1_RVT \q_reg[129]  ( .D(N132), .CLK(clk), .Q(q[129]) );
  DFFX1_RVT \q_reg[128]  ( .D(N131), .CLK(clk), .Q(q[128]) );
  DFFX1_RVT \q_reg[127]  ( .D(N130), .CLK(clk), .Q(q[127]) );
  DFFX1_RVT \q_reg[126]  ( .D(N129), .CLK(clk), .Q(q[126]) );
  DFFX1_RVT \q_reg[125]  ( .D(N128), .CLK(clk), .Q(q[125]) );
  DFFX1_RVT \q_reg[124]  ( .D(N127), .CLK(clk), .Q(q[124]) );
  DFFX1_RVT \q_reg[123]  ( .D(N126), .CLK(clk), .Q(q[123]) );
  DFFX1_RVT \q_reg[122]  ( .D(N125), .CLK(clk), .Q(q[122]) );
  DFFX1_RVT \q_reg[121]  ( .D(N124), .CLK(clk), .Q(q[121]) );
  DFFX1_RVT \q_reg[120]  ( .D(N123), .CLK(clk), .Q(q[120]) );
  DFFX1_RVT \q_reg[119]  ( .D(N122), .CLK(clk), .Q(q[119]) );
  DFFX1_RVT \q_reg[118]  ( .D(N121), .CLK(clk), .Q(q[118]) );
  DFFX1_RVT \q_reg[117]  ( .D(N120), .CLK(clk), .Q(q[117]) );
  DFFX1_RVT \q_reg[116]  ( .D(N119), .CLK(clk), .Q(q[116]) );
  DFFX1_RVT \q_reg[115]  ( .D(N118), .CLK(clk), .Q(q[115]) );
  DFFX1_RVT \q_reg[114]  ( .D(N117), .CLK(clk), .Q(q[114]) );
  DFFX1_RVT \q_reg[113]  ( .D(N116), .CLK(clk), .Q(q[113]) );
  DFFX1_RVT \q_reg[112]  ( .D(N115), .CLK(clk), .Q(q[112]) );
  DFFX1_RVT \q_reg[111]  ( .D(N114), .CLK(clk), .Q(q[111]) );
  DFFX1_RVT \q_reg[110]  ( .D(N113), .CLK(clk), .Q(q[110]) );
  DFFX1_RVT \q_reg[109]  ( .D(N112), .CLK(clk), .Q(q[109]) );
  DFFX1_RVT \q_reg[108]  ( .D(N111), .CLK(clk), .Q(q[108]) );
  DFFX1_RVT \q_reg[107]  ( .D(N110), .CLK(clk), .Q(q[107]) );
  DFFX1_RVT \q_reg[106]  ( .D(N109), .CLK(clk), .Q(q[106]) );
  DFFX1_RVT \q_reg[105]  ( .D(N108), .CLK(clk), .Q(q[105]) );
  DFFX1_RVT \q_reg[104]  ( .D(N107), .CLK(clk), .Q(q[104]) );
  DFFX1_RVT \q_reg[103]  ( .D(N106), .CLK(clk), .Q(q[103]) );
  DFFX1_RVT \q_reg[102]  ( .D(N105), .CLK(clk), .Q(q[102]) );
  DFFX1_RVT \q_reg[101]  ( .D(N104), .CLK(clk), .Q(q[101]) );
  DFFX1_RVT \q_reg[100]  ( .D(N103), .CLK(clk), .Q(q[100]) );
  DFFX1_RVT \q_reg[99]  ( .D(N102), .CLK(clk), .Q(q[99]) );
  DFFX1_RVT \q_reg[98]  ( .D(N101), .CLK(clk), .Q(q[98]) );
  DFFX1_RVT \q_reg[97]  ( .D(N100), .CLK(clk), .Q(q[97]) );
  DFFX1_RVT \q_reg[96]  ( .D(N99), .CLK(clk), .Q(q[96]) );
  DFFX1_RVT \q_reg[95]  ( .D(N98), .CLK(clk), .Q(q[95]) );
  DFFX1_RVT \q_reg[94]  ( .D(N97), .CLK(clk), .Q(q[94]) );
  DFFX1_RVT \q_reg[93]  ( .D(N96), .CLK(clk), .Q(q[93]) );
  DFFX1_RVT \q_reg[92]  ( .D(N95), .CLK(clk), .Q(q[92]) );
  DFFX1_RVT \q_reg[91]  ( .D(N94), .CLK(clk), .Q(q[91]) );
  DFFX1_RVT \q_reg[90]  ( .D(N93), .CLK(clk), .Q(q[90]) );
  DFFX1_RVT \q_reg[89]  ( .D(N92), .CLK(clk), .Q(q[89]) );
  DFFX1_RVT \q_reg[88]  ( .D(N91), .CLK(clk), .Q(q[88]) );
  DFFX1_RVT \q_reg[87]  ( .D(N90), .CLK(clk), .Q(q[87]) );
  DFFX1_RVT \q_reg[86]  ( .D(N89), .CLK(clk), .Q(q[86]) );
  DFFX1_RVT \q_reg[85]  ( .D(N88), .CLK(clk), .Q(q[85]) );
  DFFX1_RVT \q_reg[84]  ( .D(N87), .CLK(clk), .Q(q[84]) );
  DFFX1_RVT \q_reg[83]  ( .D(N86), .CLK(clk), .Q(q[83]) );
  DFFX1_RVT \q_reg[82]  ( .D(N85), .CLK(clk), .Q(q[82]) );
  DFFX1_RVT \q_reg[81]  ( .D(N84), .CLK(clk), .Q(q[81]) );
  DFFX1_RVT \q_reg[80]  ( .D(N83), .CLK(clk), .Q(q[80]) );
  DFFX1_RVT \q_reg[79]  ( .D(N82), .CLK(clk), .Q(q[79]) );
  DFFX1_RVT \q_reg[78]  ( .D(N81), .CLK(clk), .Q(q[78]) );
  DFFX1_RVT \q_reg[77]  ( .D(N80), .CLK(clk), .Q(q[77]) );
  DFFX1_RVT \q_reg[76]  ( .D(N79), .CLK(clk), .Q(q[76]) );
  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
  AND2X1_RVT U78 ( .A1(din[74]), .A2(n1), .Y(N77) );
  AND2X1_RVT U79 ( .A1(din[75]), .A2(n1), .Y(N78) );
  AND2X1_RVT U80 ( .A1(din[76]), .A2(n1), .Y(N79) );
  AND2X1_RVT U81 ( .A1(din[77]), .A2(n1), .Y(N80) );
  AND2X1_RVT U82 ( .A1(din[78]), .A2(n1), .Y(N81) );
  AND2X1_RVT U83 ( .A1(din[79]), .A2(n1), .Y(N82) );
  AND2X1_RVT U84 ( .A1(din[80]), .A2(n1), .Y(N83) );
  AND2X1_RVT U85 ( .A1(din[81]), .A2(n1), .Y(N84) );
  AND2X1_RVT U86 ( .A1(din[82]), .A2(n1), .Y(N85) );
  AND2X1_RVT U87 ( .A1(din[83]), .A2(n1), .Y(N86) );
  AND2X1_RVT U88 ( .A1(din[84]), .A2(n1), .Y(N87) );
  AND2X1_RVT U89 ( .A1(din[85]), .A2(n1), .Y(N88) );
  AND2X1_RVT U90 ( .A1(din[86]), .A2(n1), .Y(N89) );
  AND2X1_RVT U91 ( .A1(din[87]), .A2(n1), .Y(N90) );
  AND2X1_RVT U92 ( .A1(din[88]), .A2(n1), .Y(N91) );
  AND2X1_RVT U93 ( .A1(din[89]), .A2(n1), .Y(N92) );
  AND2X1_RVT U94 ( .A1(din[90]), .A2(n1), .Y(N93) );
  AND2X1_RVT U95 ( .A1(din[91]), .A2(n1), .Y(N94) );
  AND2X1_RVT U96 ( .A1(din[92]), .A2(n1), .Y(N95) );
  AND2X1_RVT U97 ( .A1(din[93]), .A2(n1), .Y(N96) );
  AND2X1_RVT U98 ( .A1(din[94]), .A2(n1), .Y(N97) );
  AND2X1_RVT U99 ( .A1(din[95]), .A2(n1), .Y(N98) );
  AND2X1_RVT U100 ( .A1(din[96]), .A2(n1), .Y(N99) );
  AND2X1_RVT U101 ( .A1(din[97]), .A2(n1), .Y(N100) );
  AND2X1_RVT U102 ( .A1(din[98]), .A2(n1), .Y(N101) );
  AND2X1_RVT U103 ( .A1(din[99]), .A2(n1), .Y(N102) );
  AND2X1_RVT U104 ( .A1(din[100]), .A2(n1), .Y(N103) );
  AND2X1_RVT U105 ( .A1(din[101]), .A2(n1), .Y(N104) );
  AND2X1_RVT U106 ( .A1(din[102]), .A2(n1), .Y(N105) );
  AND2X1_RVT U107 ( .A1(din[103]), .A2(n1), .Y(N106) );
  AND2X1_RVT U108 ( .A1(din[104]), .A2(n1), .Y(N107) );
  AND2X1_RVT U109 ( .A1(din[105]), .A2(n1), .Y(N108) );
  AND2X1_RVT U110 ( .A1(din[106]), .A2(n1), .Y(N109) );
  AND2X1_RVT U111 ( .A1(din[107]), .A2(n1), .Y(N110) );
  AND2X1_RVT U112 ( .A1(din[108]), .A2(n1), .Y(N111) );
  AND2X1_RVT U113 ( .A1(din[109]), .A2(n1), .Y(N112) );
  AND2X1_RVT U114 ( .A1(din[110]), .A2(n1), .Y(N113) );
  AND2X1_RVT U115 ( .A1(din[111]), .A2(n1), .Y(N114) );
  AND2X1_RVT U116 ( .A1(din[112]), .A2(n1), .Y(N115) );
  AND2X1_RVT U117 ( .A1(din[113]), .A2(n1), .Y(N116) );
  AND2X1_RVT U118 ( .A1(din[114]), .A2(n1), .Y(N117) );
  AND2X1_RVT U119 ( .A1(din[115]), .A2(n1), .Y(N118) );
  AND2X1_RVT U120 ( .A1(din[116]), .A2(n1), .Y(N119) );
  AND2X1_RVT U121 ( .A1(din[117]), .A2(n1), .Y(N120) );
  AND2X1_RVT U122 ( .A1(din[118]), .A2(n1), .Y(N121) );
  AND2X1_RVT U123 ( .A1(din[119]), .A2(n1), .Y(N122) );
  AND2X1_RVT U124 ( .A1(din[120]), .A2(n1), .Y(N123) );
  AND2X1_RVT U125 ( .A1(din[121]), .A2(n1), .Y(N124) );
  AND2X1_RVT U126 ( .A1(din[122]), .A2(n1), .Y(N125) );
  AND2X1_RVT U127 ( .A1(din[123]), .A2(n1), .Y(N126) );
  AND2X1_RVT U128 ( .A1(din[124]), .A2(n1), .Y(N127) );
  AND2X1_RVT U129 ( .A1(din[125]), .A2(n1), .Y(N128) );
  AND2X1_RVT U130 ( .A1(din[126]), .A2(n1), .Y(N129) );
  AND2X1_RVT U131 ( .A1(din[127]), .A2(n1), .Y(N130) );
  AND2X1_RVT U132 ( .A1(din[128]), .A2(n1), .Y(N131) );
  AND2X1_RVT U133 ( .A1(din[129]), .A2(n1), .Y(N132) );
  AND2X1_RVT U134 ( .A1(din[130]), .A2(n1), .Y(N133) );
  AND2X1_RVT U135 ( .A1(din[131]), .A2(n1), .Y(N134) );
  AND2X1_RVT U136 ( .A1(din[132]), .A2(n1), .Y(N135) );
  AND2X1_RVT U137 ( .A1(din[133]), .A2(n1), .Y(N136) );
  AND2X1_RVT U138 ( .A1(din[134]), .A2(n1), .Y(N137) );
  AND2X1_RVT U139 ( .A1(din[135]), .A2(n1), .Y(N138) );
  AND2X1_RVT U140 ( .A1(din[136]), .A2(n1), .Y(N139) );
  AND2X1_RVT U141 ( .A1(din[137]), .A2(n1), .Y(N140) );
  AND2X1_RVT U142 ( .A1(din[138]), .A2(n1), .Y(N141) );
  AND2X1_RVT U143 ( .A1(din[139]), .A2(n1), .Y(N142) );
  AND2X1_RVT U144 ( .A1(din[140]), .A2(n1), .Y(N143) );
  AND2X1_RVT U145 ( .A1(din[141]), .A2(n1), .Y(N144) );
  AND2X1_RVT U146 ( .A1(din[142]), .A2(n1), .Y(N145) );
  AND2X1_RVT U147 ( .A1(din[143]), .A2(n1), .Y(N146) );
  AND2X1_RVT U148 ( .A1(din[144]), .A2(n1), .Y(N147) );
  AND2X1_RVT U149 ( .A1(din[145]), .A2(n1), .Y(N148) );
  AND2X1_RVT U150 ( .A1(din[146]), .A2(n1), .Y(N149) );
  AND2X1_RVT U151 ( .A1(din[147]), .A2(n1), .Y(N150) );
  AND2X1_RVT U152 ( .A1(din[148]), .A2(n1), .Y(N151) );
  AND2X1_RVT U153 ( .A1(din[149]), .A2(n1), .Y(N152) );
  AND2X1_RVT U154 ( .A1(din[150]), .A2(n1), .Y(N153) );
  AND2X1_RVT U155 ( .A1(din[151]), .A2(n1), .Y(N154) );
  AND2X1_RVT U156 ( .A1(din[152]), .A2(n1), .Y(N155) );
  AND2X1_RVT U157 ( .A1(din[153]), .A2(n1), .Y(N156) );
  AND2X1_RVT U158 ( .A1(din[154]), .A2(n1), .Y(N157) );
endmodule


module fpu_in_dp ( fp_data_rdy, fpio_data_px2_116_112, fpio_data_px2_79_72, 
        fpio_data_px2_67_0, inq_fwrd, inq_fwrd_inv, inq_bp, inq_bp_inv, 
        inq_dout, rclk, fp_op_in_7in, inq_id, inq_rnd_mode, inq_fcc, inq_op, 
        inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1, inq_in2_exp_neq_ffs, 
        inq_in2_exp_eq_0, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2, fp_id_in, fp_rnd_mode_in, fp_fcc_in, 
        fp_op_in, fp_src1_in, fp_src2_in, se, si, so );
  input [116:112] fpio_data_px2_116_112;
  input [79:72] fpio_data_px2_79_72;
  input [67:0] fpio_data_px2_67_0;
  input [154:0] inq_dout;
  output [4:0] inq_id;
  output [1:0] inq_rnd_mode;
  output [1:0] inq_fcc;
  output [7:0] inq_op;
  output [63:0] inq_in1;
  output [63:0] inq_in2;
  output [4:0] fp_id_in;
  output [1:0] fp_rnd_mode_in;
  output [1:0] fp_fcc_in;
  output [7:0] fp_op_in;
  output [68:0] fp_src1_in;
  output [68:0] fp_src2_in;
  input fp_data_rdy, inq_fwrd, inq_fwrd_inv, inq_bp, inq_bp_inv, rclk, se, si;
  output fp_op_in_7in, inq_in1_exp_neq_ffs, inq_in1_exp_eq_0,
         inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in2_exp_neq_ffs, inq_in2_exp_eq_0, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, so;
  wire   fp_op_in_7in, clk, fp_srca_53_0_neq_0, fp_srca_50_0_neq_0,
         fp_srca_53_32_neq_0, n35, n36, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n37, n38;
  wire   [63:0] fp_srca_in;
  wire   [68:0] fp_srcb_in;
  wire   [154:0] inq_din_d1;
  assign fp_op_in[7] = fp_op_in_7in;
  assign so = 1'b0;

  clken_buf_0 ckbuf_in_dp ( .clk(clk), .rclk(rclk), .enb_l(1'b0), .tmb_l(1'b0)
         );
  dff_SIZE5_2 i_fp_id_in ( .din(fpio_data_px2_116_112), .clk(clk), .q(fp_id_in), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE8_4 i_fp_op_in ( .din(fpio_data_px2_79_72), .clk(clk), .q({
        fp_op_in_7in, fp_op_in[6:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE2_0 i_fp_fcc_in ( .din(fpio_data_px2_67_0[67:66]), .clk(clk), .q(
        fp_fcc_in), .se(se), .si({1'b0, 1'b0}) );
  dff_SIZE2_2 i_fp_rnd_mode_in ( .din(fpio_data_px2_67_0[65:64]), .clk(clk), 
        .q(fp_rnd_mode_in), .se(se), .si({1'b0, 1'b0}) );
  dff_SIZE64_0 i_fp_srca_in ( .din(fpio_data_px2_67_0[63:0]), .clk(clk), .q(
        fp_srca_in), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE69 i_fp_srcb_in ( .din({n35, n36, fp_srca_53_0_neq_0, 
        fp_srca_50_0_neq_0, fp_srca_53_32_neq_0, fp_srca_in}), .en(fp_data_rdy), .clk(clk), .q(fp_srcb_in), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE155 i_inq_din_d1 ( .din({fp_id_in, fp_rnd_mode_in, fp_fcc_in, 
        fp_op_in_7in, fp_op_in[6:0], fp_src1_in, fp_src2_in}), .clk(clk), .q(
        inq_din_d1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  INVX0_RVT U2 ( .A(fp_srca_50_0_neq_0), .Y(n27) );
  INVX0_RVT U3 ( .A(n28), .Y(n32) );
  OR3X1_RVT U4 ( .A1(n28), .A2(n15), .A3(n14), .Y(fp_srca_50_0_neq_0) );
  INVX0_RVT U5 ( .A(fp_srca_in[52]), .Y(n30) );
  INVX0_RVT U6 ( .A(fp_srca_in[53]), .Y(n29) );
  INVX0_RVT U7 ( .A(fp_op_in[0]), .Y(n17) );
  INVX0_RVT U8 ( .A(fp_srca_in[61]), .Y(n23) );
  INVX0_RVT U9 ( .A(fp_srca_in[62]), .Y(n24) );
  INVX1_RVT U10 ( .A(fp_op_in_7in), .Y(n34) );
  AND2X1_RVT U11 ( .A1(fp_srca_in[54]), .A2(n34), .Y(fp_src1_in[54]) );
  INVX1_RVT U12 ( .A(inq_fwrd_inv), .Y(n33) );
  NOR2X0_RVT U13 ( .A1(inq_bp_inv), .A2(n33), .Y(n38) );
  AND2X1_RVT U14 ( .A1(inq_fwrd_inv), .A2(inq_bp_inv), .Y(n37) );
  AO222X1_RVT U15 ( .A1(n33), .A2(fp_src1_in[54]), .A3(n38), .A4(
        inq_din_d1[123]), .A5(inq_dout[123]), .A6(n37), .Y(inq_in1[54]) );
  AO22X1_RVT U16 ( .A1(fp_op_in_7in), .A2(fp_srca_in[54]), .A3(n34), .A4(
        fp_srcb_in[54]), .Y(fp_src2_in[54]) );
  AO222X1_RVT U17 ( .A1(n33), .A2(fp_src2_in[54]), .A3(inq_din_d1[54]), .A4(
        n38), .A5(n37), .A6(inq_dout[54]), .Y(inq_in2[54]) );
  AO222X1_RVT U18 ( .A1(n33), .A2(fp_op_in[1]), .A3(n38), .A4(inq_din_d1[139]), 
        .A5(inq_dout[139]), .A6(n37), .Y(inq_op[1]) );
  AND2X1_RVT U19 ( .A1(fp_srca_in[52]), .A2(n34), .Y(fp_src1_in[52]) );
  AO222X1_RVT U20 ( .A1(n33), .A2(fp_src1_in[52]), .A3(n38), .A4(
        inq_din_d1[121]), .A5(inq_dout[121]), .A6(n37), .Y(inq_in1[52]) );
  AND2X1_RVT U21 ( .A1(fp_srca_in[53]), .A2(n34), .Y(fp_src1_in[53]) );
  AO222X1_RVT U22 ( .A1(n33), .A2(fp_src1_in[53]), .A3(n38), .A4(
        inq_din_d1[122]), .A5(inq_dout[122]), .A6(n37), .Y(inq_in1[53]) );
  AO222X1_RVT U23 ( .A1(n33), .A2(fp_op_in[0]), .A3(n38), .A4(inq_din_d1[138]), 
        .A5(inq_dout[138]), .A6(n37), .Y(inq_op[0]) );
  AO22X1_RVT U24 ( .A1(fp_op_in_7in), .A2(fp_srca_in[53]), .A3(n34), .A4(
        fp_srcb_in[53]), .Y(fp_src2_in[53]) );
  AO222X1_RVT U25 ( .A1(n33), .A2(fp_src2_in[53]), .A3(inq_din_d1[53]), .A4(
        n38), .A5(n37), .A6(inq_dout[53]), .Y(inq_in2[53]) );
  AO22X1_RVT U26 ( .A1(fp_op_in_7in), .A2(fp_srca_in[52]), .A3(n34), .A4(
        fp_srcb_in[52]), .Y(fp_src2_in[52]) );
  AO222X1_RVT U27 ( .A1(n33), .A2(fp_src2_in[52]), .A3(inq_din_d1[52]), .A4(
        n38), .A5(n37), .A6(inq_dout[52]), .Y(inq_in2[52]) );
  AND2X1_RVT U28 ( .A1(fp_srca_in[0]), .A2(n34), .Y(fp_src1_in[0]) );
  AND2X1_RVT U29 ( .A1(fp_srca_in[2]), .A2(n34), .Y(fp_src1_in[2]) );
  AND2X1_RVT U30 ( .A1(fp_srca_in[3]), .A2(n34), .Y(fp_src1_in[3]) );
  AND2X1_RVT U31 ( .A1(fp_srca_in[4]), .A2(n34), .Y(fp_src1_in[4]) );
  AND2X1_RVT U32 ( .A1(fp_srca_in[5]), .A2(n34), .Y(fp_src1_in[5]) );
  AND2X1_RVT U33 ( .A1(fp_srca_in[6]), .A2(n34), .Y(fp_src1_in[6]) );
  AND2X1_RVT U34 ( .A1(fp_srca_in[7]), .A2(n34), .Y(fp_src1_in[7]) );
  AND2X1_RVT U35 ( .A1(fp_srca_in[8]), .A2(n34), .Y(fp_src1_in[8]) );
  AND2X1_RVT U36 ( .A1(fp_srca_in[9]), .A2(n34), .Y(fp_src1_in[9]) );
  AND2X1_RVT U37 ( .A1(fp_srca_in[10]), .A2(n34), .Y(fp_src1_in[10]) );
  AND2X1_RVT U38 ( .A1(fp_srca_in[11]), .A2(n34), .Y(fp_src1_in[11]) );
  AND2X1_RVT U39 ( .A1(fp_srca_in[12]), .A2(n34), .Y(fp_src1_in[12]) );
  AND2X1_RVT U40 ( .A1(fp_srca_in[13]), .A2(n34), .Y(fp_src1_in[13]) );
  AND2X1_RVT U41 ( .A1(fp_srca_in[1]), .A2(n34), .Y(fp_src1_in[1]) );
  AND2X1_RVT U42 ( .A1(fp_srca_in[38]), .A2(n34), .Y(fp_src1_in[38]) );
  AND2X1_RVT U43 ( .A1(fp_srca_in[37]), .A2(n34), .Y(fp_src1_in[37]) );
  AND2X1_RVT U44 ( .A1(fp_srca_in[36]), .A2(n34), .Y(fp_src1_in[36]) );
  AND2X1_RVT U45 ( .A1(fp_srca_in[35]), .A2(n34), .Y(fp_src1_in[35]) );
  AND2X1_RVT U46 ( .A1(fp_srca_in[34]), .A2(n34), .Y(fp_src1_in[34]) );
  AND2X1_RVT U47 ( .A1(fp_srca_in[33]), .A2(n34), .Y(fp_src1_in[33]) );
  AND2X1_RVT U48 ( .A1(fp_srca_in[32]), .A2(n34), .Y(fp_src1_in[32]) );
  AND2X1_RVT U49 ( .A1(fp_srca_in[31]), .A2(n34), .Y(fp_src1_in[31]) );
  AND2X1_RVT U50 ( .A1(fp_srca_in[30]), .A2(n34), .Y(fp_src1_in[30]) );
  AND2X1_RVT U51 ( .A1(fp_srca_in[29]), .A2(n34), .Y(fp_src1_in[29]) );
  AND2X1_RVT U52 ( .A1(fp_srca_in[28]), .A2(n34), .Y(fp_src1_in[28]) );
  AND2X1_RVT U53 ( .A1(fp_srca_in[27]), .A2(n34), .Y(fp_src1_in[27]) );
  AND2X1_RVT U54 ( .A1(fp_srca_in[26]), .A2(n34), .Y(fp_src1_in[26]) );
  AND2X1_RVT U55 ( .A1(fp_srca_in[25]), .A2(n34), .Y(fp_src1_in[25]) );
  AND2X1_RVT U56 ( .A1(fp_srca_in[24]), .A2(n34), .Y(fp_src1_in[24]) );
  AND2X1_RVT U57 ( .A1(fp_srca_in[23]), .A2(n34), .Y(fp_src1_in[23]) );
  AND2X1_RVT U58 ( .A1(fp_srca_in[22]), .A2(n34), .Y(fp_src1_in[22]) );
  AND2X1_RVT U59 ( .A1(fp_srca_in[21]), .A2(n34), .Y(fp_src1_in[21]) );
  AND2X1_RVT U60 ( .A1(fp_srca_in[20]), .A2(n34), .Y(fp_src1_in[20]) );
  AND2X1_RVT U61 ( .A1(fp_srca_in[19]), .A2(n34), .Y(fp_src1_in[19]) );
  AND2X1_RVT U62 ( .A1(fp_srca_in[18]), .A2(n34), .Y(fp_src1_in[18]) );
  AND2X1_RVT U63 ( .A1(fp_srca_in[17]), .A2(n34), .Y(fp_src1_in[17]) );
  AND2X1_RVT U64 ( .A1(fp_srca_in[16]), .A2(n34), .Y(fp_src1_in[16]) );
  AND2X1_RVT U65 ( .A1(fp_srca_in[15]), .A2(n34), .Y(fp_src1_in[15]) );
  AND2X1_RVT U66 ( .A1(fp_srca_in[14]), .A2(n34), .Y(fp_src1_in[14]) );
  AND2X1_RVT U67 ( .A1(fp_srca_in[39]), .A2(n34), .Y(fp_src1_in[39]) );
  AND2X1_RVT U68 ( .A1(fp_srca_in[47]), .A2(n34), .Y(fp_src1_in[47]) );
  AND2X1_RVT U69 ( .A1(fp_srca_in[40]), .A2(n34), .Y(fp_src1_in[40]) );
  AND2X1_RVT U70 ( .A1(fp_srca_in[41]), .A2(n34), .Y(fp_src1_in[41]) );
  AND2X1_RVT U71 ( .A1(fp_srca_in[42]), .A2(n34), .Y(fp_src1_in[42]) );
  AND2X1_RVT U72 ( .A1(fp_srca_in[43]), .A2(n34), .Y(fp_src1_in[43]) );
  AND2X1_RVT U73 ( .A1(fp_srca_in[44]), .A2(n34), .Y(fp_src1_in[44]) );
  AND2X1_RVT U74 ( .A1(fp_srca_in[45]), .A2(n34), .Y(fp_src1_in[45]) );
  AND2X1_RVT U75 ( .A1(fp_srca_in[46]), .A2(n34), .Y(fp_src1_in[46]) );
  AND2X1_RVT U76 ( .A1(fp_srca_in[48]), .A2(n34), .Y(fp_src1_in[48]) );
  AND2X1_RVT U77 ( .A1(fp_srca_in[49]), .A2(n34), .Y(fp_src1_in[49]) );
  AND2X1_RVT U78 ( .A1(fp_srca_in[50]), .A2(n34), .Y(fp_src1_in[50]) );
  AND2X1_RVT U79 ( .A1(fp_srca_in[59]), .A2(n34), .Y(fp_src1_in[59]) );
  AND2X1_RVT U80 ( .A1(fp_srca_in[58]), .A2(n34), .Y(fp_src1_in[58]) );
  AND2X1_RVT U81 ( .A1(fp_srca_in[62]), .A2(n34), .Y(fp_src1_in[62]) );
  AND2X1_RVT U82 ( .A1(fp_srca_in[57]), .A2(n34), .Y(fp_src1_in[57]) );
  AND2X1_RVT U83 ( .A1(fp_srca_in[56]), .A2(n34), .Y(fp_src1_in[56]) );
  AND2X1_RVT U84 ( .A1(fp_srca_in[55]), .A2(n34), .Y(fp_src1_in[55]) );
  AND2X1_RVT U85 ( .A1(fp_srca_in[61]), .A2(n34), .Y(fp_src1_in[61]) );
  AND2X1_RVT U86 ( .A1(fp_srca_in[60]), .A2(n34), .Y(fp_src1_in[60]) );
  AND2X1_RVT U87 ( .A1(fp_srca_in[63]), .A2(n34), .Y(fp_src1_in[63]) );
  AND2X1_RVT U88 ( .A1(fp_srca_in[51]), .A2(n34), .Y(fp_src1_in[51]) );
  NOR4X1_RVT U89 ( .A1(fp_srca_in[38]), .A2(fp_srca_in[39]), .A3(
        fp_srca_in[40]), .A4(fp_srca_in[41]), .Y(n5) );
  NOR4X1_RVT U90 ( .A1(fp_srca_in[42]), .A2(fp_srca_in[43]), .A3(
        fp_srca_in[44]), .A4(fp_srca_in[45]), .Y(n4) );
  NOR4X1_RVT U91 ( .A1(fp_srca_in[46]), .A2(fp_srca_in[47]), .A3(
        fp_srca_in[48]), .A4(fp_srca_in[49]), .Y(n3) );
  OR4X1_RVT U92 ( .A1(fp_srca_in[34]), .A2(fp_srca_in[35]), .A3(fp_srca_in[36]), .A4(fp_srca_in[37]), .Y(n1) );
  NOR4X1_RVT U93 ( .A1(fp_srca_in[50]), .A2(fp_srca_in[32]), .A3(
        fp_srca_in[33]), .A4(n1), .Y(n2) );
  NAND4X0_RVT U94 ( .A1(n5), .A2(n4), .A3(n3), .A4(n2), .Y(n28) );
  NOR4X1_RVT U95 ( .A1(fp_srca_in[0]), .A2(fp_srca_in[1]), .A3(fp_srca_in[2]), 
        .A4(fp_srca_in[3]), .Y(n9) );
  NOR4X1_RVT U96 ( .A1(fp_srca_in[4]), .A2(fp_srca_in[5]), .A3(fp_srca_in[6]), 
        .A4(fp_srca_in[7]), .Y(n8) );
  NOR4X1_RVT U97 ( .A1(fp_srca_in[8]), .A2(fp_srca_in[9]), .A3(fp_srca_in[10]), 
        .A4(fp_srca_in[11]), .Y(n7) );
  NOR4X1_RVT U98 ( .A1(fp_srca_in[12]), .A2(fp_srca_in[13]), .A3(
        fp_srca_in[14]), .A4(fp_srca_in[15]), .Y(n6) );
  NAND4X0_RVT U99 ( .A1(n9), .A2(n8), .A3(n7), .A4(n6), .Y(n15) );
  NOR4X1_RVT U100 ( .A1(fp_srca_in[20]), .A2(fp_srca_in[21]), .A3(
        fp_srca_in[22]), .A4(fp_srca_in[23]), .Y(n13) );
  NOR4X1_RVT U101 ( .A1(fp_srca_in[16]), .A2(fp_srca_in[17]), .A3(
        fp_srca_in[18]), .A4(fp_srca_in[19]), .Y(n12) );
  NOR4X1_RVT U102 ( .A1(fp_srca_in[28]), .A2(fp_srca_in[29]), .A3(
        fp_srca_in[30]), .A4(fp_srca_in[31]), .Y(n11) );
  NOR4X1_RVT U103 ( .A1(fp_srca_in[24]), .A2(fp_srca_in[25]), .A3(
        fp_srca_in[26]), .A4(fp_srca_in[27]), .Y(n10) );
  NAND4X0_RVT U104 ( .A1(n13), .A2(n12), .A3(n11), .A4(n10), .Y(n14) );
  AND4X1_RVT U105 ( .A1(fp_srca_in[59]), .A2(fp_srca_in[60]), .A3(
        fp_srca_in[61]), .A4(fp_srca_in[62]), .Y(n20) );
  AND4X1_RVT U106 ( .A1(fp_srca_in[55]), .A2(fp_srca_in[56]), .A3(
        fp_srca_in[57]), .A4(fp_srca_in[58]), .Y(n19) );
  NAND3X0_RVT U107 ( .A1(fp_srca_in[52]), .A2(fp_srca_in[53]), .A3(
        fp_srca_in[54]), .Y(n16) );
  NAND2X0_RVT U108 ( .A1(n17), .A2(n16), .Y(n18) );
  NAND3X0_RVT U109 ( .A1(n20), .A2(n19), .A3(n18), .Y(n35) );
  AO222X1_RVT U111 ( .A1(n33), .A2(fp_id_in[4]), .A3(n38), .A4(inq_din_d1[154]), .A5(inq_dout[154]), .A6(n37), .Y(inq_id[4]) );
  AO222X1_RVT U112 ( .A1(n33), .A2(fp_id_in[3]), .A3(n38), .A4(inq_din_d1[153]), .A5(inq_dout[153]), .A6(n37), .Y(inq_id[3]) );
  AO222X1_RVT U113 ( .A1(n33), .A2(fp_id_in[2]), .A3(n38), .A4(inq_din_d1[152]), .A5(inq_dout[152]), .A6(n37), .Y(inq_id[2]) );
  AO222X1_RVT U114 ( .A1(n33), .A2(fp_id_in[1]), .A3(n38), .A4(inq_din_d1[151]), .A5(inq_dout[151]), .A6(n37), .Y(inq_id[1]) );
  AO222X1_RVT U115 ( .A1(n33), .A2(fp_id_in[0]), .A3(n38), .A4(inq_din_d1[150]), .A5(inq_dout[150]), .A6(n37), .Y(inq_id[0]) );
  AO222X1_RVT U116 ( .A1(n33), .A2(fp_rnd_mode_in[1]), .A3(n38), .A4(
        inq_din_d1[149]), .A5(inq_dout[149]), .A6(n37), .Y(inq_rnd_mode[1]) );
  AO222X1_RVT U117 ( .A1(n33), .A2(fp_rnd_mode_in[0]), .A3(n38), .A4(
        inq_din_d1[148]), .A5(inq_dout[148]), .A6(n37), .Y(inq_rnd_mode[0]) );
  AO222X1_RVT U118 ( .A1(n33), .A2(fp_fcc_in[1]), .A3(n38), .A4(
        inq_din_d1[147]), .A5(inq_dout[147]), .A6(n37), .Y(inq_fcc[1]) );
  AO222X1_RVT U119 ( .A1(n33), .A2(fp_fcc_in[0]), .A3(n38), .A4(
        inq_din_d1[146]), .A5(inq_dout[146]), .A6(n37), .Y(inq_fcc[0]) );
  AO222X1_RVT U120 ( .A1(n33), .A2(fp_op_in_7in), .A3(n38), .A4(
        inq_din_d1[145]), .A5(inq_dout[145]), .A6(n37), .Y(inq_op[7]) );
  AO222X1_RVT U121 ( .A1(n33), .A2(fp_op_in[6]), .A3(n38), .A4(inq_din_d1[144]), .A5(inq_dout[144]), .A6(n37), .Y(inq_op[6]) );
  AO222X1_RVT U122 ( .A1(n33), .A2(fp_op_in[5]), .A3(n38), .A4(inq_din_d1[143]), .A5(inq_dout[143]), .A6(n37), .Y(inq_op[5]) );
  AO222X1_RVT U123 ( .A1(n33), .A2(fp_op_in[4]), .A3(n38), .A4(inq_din_d1[142]), .A5(inq_dout[142]), .A6(n37), .Y(inq_op[4]) );
  AO222X1_RVT U124 ( .A1(n33), .A2(fp_op_in[3]), .A3(n38), .A4(inq_din_d1[141]), .A5(inq_dout[141]), .A6(n37), .Y(inq_op[3]) );
  AO222X1_RVT U125 ( .A1(n33), .A2(fp_op_in[2]), .A3(n38), .A4(inq_din_d1[140]), .A5(inq_dout[140]), .A6(n37), .Y(inq_op[2]) );
  OR2X1_RVT U126 ( .A1(n35), .A2(fp_op_in_7in), .Y(fp_src1_in[68]) );
  AO222X1_RVT U127 ( .A1(n33), .A2(fp_src1_in[68]), .A3(inq_din_d1[137]), .A4(
        n38), .A5(n37), .A6(inq_dout[137]), .Y(inq_in1_exp_neq_ffs) );
  OR4X1_RVT U128 ( .A1(fp_srca_in[55]), .A2(fp_srca_in[56]), .A3(
        fp_srca_in[57]), .A4(fp_srca_in[58]), .Y(n26) );
  OR3X2_RVT U129 ( .A1(fp_srca_in[52]), .A2(fp_srca_in[53]), .A3(
        fp_srca_in[54]), .Y(n21) );
  NAND2X0_RVT U130 ( .A1(fp_op_in[1]), .A2(n21), .Y(n22) );
  NAND3X0_RVT U131 ( .A1(n24), .A2(n23), .A3(n22), .Y(n25) );
  NOR4X1_RVT U132 ( .A1(fp_srca_in[59]), .A2(fp_srca_in[60]), .A3(n26), .A4(
        n25), .Y(n36) );
  OR2X1_RVT U133 ( .A1(fp_op_in_7in), .A2(n36), .Y(fp_src1_in[67]) );
  AO222X1_RVT U134 ( .A1(n33), .A2(fp_src1_in[67]), .A3(inq_din_d1[136]), .A4(
        n38), .A5(n37), .A6(inq_dout[136]), .Y(inq_in1_exp_eq_0) );
  INVX1_RVT U135 ( .A(fp_srca_in[51]), .Y(n31) );
  NAND4X0_RVT U136 ( .A1(n27), .A2(n31), .A3(n30), .A4(n29), .Y(
        fp_srca_53_0_neq_0) );
  AND2X1_RVT U137 ( .A1(n34), .A2(fp_srca_53_0_neq_0), .Y(fp_src1_in[66]) );
  AO222X1_RVT U138 ( .A1(n33), .A2(fp_src1_in[66]), .A3(n38), .A4(
        inq_din_d1[135]), .A5(inq_dout[135]), .A6(n37), .Y(inq_in1_53_0_neq_0)
         );
  AND2X1_RVT U139 ( .A1(n34), .A2(fp_srca_50_0_neq_0), .Y(fp_src1_in[65]) );
  AO222X1_RVT U140 ( .A1(n33), .A2(fp_src1_in[65]), .A3(n38), .A4(
        inq_din_d1[134]), .A5(inq_dout[134]), .A6(n37), .Y(inq_in1_50_0_neq_0)
         );
  NAND4X0_RVT U141 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .Y(
        fp_srca_53_32_neq_0) );
  AND2X1_RVT U142 ( .A1(n34), .A2(fp_srca_53_32_neq_0), .Y(fp_src1_in[64]) );
  AO222X1_RVT U143 ( .A1(n33), .A2(fp_src1_in[64]), .A3(n38), .A4(
        inq_din_d1[133]), .A5(inq_dout[133]), .A6(n37), .Y(inq_in1_53_32_neq_0) );
  AO222X1_RVT U144 ( .A1(n33), .A2(fp_src1_in[63]), .A3(n38), .A4(
        inq_din_d1[132]), .A5(inq_dout[132]), .A6(n37), .Y(inq_in1[63]) );
  AO222X1_RVT U145 ( .A1(n33), .A2(fp_src1_in[62]), .A3(n38), .A4(
        inq_din_d1[131]), .A5(inq_dout[131]), .A6(n37), .Y(inq_in1[62]) );
  AO222X1_RVT U146 ( .A1(n33), .A2(fp_src1_in[61]), .A3(n38), .A4(
        inq_din_d1[130]), .A5(inq_dout[130]), .A6(n37), .Y(inq_in1[61]) );
  AO222X1_RVT U147 ( .A1(n33), .A2(fp_src1_in[60]), .A3(n38), .A4(
        inq_din_d1[129]), .A5(inq_dout[129]), .A6(n37), .Y(inq_in1[60]) );
  AO222X1_RVT U148 ( .A1(n33), .A2(fp_src1_in[59]), .A3(n38), .A4(
        inq_din_d1[128]), .A5(inq_dout[128]), .A6(n37), .Y(inq_in1[59]) );
  AO222X1_RVT U149 ( .A1(n33), .A2(fp_src1_in[58]), .A3(n38), .A4(
        inq_din_d1[127]), .A5(inq_dout[127]), .A6(n37), .Y(inq_in1[58]) );
  AO222X1_RVT U150 ( .A1(n33), .A2(fp_src1_in[57]), .A3(n38), .A4(
        inq_din_d1[126]), .A5(inq_dout[126]), .A6(n37), .Y(inq_in1[57]) );
  AO222X1_RVT U151 ( .A1(n33), .A2(fp_src1_in[56]), .A3(n38), .A4(
        inq_din_d1[125]), .A5(inq_dout[125]), .A6(n37), .Y(inq_in1[56]) );
  AO222X1_RVT U152 ( .A1(n33), .A2(fp_src1_in[55]), .A3(n38), .A4(
        inq_din_d1[124]), .A5(inq_dout[124]), .A6(n37), .Y(inq_in1[55]) );
  AO222X1_RVT U153 ( .A1(n33), .A2(fp_src1_in[51]), .A3(n38), .A4(
        inq_din_d1[120]), .A5(inq_dout[120]), .A6(n37), .Y(inq_in1[51]) );
  AO222X1_RVT U154 ( .A1(n33), .A2(fp_src1_in[50]), .A3(n38), .A4(
        inq_din_d1[119]), .A5(inq_dout[119]), .A6(n37), .Y(inq_in1[50]) );
  AO222X1_RVT U155 ( .A1(n33), .A2(fp_src1_in[49]), .A3(n38), .A4(
        inq_din_d1[118]), .A5(inq_dout[118]), .A6(n37), .Y(inq_in1[49]) );
  AO222X1_RVT U156 ( .A1(n33), .A2(fp_src1_in[48]), .A3(n38), .A4(
        inq_din_d1[117]), .A5(inq_dout[117]), .A6(n37), .Y(inq_in1[48]) );
  AO222X1_RVT U157 ( .A1(n33), .A2(fp_src1_in[47]), .A3(n38), .A4(
        inq_din_d1[116]), .A5(inq_dout[116]), .A6(n37), .Y(inq_in1[47]) );
  AO222X1_RVT U158 ( .A1(n33), .A2(fp_src1_in[46]), .A3(n38), .A4(
        inq_din_d1[115]), .A5(inq_dout[115]), .A6(n37), .Y(inq_in1[46]) );
  AO222X1_RVT U159 ( .A1(n33), .A2(fp_src1_in[45]), .A3(n38), .A4(
        inq_din_d1[114]), .A5(inq_dout[114]), .A6(n37), .Y(inq_in1[45]) );
  AO222X1_RVT U160 ( .A1(n33), .A2(fp_src1_in[44]), .A3(n38), .A4(
        inq_din_d1[113]), .A5(inq_dout[113]), .A6(n37), .Y(inq_in1[44]) );
  AO222X1_RVT U161 ( .A1(n33), .A2(fp_src1_in[43]), .A3(n38), .A4(
        inq_din_d1[112]), .A5(inq_dout[112]), .A6(n37), .Y(inq_in1[43]) );
  AO222X1_RVT U162 ( .A1(n33), .A2(fp_src1_in[42]), .A3(n38), .A4(
        inq_din_d1[111]), .A5(inq_dout[111]), .A6(n37), .Y(inq_in1[42]) );
  AO222X1_RVT U163 ( .A1(n33), .A2(fp_src1_in[41]), .A3(n38), .A4(
        inq_din_d1[110]), .A5(inq_dout[110]), .A6(n37), .Y(inq_in1[41]) );
  AO222X1_RVT U164 ( .A1(n33), .A2(fp_src1_in[40]), .A3(n38), .A4(
        inq_din_d1[109]), .A5(inq_dout[109]), .A6(n37), .Y(inq_in1[40]) );
  AO222X1_RVT U165 ( .A1(n33), .A2(fp_src1_in[39]), .A3(n38), .A4(
        inq_din_d1[108]), .A5(inq_dout[108]), .A6(n37), .Y(inq_in1[39]) );
  AO222X1_RVT U166 ( .A1(n33), .A2(fp_src1_in[38]), .A3(n38), .A4(
        inq_din_d1[107]), .A5(inq_dout[107]), .A6(n37), .Y(inq_in1[38]) );
  AO222X1_RVT U167 ( .A1(n33), .A2(fp_src1_in[37]), .A3(n38), .A4(
        inq_din_d1[106]), .A5(inq_dout[106]), .A6(n37), .Y(inq_in1[37]) );
  AO222X1_RVT U168 ( .A1(n33), .A2(fp_src1_in[36]), .A3(n38), .A4(
        inq_din_d1[105]), .A5(inq_dout[105]), .A6(n37), .Y(inq_in1[36]) );
  AO222X1_RVT U169 ( .A1(n33), .A2(fp_src1_in[35]), .A3(n38), .A4(
        inq_din_d1[104]), .A5(inq_dout[104]), .A6(n37), .Y(inq_in1[35]) );
  AO222X1_RVT U170 ( .A1(n33), .A2(fp_src1_in[34]), .A3(n38), .A4(
        inq_din_d1[103]), .A5(inq_dout[103]), .A6(n37), .Y(inq_in1[34]) );
  AO222X1_RVT U171 ( .A1(n33), .A2(fp_src1_in[33]), .A3(n38), .A4(
        inq_din_d1[102]), .A5(inq_dout[102]), .A6(n37), .Y(inq_in1[33]) );
  AO222X1_RVT U172 ( .A1(n33), .A2(fp_src1_in[32]), .A3(n38), .A4(
        inq_din_d1[101]), .A5(inq_dout[101]), .A6(n37), .Y(inq_in1[32]) );
  AO222X1_RVT U173 ( .A1(n33), .A2(fp_src1_in[31]), .A3(n38), .A4(
        inq_din_d1[100]), .A5(inq_dout[100]), .A6(n37), .Y(inq_in1[31]) );
  AO222X1_RVT U174 ( .A1(n33), .A2(fp_src1_in[30]), .A3(n38), .A4(
        inq_din_d1[99]), .A5(inq_dout[99]), .A6(n37), .Y(inq_in1[30]) );
  AO222X1_RVT U175 ( .A1(n33), .A2(fp_src1_in[29]), .A3(n38), .A4(
        inq_din_d1[98]), .A5(inq_dout[98]), .A6(n37), .Y(inq_in1[29]) );
  AO222X1_RVT U176 ( .A1(n33), .A2(fp_src1_in[28]), .A3(n38), .A4(
        inq_din_d1[97]), .A5(inq_dout[97]), .A6(n37), .Y(inq_in1[28]) );
  AO222X1_RVT U177 ( .A1(n33), .A2(fp_src1_in[27]), .A3(n38), .A4(
        inq_din_d1[96]), .A5(inq_dout[96]), .A6(n37), .Y(inq_in1[27]) );
  AO222X1_RVT U178 ( .A1(n33), .A2(fp_src1_in[26]), .A3(n38), .A4(
        inq_din_d1[95]), .A5(inq_dout[95]), .A6(n37), .Y(inq_in1[26]) );
  AO222X1_RVT U179 ( .A1(n33), .A2(fp_src1_in[25]), .A3(n38), .A4(
        inq_din_d1[94]), .A5(inq_dout[94]), .A6(n37), .Y(inq_in1[25]) );
  AO222X1_RVT U180 ( .A1(n33), .A2(fp_src1_in[24]), .A3(n38), .A4(
        inq_din_d1[93]), .A5(inq_dout[93]), .A6(n37), .Y(inq_in1[24]) );
  AO222X1_RVT U181 ( .A1(n33), .A2(fp_src1_in[23]), .A3(n38), .A4(
        inq_din_d1[92]), .A5(inq_dout[92]), .A6(n37), .Y(inq_in1[23]) );
  AO222X1_RVT U182 ( .A1(n33), .A2(fp_src1_in[22]), .A3(n38), .A4(
        inq_din_d1[91]), .A5(inq_dout[91]), .A6(n37), .Y(inq_in1[22]) );
  AO222X1_RVT U183 ( .A1(n33), .A2(fp_src1_in[21]), .A3(n38), .A4(
        inq_din_d1[90]), .A5(inq_dout[90]), .A6(n37), .Y(inq_in1[21]) );
  AO222X1_RVT U184 ( .A1(n33), .A2(fp_src1_in[20]), .A3(n38), .A4(
        inq_din_d1[89]), .A5(inq_dout[89]), .A6(n37), .Y(inq_in1[20]) );
  AO222X1_RVT U185 ( .A1(n33), .A2(fp_src1_in[19]), .A3(n38), .A4(
        inq_din_d1[88]), .A5(inq_dout[88]), .A6(n37), .Y(inq_in1[19]) );
  AO222X1_RVT U186 ( .A1(n33), .A2(fp_src1_in[18]), .A3(n38), .A4(
        inq_din_d1[87]), .A5(inq_dout[87]), .A6(n37), .Y(inq_in1[18]) );
  AO222X1_RVT U187 ( .A1(n33), .A2(fp_src1_in[17]), .A3(n38), .A4(
        inq_din_d1[86]), .A5(inq_dout[86]), .A6(n37), .Y(inq_in1[17]) );
  AO222X1_RVT U188 ( .A1(n33), .A2(fp_src1_in[16]), .A3(n38), .A4(
        inq_din_d1[85]), .A5(inq_dout[85]), .A6(n37), .Y(inq_in1[16]) );
  AO222X1_RVT U189 ( .A1(n33), .A2(fp_src1_in[15]), .A3(n38), .A4(
        inq_din_d1[84]), .A5(inq_dout[84]), .A6(n37), .Y(inq_in1[15]) );
  AO222X1_RVT U190 ( .A1(n33), .A2(fp_src1_in[14]), .A3(n38), .A4(
        inq_din_d1[83]), .A5(inq_dout[83]), .A6(n37), .Y(inq_in1[14]) );
  AO222X1_RVT U191 ( .A1(n33), .A2(fp_src1_in[13]), .A3(n38), .A4(
        inq_din_d1[82]), .A5(inq_dout[82]), .A6(n37), .Y(inq_in1[13]) );
  AO222X1_RVT U192 ( .A1(n33), .A2(fp_src1_in[12]), .A3(n38), .A4(
        inq_din_d1[81]), .A5(inq_dout[81]), .A6(n37), .Y(inq_in1[12]) );
  AO222X1_RVT U193 ( .A1(n33), .A2(fp_src1_in[11]), .A3(n38), .A4(
        inq_din_d1[80]), .A5(inq_dout[80]), .A6(n37), .Y(inq_in1[11]) );
  AO222X1_RVT U194 ( .A1(n33), .A2(fp_src1_in[10]), .A3(n38), .A4(
        inq_din_d1[79]), .A5(inq_dout[79]), .A6(n37), .Y(inq_in1[10]) );
  AO222X1_RVT U195 ( .A1(n33), .A2(fp_src1_in[9]), .A3(n38), .A4(
        inq_din_d1[78]), .A5(inq_dout[78]), .A6(n37), .Y(inq_in1[9]) );
  AO222X1_RVT U196 ( .A1(n33), .A2(fp_src1_in[8]), .A3(n38), .A4(
        inq_din_d1[77]), .A5(inq_dout[77]), .A6(n37), .Y(inq_in1[8]) );
  AO222X1_RVT U197 ( .A1(n33), .A2(fp_src1_in[7]), .A3(n38), .A4(
        inq_din_d1[76]), .A5(inq_dout[76]), .A6(n37), .Y(inq_in1[7]) );
  AO222X1_RVT U198 ( .A1(n33), .A2(fp_src1_in[6]), .A3(n38), .A4(
        inq_din_d1[75]), .A5(inq_dout[75]), .A6(n37), .Y(inq_in1[6]) );
  AO222X1_RVT U199 ( .A1(n33), .A2(fp_src1_in[5]), .A3(n38), .A4(
        inq_din_d1[74]), .A5(inq_dout[74]), .A6(n37), .Y(inq_in1[5]) );
  AO222X1_RVT U200 ( .A1(n33), .A2(fp_src1_in[4]), .A3(n38), .A4(
        inq_din_d1[73]), .A5(inq_dout[73]), .A6(n37), .Y(inq_in1[4]) );
  AO222X1_RVT U201 ( .A1(n33), .A2(fp_src1_in[3]), .A3(n38), .A4(
        inq_din_d1[72]), .A5(inq_dout[72]), .A6(n37), .Y(inq_in1[3]) );
  AO222X1_RVT U202 ( .A1(n33), .A2(fp_src1_in[2]), .A3(n38), .A4(
        inq_din_d1[71]), .A5(inq_dout[71]), .A6(n37), .Y(inq_in1[2]) );
  AO222X1_RVT U203 ( .A1(n33), .A2(fp_src1_in[1]), .A3(n38), .A4(
        inq_din_d1[70]), .A5(inq_dout[70]), .A6(n37), .Y(inq_in1[1]) );
  AO222X1_RVT U204 ( .A1(n33), .A2(fp_src1_in[0]), .A3(n38), .A4(
        inq_din_d1[69]), .A5(inq_dout[69]), .A6(n37), .Y(inq_in1[0]) );
  AO22X1_RVT U205 ( .A1(fp_op_in_7in), .A2(n35), .A3(n34), .A4(fp_srcb_in[68]), 
        .Y(fp_src2_in[68]) );
  AO222X1_RVT U206 ( .A1(n33), .A2(fp_src2_in[68]), .A3(n38), .A4(
        inq_din_d1[68]), .A5(inq_dout[68]), .A6(n37), .Y(inq_in2_exp_neq_ffs)
         );
  AO22X1_RVT U207 ( .A1(fp_op_in_7in), .A2(n36), .A3(n34), .A4(fp_srcb_in[67]), 
        .Y(fp_src2_in[67]) );
  AO222X1_RVT U208 ( .A1(n33), .A2(fp_src2_in[67]), .A3(inq_din_d1[67]), .A4(
        n38), .A5(n37), .A6(inq_dout[67]), .Y(inq_in2_exp_eq_0) );
  AO22X1_RVT U209 ( .A1(fp_op_in_7in), .A2(fp_srca_53_0_neq_0), .A3(n34), .A4(
        fp_srcb_in[66]), .Y(fp_src2_in[66]) );
  AO222X1_RVT U210 ( .A1(n33), .A2(fp_src2_in[66]), .A3(n37), .A4(inq_dout[66]), .A5(n38), .A6(inq_din_d1[66]), .Y(inq_in2_53_0_neq_0) );
  AO22X1_RVT U211 ( .A1(fp_op_in_7in), .A2(fp_srca_50_0_neq_0), .A3(n34), .A4(
        fp_srcb_in[65]), .Y(fp_src2_in[65]) );
  AO222X1_RVT U212 ( .A1(n33), .A2(fp_src2_in[65]), .A3(n38), .A4(
        inq_din_d1[65]), .A5(inq_dout[65]), .A6(n37), .Y(inq_in2_50_0_neq_0)
         );
  AO22X1_RVT U213 ( .A1(fp_op_in_7in), .A2(fp_srca_53_32_neq_0), .A3(n34), 
        .A4(fp_srcb_in[64]), .Y(fp_src2_in[64]) );
  AO222X1_RVT U214 ( .A1(n33), .A2(fp_src2_in[64]), .A3(n38), .A4(
        inq_din_d1[64]), .A5(inq_dout[64]), .A6(n37), .Y(inq_in2_53_32_neq_0)
         );
  AO22X1_RVT U215 ( .A1(fp_op_in_7in), .A2(fp_srca_in[63]), .A3(n34), .A4(
        fp_srcb_in[63]), .Y(fp_src2_in[63]) );
  AO222X1_RVT U216 ( .A1(n33), .A2(fp_src2_in[63]), .A3(inq_din_d1[63]), .A4(
        n38), .A5(n37), .A6(inq_dout[63]), .Y(inq_in2[63]) );
  AO22X1_RVT U217 ( .A1(fp_op_in_7in), .A2(fp_srca_in[62]), .A3(n34), .A4(
        fp_srcb_in[62]), .Y(fp_src2_in[62]) );
  AO222X1_RVT U218 ( .A1(n33), .A2(fp_src2_in[62]), .A3(inq_din_d1[62]), .A4(
        n38), .A5(n37), .A6(inq_dout[62]), .Y(inq_in2[62]) );
  AO22X1_RVT U219 ( .A1(fp_op_in_7in), .A2(fp_srca_in[61]), .A3(n34), .A4(
        fp_srcb_in[61]), .Y(fp_src2_in[61]) );
  AO222X1_RVT U220 ( .A1(n33), .A2(fp_src2_in[61]), .A3(inq_din_d1[61]), .A4(
        n38), .A5(n37), .A6(inq_dout[61]), .Y(inq_in2[61]) );
  AO22X1_RVT U221 ( .A1(fp_op_in_7in), .A2(fp_srca_in[60]), .A3(n34), .A4(
        fp_srcb_in[60]), .Y(fp_src2_in[60]) );
  AO222X1_RVT U222 ( .A1(n33), .A2(fp_src2_in[60]), .A3(inq_din_d1[60]), .A4(
        n38), .A5(n37), .A6(inq_dout[60]), .Y(inq_in2[60]) );
  AO22X1_RVT U223 ( .A1(fp_op_in_7in), .A2(fp_srca_in[59]), .A3(n34), .A4(
        fp_srcb_in[59]), .Y(fp_src2_in[59]) );
  AO222X1_RVT U224 ( .A1(n33), .A2(fp_src2_in[59]), .A3(inq_din_d1[59]), .A4(
        n38), .A5(n37), .A6(inq_dout[59]), .Y(inq_in2[59]) );
  AO22X1_RVT U225 ( .A1(fp_op_in_7in), .A2(fp_srca_in[58]), .A3(n34), .A4(
        fp_srcb_in[58]), .Y(fp_src2_in[58]) );
  AO222X1_RVT U226 ( .A1(n33), .A2(fp_src2_in[58]), .A3(inq_din_d1[58]), .A4(
        n38), .A5(n37), .A6(inq_dout[58]), .Y(inq_in2[58]) );
  AO22X1_RVT U227 ( .A1(fp_op_in_7in), .A2(fp_srca_in[57]), .A3(n34), .A4(
        fp_srcb_in[57]), .Y(fp_src2_in[57]) );
  AO222X1_RVT U228 ( .A1(n33), .A2(fp_src2_in[57]), .A3(inq_din_d1[57]), .A4(
        n38), .A5(n37), .A6(inq_dout[57]), .Y(inq_in2[57]) );
  AO22X1_RVT U229 ( .A1(fp_op_in_7in), .A2(fp_srca_in[56]), .A3(n34), .A4(
        fp_srcb_in[56]), .Y(fp_src2_in[56]) );
  AO222X1_RVT U230 ( .A1(n33), .A2(fp_src2_in[56]), .A3(inq_din_d1[56]), .A4(
        n38), .A5(n37), .A6(inq_dout[56]), .Y(inq_in2[56]) );
  AO22X1_RVT U231 ( .A1(fp_op_in_7in), .A2(fp_srca_in[55]), .A3(n34), .A4(
        fp_srcb_in[55]), .Y(fp_src2_in[55]) );
  AO222X1_RVT U232 ( .A1(n33), .A2(fp_src2_in[55]), .A3(inq_din_d1[55]), .A4(
        n38), .A5(n37), .A6(inq_dout[55]), .Y(inq_in2[55]) );
  AO22X1_RVT U233 ( .A1(fp_op_in_7in), .A2(fp_srca_in[51]), .A3(n34), .A4(
        fp_srcb_in[51]), .Y(fp_src2_in[51]) );
  AO222X1_RVT U234 ( .A1(n33), .A2(fp_src2_in[51]), .A3(inq_din_d1[51]), .A4(
        n38), .A5(n37), .A6(inq_dout[51]), .Y(inq_in2[51]) );
  AO22X1_RVT U235 ( .A1(fp_op_in_7in), .A2(fp_srca_in[50]), .A3(n34), .A4(
        fp_srcb_in[50]), .Y(fp_src2_in[50]) );
  AO222X1_RVT U236 ( .A1(n33), .A2(fp_src2_in[50]), .A3(inq_din_d1[50]), .A4(
        n38), .A5(n37), .A6(inq_dout[50]), .Y(inq_in2[50]) );
  AO22X1_RVT U237 ( .A1(fp_op_in_7in), .A2(fp_srca_in[49]), .A3(n34), .A4(
        fp_srcb_in[49]), .Y(fp_src2_in[49]) );
  AO222X1_RVT U238 ( .A1(n33), .A2(fp_src2_in[49]), .A3(inq_din_d1[49]), .A4(
        n38), .A5(n37), .A6(inq_dout[49]), .Y(inq_in2[49]) );
  AO22X1_RVT U239 ( .A1(fp_op_in_7in), .A2(fp_srca_in[48]), .A3(n34), .A4(
        fp_srcb_in[48]), .Y(fp_src2_in[48]) );
  AO222X1_RVT U240 ( .A1(n33), .A2(fp_src2_in[48]), .A3(inq_din_d1[48]), .A4(
        n38), .A5(n37), .A6(inq_dout[48]), .Y(inq_in2[48]) );
  AO22X1_RVT U241 ( .A1(fp_op_in_7in), .A2(fp_srca_in[47]), .A3(n34), .A4(
        fp_srcb_in[47]), .Y(fp_src2_in[47]) );
  AO222X1_RVT U242 ( .A1(n33), .A2(fp_src2_in[47]), .A3(inq_din_d1[47]), .A4(
        n38), .A5(n37), .A6(inq_dout[47]), .Y(inq_in2[47]) );
  AO22X1_RVT U243 ( .A1(fp_op_in_7in), .A2(fp_srca_in[46]), .A3(n34), .A4(
        fp_srcb_in[46]), .Y(fp_src2_in[46]) );
  AO222X1_RVT U244 ( .A1(n33), .A2(fp_src2_in[46]), .A3(inq_din_d1[46]), .A4(
        n38), .A5(n37), .A6(inq_dout[46]), .Y(inq_in2[46]) );
  AO22X1_RVT U245 ( .A1(fp_op_in_7in), .A2(fp_srca_in[45]), .A3(n34), .A4(
        fp_srcb_in[45]), .Y(fp_src2_in[45]) );
  AO222X1_RVT U246 ( .A1(n33), .A2(fp_src2_in[45]), .A3(inq_din_d1[45]), .A4(
        n38), .A5(n37), .A6(inq_dout[45]), .Y(inq_in2[45]) );
  AO22X1_RVT U247 ( .A1(fp_op_in_7in), .A2(fp_srca_in[44]), .A3(n34), .A4(
        fp_srcb_in[44]), .Y(fp_src2_in[44]) );
  AO222X1_RVT U248 ( .A1(n33), .A2(fp_src2_in[44]), .A3(inq_din_d1[44]), .A4(
        n38), .A5(n37), .A6(inq_dout[44]), .Y(inq_in2[44]) );
  AO22X1_RVT U249 ( .A1(fp_op_in_7in), .A2(fp_srca_in[43]), .A3(n34), .A4(
        fp_srcb_in[43]), .Y(fp_src2_in[43]) );
  AO222X1_RVT U250 ( .A1(n33), .A2(fp_src2_in[43]), .A3(inq_din_d1[43]), .A4(
        n38), .A5(n37), .A6(inq_dout[43]), .Y(inq_in2[43]) );
  AO22X1_RVT U251 ( .A1(fp_op_in_7in), .A2(fp_srca_in[42]), .A3(n34), .A4(
        fp_srcb_in[42]), .Y(fp_src2_in[42]) );
  AO222X1_RVT U252 ( .A1(n33), .A2(fp_src2_in[42]), .A3(inq_din_d1[42]), .A4(
        n38), .A5(n37), .A6(inq_dout[42]), .Y(inq_in2[42]) );
  AO22X1_RVT U253 ( .A1(fp_op_in_7in), .A2(fp_srca_in[41]), .A3(n34), .A4(
        fp_srcb_in[41]), .Y(fp_src2_in[41]) );
  AO222X1_RVT U254 ( .A1(n33), .A2(fp_src2_in[41]), .A3(inq_din_d1[41]), .A4(
        n38), .A5(n37), .A6(inq_dout[41]), .Y(inq_in2[41]) );
  AO22X1_RVT U255 ( .A1(fp_op_in_7in), .A2(fp_srca_in[40]), .A3(n34), .A4(
        fp_srcb_in[40]), .Y(fp_src2_in[40]) );
  AO222X1_RVT U256 ( .A1(n33), .A2(fp_src2_in[40]), .A3(inq_din_d1[40]), .A4(
        n38), .A5(n37), .A6(inq_dout[40]), .Y(inq_in2[40]) );
  AO22X1_RVT U257 ( .A1(fp_op_in_7in), .A2(fp_srca_in[39]), .A3(n34), .A4(
        fp_srcb_in[39]), .Y(fp_src2_in[39]) );
  AO222X1_RVT U258 ( .A1(n33), .A2(fp_src2_in[39]), .A3(inq_din_d1[39]), .A4(
        n38), .A5(n37), .A6(inq_dout[39]), .Y(inq_in2[39]) );
  AO22X1_RVT U259 ( .A1(fp_op_in_7in), .A2(fp_srca_in[38]), .A3(n34), .A4(
        fp_srcb_in[38]), .Y(fp_src2_in[38]) );
  AO222X1_RVT U260 ( .A1(n33), .A2(fp_src2_in[38]), .A3(inq_din_d1[38]), .A4(
        n38), .A5(n37), .A6(inq_dout[38]), .Y(inq_in2[38]) );
  AO22X1_RVT U261 ( .A1(fp_op_in_7in), .A2(fp_srca_in[37]), .A3(n34), .A4(
        fp_srcb_in[37]), .Y(fp_src2_in[37]) );
  AO222X1_RVT U262 ( .A1(n33), .A2(fp_src2_in[37]), .A3(inq_din_d1[37]), .A4(
        n38), .A5(n37), .A6(inq_dout[37]), .Y(inq_in2[37]) );
  AO22X1_RVT U263 ( .A1(fp_op_in_7in), .A2(fp_srca_in[36]), .A3(n34), .A4(
        fp_srcb_in[36]), .Y(fp_src2_in[36]) );
  AO222X1_RVT U264 ( .A1(n33), .A2(fp_src2_in[36]), .A3(inq_din_d1[36]), .A4(
        n38), .A5(n37), .A6(inq_dout[36]), .Y(inq_in2[36]) );
  AO22X1_RVT U265 ( .A1(fp_op_in_7in), .A2(fp_srca_in[35]), .A3(n34), .A4(
        fp_srcb_in[35]), .Y(fp_src2_in[35]) );
  AO222X1_RVT U266 ( .A1(n33), .A2(fp_src2_in[35]), .A3(inq_din_d1[35]), .A4(
        n38), .A5(n37), .A6(inq_dout[35]), .Y(inq_in2[35]) );
  AO22X1_RVT U267 ( .A1(fp_op_in_7in), .A2(fp_srca_in[34]), .A3(n34), .A4(
        fp_srcb_in[34]), .Y(fp_src2_in[34]) );
  AO222X1_RVT U268 ( .A1(n33), .A2(fp_src2_in[34]), .A3(inq_din_d1[34]), .A4(
        n38), .A5(n37), .A6(inq_dout[34]), .Y(inq_in2[34]) );
  AO22X1_RVT U269 ( .A1(fp_op_in_7in), .A2(fp_srca_in[33]), .A3(n34), .A4(
        fp_srcb_in[33]), .Y(fp_src2_in[33]) );
  AO222X1_RVT U270 ( .A1(n33), .A2(fp_src2_in[33]), .A3(inq_din_d1[33]), .A4(
        n38), .A5(n37), .A6(inq_dout[33]), .Y(inq_in2[33]) );
  AO22X1_RVT U271 ( .A1(fp_op_in_7in), .A2(fp_srca_in[32]), .A3(n34), .A4(
        fp_srcb_in[32]), .Y(fp_src2_in[32]) );
  AO222X1_RVT U272 ( .A1(n33), .A2(fp_src2_in[32]), .A3(inq_din_d1[32]), .A4(
        n38), .A5(n37), .A6(inq_dout[32]), .Y(inq_in2[32]) );
  AO22X1_RVT U273 ( .A1(fp_op_in_7in), .A2(fp_srca_in[31]), .A3(n34), .A4(
        fp_srcb_in[31]), .Y(fp_src2_in[31]) );
  AO222X1_RVT U274 ( .A1(n33), .A2(fp_src2_in[31]), .A3(inq_din_d1[31]), .A4(
        n38), .A5(n37), .A6(inq_dout[31]), .Y(inq_in2[31]) );
  AO22X1_RVT U275 ( .A1(fp_op_in_7in), .A2(fp_srca_in[30]), .A3(n34), .A4(
        fp_srcb_in[30]), .Y(fp_src2_in[30]) );
  AO222X1_RVT U276 ( .A1(n33), .A2(fp_src2_in[30]), .A3(inq_din_d1[30]), .A4(
        n38), .A5(n37), .A6(inq_dout[30]), .Y(inq_in2[30]) );
  AO22X1_RVT U277 ( .A1(fp_op_in_7in), .A2(fp_srca_in[29]), .A3(n34), .A4(
        fp_srcb_in[29]), .Y(fp_src2_in[29]) );
  AO222X1_RVT U278 ( .A1(n33), .A2(fp_src2_in[29]), .A3(inq_din_d1[29]), .A4(
        n38), .A5(n37), .A6(inq_dout[29]), .Y(inq_in2[29]) );
  AO22X1_RVT U279 ( .A1(fp_op_in_7in), .A2(fp_srca_in[28]), .A3(n34), .A4(
        fp_srcb_in[28]), .Y(fp_src2_in[28]) );
  AO222X1_RVT U280 ( .A1(n33), .A2(fp_src2_in[28]), .A3(inq_din_d1[28]), .A4(
        n38), .A5(n37), .A6(inq_dout[28]), .Y(inq_in2[28]) );
  AO22X1_RVT U281 ( .A1(fp_op_in_7in), .A2(fp_srca_in[27]), .A3(n34), .A4(
        fp_srcb_in[27]), .Y(fp_src2_in[27]) );
  AO222X1_RVT U282 ( .A1(n33), .A2(fp_src2_in[27]), .A3(inq_din_d1[27]), .A4(
        n38), .A5(n37), .A6(inq_dout[27]), .Y(inq_in2[27]) );
  AO22X1_RVT U283 ( .A1(fp_op_in_7in), .A2(fp_srca_in[26]), .A3(n34), .A4(
        fp_srcb_in[26]), .Y(fp_src2_in[26]) );
  AO222X1_RVT U284 ( .A1(n33), .A2(fp_src2_in[26]), .A3(inq_din_d1[26]), .A4(
        n38), .A5(n37), .A6(inq_dout[26]), .Y(inq_in2[26]) );
  AO22X1_RVT U285 ( .A1(fp_op_in_7in), .A2(fp_srca_in[25]), .A3(n34), .A4(
        fp_srcb_in[25]), .Y(fp_src2_in[25]) );
  AO222X1_RVT U286 ( .A1(n33), .A2(fp_src2_in[25]), .A3(inq_din_d1[25]), .A4(
        n38), .A5(n37), .A6(inq_dout[25]), .Y(inq_in2[25]) );
  AO22X1_RVT U287 ( .A1(fp_op_in_7in), .A2(fp_srca_in[24]), .A3(n34), .A4(
        fp_srcb_in[24]), .Y(fp_src2_in[24]) );
  AO222X1_RVT U288 ( .A1(n33), .A2(fp_src2_in[24]), .A3(inq_din_d1[24]), .A4(
        n38), .A5(n37), .A6(inq_dout[24]), .Y(inq_in2[24]) );
  AO22X1_RVT U289 ( .A1(fp_op_in_7in), .A2(fp_srca_in[23]), .A3(n34), .A4(
        fp_srcb_in[23]), .Y(fp_src2_in[23]) );
  AO222X1_RVT U290 ( .A1(n33), .A2(fp_src2_in[23]), .A3(inq_din_d1[23]), .A4(
        n38), .A5(n37), .A6(inq_dout[23]), .Y(inq_in2[23]) );
  AO22X1_RVT U291 ( .A1(fp_op_in_7in), .A2(fp_srca_in[22]), .A3(n34), .A4(
        fp_srcb_in[22]), .Y(fp_src2_in[22]) );
  AO222X1_RVT U292 ( .A1(n33), .A2(fp_src2_in[22]), .A3(inq_din_d1[22]), .A4(
        n38), .A5(n37), .A6(inq_dout[22]), .Y(inq_in2[22]) );
  AO22X1_RVT U293 ( .A1(fp_op_in_7in), .A2(fp_srca_in[21]), .A3(n34), .A4(
        fp_srcb_in[21]), .Y(fp_src2_in[21]) );
  AO222X1_RVT U294 ( .A1(n33), .A2(fp_src2_in[21]), .A3(inq_din_d1[21]), .A4(
        n38), .A5(n37), .A6(inq_dout[21]), .Y(inq_in2[21]) );
  AO22X1_RVT U295 ( .A1(fp_op_in_7in), .A2(fp_srca_in[20]), .A3(n34), .A4(
        fp_srcb_in[20]), .Y(fp_src2_in[20]) );
  AO222X1_RVT U296 ( .A1(n33), .A2(fp_src2_in[20]), .A3(inq_din_d1[20]), .A4(
        n38), .A5(n37), .A6(inq_dout[20]), .Y(inq_in2[20]) );
  AO22X1_RVT U297 ( .A1(fp_op_in_7in), .A2(fp_srca_in[19]), .A3(n34), .A4(
        fp_srcb_in[19]), .Y(fp_src2_in[19]) );
  AO222X1_RVT U298 ( .A1(n33), .A2(fp_src2_in[19]), .A3(inq_din_d1[19]), .A4(
        n38), .A5(n37), .A6(inq_dout[19]), .Y(inq_in2[19]) );
  AO22X1_RVT U299 ( .A1(fp_op_in_7in), .A2(fp_srca_in[18]), .A3(n34), .A4(
        fp_srcb_in[18]), .Y(fp_src2_in[18]) );
  AO222X1_RVT U300 ( .A1(n33), .A2(fp_src2_in[18]), .A3(inq_din_d1[18]), .A4(
        n38), .A5(n37), .A6(inq_dout[18]), .Y(inq_in2[18]) );
  AO22X1_RVT U301 ( .A1(fp_op_in_7in), .A2(fp_srca_in[17]), .A3(n34), .A4(
        fp_srcb_in[17]), .Y(fp_src2_in[17]) );
  AO222X1_RVT U302 ( .A1(n33), .A2(fp_src2_in[17]), .A3(inq_din_d1[17]), .A4(
        n38), .A5(n37), .A6(inq_dout[17]), .Y(inq_in2[17]) );
  AO22X1_RVT U303 ( .A1(fp_op_in_7in), .A2(fp_srca_in[16]), .A3(n34), .A4(
        fp_srcb_in[16]), .Y(fp_src2_in[16]) );
  AO222X1_RVT U304 ( .A1(n33), .A2(fp_src2_in[16]), .A3(inq_din_d1[16]), .A4(
        n38), .A5(n37), .A6(inq_dout[16]), .Y(inq_in2[16]) );
  AO22X1_RVT U305 ( .A1(fp_op_in_7in), .A2(fp_srca_in[15]), .A3(n34), .A4(
        fp_srcb_in[15]), .Y(fp_src2_in[15]) );
  AO222X1_RVT U306 ( .A1(n33), .A2(fp_src2_in[15]), .A3(inq_din_d1[15]), .A4(
        n38), .A5(n37), .A6(inq_dout[15]), .Y(inq_in2[15]) );
  AO22X1_RVT U307 ( .A1(fp_op_in_7in), .A2(fp_srca_in[14]), .A3(n34), .A4(
        fp_srcb_in[14]), .Y(fp_src2_in[14]) );
  AO222X1_RVT U308 ( .A1(n33), .A2(fp_src2_in[14]), .A3(inq_din_d1[14]), .A4(
        n38), .A5(n37), .A6(inq_dout[14]), .Y(inq_in2[14]) );
  AO22X1_RVT U309 ( .A1(fp_op_in_7in), .A2(fp_srca_in[13]), .A3(n34), .A4(
        fp_srcb_in[13]), .Y(fp_src2_in[13]) );
  AO222X1_RVT U310 ( .A1(n33), .A2(fp_src2_in[13]), .A3(inq_din_d1[13]), .A4(
        n38), .A5(n37), .A6(inq_dout[13]), .Y(inq_in2[13]) );
  AO22X1_RVT U311 ( .A1(fp_op_in_7in), .A2(fp_srca_in[12]), .A3(n34), .A4(
        fp_srcb_in[12]), .Y(fp_src2_in[12]) );
  AO222X1_RVT U312 ( .A1(n33), .A2(fp_src2_in[12]), .A3(inq_din_d1[12]), .A4(
        n38), .A5(n37), .A6(inq_dout[12]), .Y(inq_in2[12]) );
  AO22X1_RVT U313 ( .A1(fp_op_in_7in), .A2(fp_srca_in[11]), .A3(n34), .A4(
        fp_srcb_in[11]), .Y(fp_src2_in[11]) );
  AO222X1_RVT U314 ( .A1(n33), .A2(fp_src2_in[11]), .A3(inq_din_d1[11]), .A4(
        n38), .A5(n37), .A6(inq_dout[11]), .Y(inq_in2[11]) );
  AO22X1_RVT U315 ( .A1(fp_op_in_7in), .A2(fp_srca_in[10]), .A3(n34), .A4(
        fp_srcb_in[10]), .Y(fp_src2_in[10]) );
  AO222X1_RVT U316 ( .A1(n33), .A2(fp_src2_in[10]), .A3(inq_din_d1[10]), .A4(
        n38), .A5(n37), .A6(inq_dout[10]), .Y(inq_in2[10]) );
  AO22X1_RVT U317 ( .A1(fp_op_in_7in), .A2(fp_srca_in[9]), .A3(n34), .A4(
        fp_srcb_in[9]), .Y(fp_src2_in[9]) );
  AO222X1_RVT U318 ( .A1(n33), .A2(fp_src2_in[9]), .A3(inq_din_d1[9]), .A4(n38), .A5(n37), .A6(inq_dout[9]), .Y(inq_in2[9]) );
  AO22X1_RVT U319 ( .A1(fp_op_in_7in), .A2(fp_srca_in[8]), .A3(n34), .A4(
        fp_srcb_in[8]), .Y(fp_src2_in[8]) );
  AO222X1_RVT U320 ( .A1(n33), .A2(fp_src2_in[8]), .A3(inq_din_d1[8]), .A4(n38), .A5(n37), .A6(inq_dout[8]), .Y(inq_in2[8]) );
  AO22X1_RVT U321 ( .A1(fp_op_in_7in), .A2(fp_srca_in[7]), .A3(n34), .A4(
        fp_srcb_in[7]), .Y(fp_src2_in[7]) );
  AO222X1_RVT U322 ( .A1(n33), .A2(fp_src2_in[7]), .A3(inq_din_d1[7]), .A4(n38), .A5(n37), .A6(inq_dout[7]), .Y(inq_in2[7]) );
  AO22X1_RVT U323 ( .A1(fp_op_in_7in), .A2(fp_srca_in[6]), .A3(n34), .A4(
        fp_srcb_in[6]), .Y(fp_src2_in[6]) );
  AO222X1_RVT U324 ( .A1(n33), .A2(fp_src2_in[6]), .A3(inq_din_d1[6]), .A4(n38), .A5(n37), .A6(inq_dout[6]), .Y(inq_in2[6]) );
  AO22X1_RVT U325 ( .A1(fp_op_in_7in), .A2(fp_srca_in[5]), .A3(n34), .A4(
        fp_srcb_in[5]), .Y(fp_src2_in[5]) );
  AO222X1_RVT U326 ( .A1(n33), .A2(fp_src2_in[5]), .A3(inq_din_d1[5]), .A4(n38), .A5(n37), .A6(inq_dout[5]), .Y(inq_in2[5]) );
  AO22X1_RVT U327 ( .A1(fp_op_in_7in), .A2(fp_srca_in[4]), .A3(n34), .A4(
        fp_srcb_in[4]), .Y(fp_src2_in[4]) );
  AO222X1_RVT U328 ( .A1(n33), .A2(fp_src2_in[4]), .A3(inq_din_d1[4]), .A4(n38), .A5(n37), .A6(inq_dout[4]), .Y(inq_in2[4]) );
  AO22X1_RVT U329 ( .A1(fp_op_in_7in), .A2(fp_srca_in[3]), .A3(n34), .A4(
        fp_srcb_in[3]), .Y(fp_src2_in[3]) );
  AO222X1_RVT U330 ( .A1(n33), .A2(fp_src2_in[3]), .A3(inq_din_d1[3]), .A4(n38), .A5(n37), .A6(inq_dout[3]), .Y(inq_in2[3]) );
  AO22X1_RVT U331 ( .A1(fp_op_in_7in), .A2(fp_srca_in[2]), .A3(n34), .A4(
        fp_srcb_in[2]), .Y(fp_src2_in[2]) );
  AO222X1_RVT U332 ( .A1(n33), .A2(fp_src2_in[2]), .A3(inq_din_d1[2]), .A4(n38), .A5(n37), .A6(inq_dout[2]), .Y(inq_in2[2]) );
  AO22X1_RVT U333 ( .A1(fp_op_in_7in), .A2(fp_srca_in[1]), .A3(n34), .A4(
        fp_srcb_in[1]), .Y(fp_src2_in[1]) );
  AO222X1_RVT U334 ( .A1(n33), .A2(fp_src2_in[1]), .A3(inq_din_d1[1]), .A4(n38), .A5(n37), .A6(inq_dout[1]), .Y(inq_in2[1]) );
  AO22X1_RVT U335 ( .A1(fp_op_in_7in), .A2(fp_srca_in[0]), .A3(n34), .A4(
        fp_srcb_in[0]), .Y(fp_src2_in[0]) );
  AO222X1_RVT U336 ( .A1(n33), .A2(fp_src2_in[0]), .A3(inq_din_d1[0]), .A4(n38), .A5(n37), .A6(inq_dout[0]), .Y(inq_in2[0]) );
endmodule


module fpu_in ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, a1stg_step, 
        m1stg_step, d1stg_step, add_pipe_active, mul_pipe_active, 
        div_pipe_active, inq_dout, sehold, arst_l, grst_l, rclk, fadd_clken_l, 
        fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div, inq_id, 
        inq_rnd_mode, inq_fcc, inq_op, inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, 
        inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1, 
        inq_in2_exp_neq_ffs, inq_in2_exp_eq_0, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2, fp_id_in, 
        fp_rnd_mode_in, fp_fcc_in, fp_op_in, fp_src1_in, fp_src2_in, 
        inq_rdaddr, inq_wraddr, inq_read_en, inq_we, se, si, so );
  input [123:0] pcx_fpio_data_px2;
  input [154:0] inq_dout;
  output [4:0] inq_id;
  output [1:0] inq_rnd_mode;
  output [1:0] inq_fcc;
  output [7:0] inq_op;
  output [63:0] inq_in1;
  output [63:0] inq_in2;
  output [4:0] fp_id_in;
  output [1:0] fp_rnd_mode_in;
  output [1:0] fp_fcc_in;
  output [7:0] fp_op_in;
  output [68:0] fp_src1_in;
  output [68:0] fp_src2_in;
  output [3:0] inq_rdaddr;
  output [3:0] inq_wraddr;
  input pcx_fpio_data_rdy_px2, a1stg_step, m1stg_step, d1stg_step,
         add_pipe_active, mul_pipe_active, div_pipe_active, sehold, arst_l,
         grst_l, rclk, se, si;
  output fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div,
         inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, inq_in1_53_0_neq_0,
         inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in2_exp_neq_ffs,
         inq_in2_exp_eq_0, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_read_en, inq_we, so;
  wire   pcx_fpio_data_px2_123, pcx_fpio_data_px2_122, pcx_fpio_data_px2_121,
         pcx_fpio_data_px2_120, pcx_fpio_data_px2_119, pcx_fpio_data_px2_118,
         pcx_fpio_data_px2_116, pcx_fpio_data_px2_115, pcx_fpio_data_px2_114,
         pcx_fpio_data_px2_113, pcx_fpio_data_px2_112, pcx_fpio_data_px2_79,
         pcx_fpio_data_px2_78, pcx_fpio_data_px2_77, pcx_fpio_data_px2_76,
         pcx_fpio_data_px2_75, pcx_fpio_data_px2_74, pcx_fpio_data_px2_73,
         pcx_fpio_data_px2_72, fp_op_in_7in, fp_data_rdy, inq_bp_inv,
         inq_fwrd_inv, net211165, net211166, net211167, net211168;
  assign pcx_fpio_data_px2_123 = pcx_fpio_data_px2[123];
  assign pcx_fpio_data_px2_122 = pcx_fpio_data_px2[122];
  assign pcx_fpio_data_px2_121 = pcx_fpio_data_px2[121];
  assign pcx_fpio_data_px2_120 = pcx_fpio_data_px2[120];
  assign pcx_fpio_data_px2_119 = pcx_fpio_data_px2[119];
  assign pcx_fpio_data_px2_118 = pcx_fpio_data_px2[118];
  assign pcx_fpio_data_px2_116 = pcx_fpio_data_px2[116];
  assign pcx_fpio_data_px2_115 = pcx_fpio_data_px2[115];
  assign pcx_fpio_data_px2_114 = pcx_fpio_data_px2[114];
  assign pcx_fpio_data_px2_113 = pcx_fpio_data_px2[113];
  assign pcx_fpio_data_px2_112 = pcx_fpio_data_px2[112];
  assign pcx_fpio_data_px2_79 = pcx_fpio_data_px2[79];
  assign pcx_fpio_data_px2_78 = pcx_fpio_data_px2[78];
  assign pcx_fpio_data_px2_77 = pcx_fpio_data_px2[77];
  assign pcx_fpio_data_px2_76 = pcx_fpio_data_px2[76];
  assign pcx_fpio_data_px2_75 = pcx_fpio_data_px2[75];
  assign pcx_fpio_data_px2_74 = pcx_fpio_data_px2[74];
  assign pcx_fpio_data_px2_73 = pcx_fpio_data_px2[73];
  assign pcx_fpio_data_px2_72 = pcx_fpio_data_px2[72];

  fpu_in_ctl fpu_in_ctl ( .pcx_fpio_data_rdy_px2(pcx_fpio_data_rdy_px2), 
        .pcx_fpio_data_px2({pcx_fpio_data_px2_123, pcx_fpio_data_px2_122, 
        pcx_fpio_data_px2_121, pcx_fpio_data_px2_120, pcx_fpio_data_px2_119, 
        pcx_fpio_data_px2_118}), .fp_op_in(fp_op_in[3:2]), .fp_op_in_7in(
        fp_op_in_7in), .a1stg_step(a1stg_step), .m1stg_step(m1stg_step), 
        .d1stg_step(d1stg_step), .add_pipe_active(add_pipe_active), 
        .mul_pipe_active(mul_pipe_active), .div_pipe_active(div_pipe_active), 
        .sehold(sehold), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), 
        .fp_data_rdy(fp_data_rdy), .fadd_clken_l(fadd_clken_l), .fmul_clken_l(
        fmul_clken_l), .fdiv_clken_l(fdiv_clken_l), .inq_we(inq_we), 
        .inq_wraddr(inq_wraddr), .inq_read_en(inq_read_en), .inq_rdaddr(
        inq_rdaddr), .inq_bp_inv(inq_bp_inv), .inq_fwrd_inv(inq_fwrd_inv), 
        .inq_add(inq_add), .inq_mul(inq_mul), .inq_div(inq_div), .se(se), .si(
        net211168) );
  fpu_in_dp fpu_in_dp ( .fp_data_rdy(fp_data_rdy), .fpio_data_px2_116_112({
        pcx_fpio_data_px2_116, pcx_fpio_data_px2_115, pcx_fpio_data_px2_114, 
        pcx_fpio_data_px2_113, pcx_fpio_data_px2_112}), .fpio_data_px2_79_72({
        pcx_fpio_data_px2_79, pcx_fpio_data_px2_78, pcx_fpio_data_px2_77, 
        pcx_fpio_data_px2_76, pcx_fpio_data_px2_75, pcx_fpio_data_px2_74, 
        pcx_fpio_data_px2_73, pcx_fpio_data_px2_72}), .fpio_data_px2_67_0(
        pcx_fpio_data_px2[67:0]), .inq_fwrd(net211165), .inq_fwrd_inv(
        inq_fwrd_inv), .inq_bp(net211166), .inq_bp_inv(inq_bp_inv), .inq_dout(
        inq_dout), .rclk(rclk), .fp_op_in_7in(fp_op_in_7in), .inq_id(inq_id), 
        .inq_rnd_mode(inq_rnd_mode), .inq_fcc(inq_fcc), .inq_op(inq_op), 
        .inq_in1_exp_neq_ffs(inq_in1_exp_neq_ffs), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(
        inq_in1_53_32_neq_0), .inq_in1(inq_in1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), 
        .inq_in2(inq_in2), .fp_id_in(fp_id_in), .fp_rnd_mode_in(fp_rnd_mode_in), .fp_fcc_in(fp_fcc_in), .fp_op_in(fp_op_in), .fp_src1_in(fp_src1_in), 
        .fp_src2_in(fp_src2_in), .se(se), .si(net211167) );
endmodule


module dffrl_async_SIZE1_4 ( din, clk, rst_l, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  wire   N4, n1;

  DFFARX1_RVT \q_reg[0]  ( .D(N4), .CLK(clk), .RSTB(rst_l), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
endmodule


module dffe_SIZE1_0 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n4, n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n4), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n4)
         );
endmodule


module dffe_SIZE1_141 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_140 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_139 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_138 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_137 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_136 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_135 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_134 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_133 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_132 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_131 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_130 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_129 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE8 ( din, rst, en, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input rst, en, clk, se;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, net24642, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE8 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24642), .TE(1'b0) );
  DFFX1_RVT \q_reg[7]  ( .D(N21), .CLK(net24642), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N20), .CLK(net24642), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N19), .CLK(net24642), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N18), .CLK(net24642), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N17), .CLK(net24642), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N16), .CLK(net24642), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N15), .CLK(net24642), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N14), .CLK(net24642), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N14) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N15) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N16) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N17) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N18) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N19) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[6]), .Y(N20) );
  AND2X1_RVT U12 ( .A1(n1), .A2(din[7]), .Y(N21) );
  NAND2X0_RVT U14 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dffe_SIZE1_128 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE4_0 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N4, net24462, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24462), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24462), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24462), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24462), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24462), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module dffe_SIZE1_127 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE4_4 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N4, net24462, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_4 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24462), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24462), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24462), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24462), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24462), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE2_0 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n6, n7, n1, n2, n3;

  DFFX1_RVT \q_reg[1]  ( .D(n7), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n6), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n7) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_0 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module dffe_SIZE2_21 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE31 ( din, rst, en, clk, q, se, si, so );
  input [30:0] din;
  output [30:0] q;
  input [30:0] si;
  output [30:0] so;
  input rst, en, clk, se;
  wire   N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, net24624, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE31 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24624), .TE(1'b0) );
  DFFX1_RVT \q_reg[30]  ( .D(N67), .CLK(net24624), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N66), .CLK(net24624), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N65), .CLK(net24624), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N64), .CLK(net24624), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N63), .CLK(net24624), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N62), .CLK(net24624), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N61), .CLK(net24624), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N60), .CLK(net24624), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N59), .CLK(net24624), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N58), .CLK(net24624), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N57), .CLK(net24624), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N56), .CLK(net24624), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N55), .CLK(net24624), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N54), .CLK(net24624), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N53), .CLK(net24624), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N52), .CLK(net24624), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N51), .CLK(net24624), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N50), .CLK(net24624), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N49), .CLK(net24624), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N48), .CLK(net24624), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N47), .CLK(net24624), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N46), .CLK(net24624), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N45), .CLK(net24624), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N44), .CLK(net24624), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N43), .CLK(net24624), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N42), .CLK(net24624), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N41), .CLK(net24624), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N40), .CLK(net24624), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N39), .CLK(net24624), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N38), .CLK(net24624), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N37), .CLK(net24624), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N37) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N38) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N39) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N40) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N41) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N42) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[6]), .Y(N43) );
  AND2X1_RVT U12 ( .A1(n1), .A2(din[7]), .Y(N44) );
  AND2X1_RVT U13 ( .A1(n1), .A2(din[8]), .Y(N45) );
  AND2X1_RVT U14 ( .A1(n1), .A2(din[9]), .Y(N46) );
  AND2X1_RVT U15 ( .A1(n1), .A2(din[10]), .Y(N47) );
  AND2X1_RVT U16 ( .A1(n1), .A2(din[11]), .Y(N48) );
  AND2X1_RVT U17 ( .A1(n1), .A2(din[12]), .Y(N49) );
  AND2X1_RVT U18 ( .A1(n1), .A2(din[13]), .Y(N50) );
  AND2X1_RVT U19 ( .A1(n1), .A2(din[14]), .Y(N51) );
  AND2X1_RVT U20 ( .A1(n1), .A2(din[15]), .Y(N52) );
  AND2X1_RVT U21 ( .A1(n1), .A2(din[16]), .Y(N53) );
  AND2X1_RVT U22 ( .A1(n1), .A2(din[17]), .Y(N54) );
  AND2X1_RVT U23 ( .A1(n1), .A2(din[18]), .Y(N55) );
  AND2X1_RVT U24 ( .A1(n1), .A2(din[19]), .Y(N56) );
  AND2X1_RVT U25 ( .A1(n1), .A2(din[20]), .Y(N57) );
  AND2X1_RVT U26 ( .A1(n1), .A2(din[21]), .Y(N58) );
  AND2X1_RVT U27 ( .A1(n1), .A2(din[22]), .Y(N59) );
  AND2X1_RVT U28 ( .A1(n1), .A2(din[23]), .Y(N60) );
  AND2X1_RVT U29 ( .A1(n1), .A2(din[24]), .Y(N61) );
  AND2X1_RVT U30 ( .A1(n1), .A2(din[25]), .Y(N62) );
  AND2X1_RVT U31 ( .A1(n1), .A2(din[26]), .Y(N63) );
  AND2X1_RVT U32 ( .A1(n1), .A2(din[27]), .Y(N64) );
  AND2X1_RVT U33 ( .A1(n1), .A2(din[28]), .Y(N65) );
  AND2X1_RVT U34 ( .A1(n1), .A2(din[29]), .Y(N66) );
  AND2X1_RVT U35 ( .A1(n1), .A2(din[30]), .Y(N67) );
  NAND2X0_RVT U37 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dffe_SIZE2_20 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_12 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_12 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE2_19 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE19 ( din, rst, en, clk, q, se, si, so );
  input [18:0] din;
  output [18:0] q;
  input [18:0] si;
  output [18:0] so;
  input rst, en, clk, se;
  wire   N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, net24606, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE19 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24606), .TE(1'b0) );
  DFFX1_RVT \q_reg[18]  ( .D(N43), .CLK(net24606), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N42), .CLK(net24606), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N41), .CLK(net24606), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N40), .CLK(net24606), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N39), .CLK(net24606), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N38), .CLK(net24606), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N37), .CLK(net24606), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N36), .CLK(net24606), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N35), .CLK(net24606), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N34), .CLK(net24606), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N33), .CLK(net24606), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N32), .CLK(net24606), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N31), .CLK(net24606), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N30), .CLK(net24606), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N29), .CLK(net24606), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N28), .CLK(net24606), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N27), .CLK(net24606), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N26), .CLK(net24606), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N25), .CLK(net24606), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N25) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N26) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N27) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N28) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N29) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N30) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[6]), .Y(N31) );
  AND2X1_RVT U12 ( .A1(n1), .A2(din[7]), .Y(N32) );
  AND2X1_RVT U13 ( .A1(n1), .A2(din[8]), .Y(N33) );
  AND2X1_RVT U14 ( .A1(n1), .A2(din[9]), .Y(N34) );
  AND2X1_RVT U15 ( .A1(n1), .A2(din[10]), .Y(N35) );
  AND2X1_RVT U16 ( .A1(n1), .A2(din[11]), .Y(N36) );
  AND2X1_RVT U17 ( .A1(n1), .A2(din[12]), .Y(N37) );
  AND2X1_RVT U18 ( .A1(n1), .A2(din[13]), .Y(N38) );
  AND2X1_RVT U19 ( .A1(n1), .A2(din[14]), .Y(N39) );
  AND2X1_RVT U20 ( .A1(n1), .A2(din[15]), .Y(N40) );
  AND2X1_RVT U21 ( .A1(n1), .A2(din[16]), .Y(N41) );
  AND2X1_RVT U22 ( .A1(n1), .A2(din[17]), .Y(N42) );
  AND2X1_RVT U23 ( .A1(n1), .A2(din[18]), .Y(N43) );
  NAND2X0_RVT U25 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dffre_SIZE2 ( din, rst, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input rst, en, clk, se;
  wire   n4, n5, n1, n2;

  DFFX1_RVT \q_reg[1]  ( .D(n5), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n4), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n4)
         );
  OA221X1_RVT U5 ( .A1(en), .A2(q[1]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE2_18 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_11 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_11 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE2_17 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE18 ( din, rst, en, clk, se, si, so, \q[17] , \q[16] , \q[15] , 
        \q[14] , \q[13] , \q[12] , \q[11] , \q[10]_BAR , \q[9] , \q[8] , 
        \q[7] , \q[6] , \q[5] , \q[4] , \q[3] , \q[2] , \q[1] , \q[0]  );
  input [17:0] din;
  input [17:0] si;
  output [17:0] so;
  input rst, en, clk, se;
  output \q[17] , \q[16] , \q[15] , \q[14] , \q[13] , \q[12] , \q[11] ,
         \q[10]_BAR , \q[9] , \q[8] , \q[7] , \q[6] , \q[5] , \q[4] , \q[3] ,
         \q[2] , \q[1] , \q[0] ;
  wire   N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, net24588, n4, n1, n2, n3;
  wire   [17:0] q;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE18 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24588), .TE(1'b0) );
  DFFX1_RVT \q_reg[17]  ( .D(N41), .CLK(net24588), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N40), .CLK(net24588), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N39), .CLK(net24588), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N38), .CLK(net24588), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N37), .CLK(net24588), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N36), .CLK(net24588), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N35), .CLK(net24588), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N34), .CLK(net24588), .QN(\q[10]_BAR ) );
  DFFX1_RVT \q_reg[9]  ( .D(N33), .CLK(net24588), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N32), .CLK(net24588), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N31), .CLK(net24588), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N30), .CLK(net24588), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N29), .CLK(net24588), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N28), .CLK(net24588), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N27), .CLK(net24588), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N26), .CLK(net24588), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N25), .CLK(net24588), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N24), .CLK(net24588), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N24) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N25) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N26) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N27) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N28) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N29) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[6]), .Y(N30) );
  AND2X1_RVT U12 ( .A1(n1), .A2(din[7]), .Y(N31) );
  AND2X1_RVT U13 ( .A1(n1), .A2(din[8]), .Y(N32) );
  AND2X1_RVT U14 ( .A1(n1), .A2(din[9]), .Y(N33) );
  AND2X1_RVT U15 ( .A1(n1), .A2(din[10]), .Y(N34) );
  AND2X1_RVT U16 ( .A1(n1), .A2(din[11]), .Y(N35) );
  AND2X1_RVT U17 ( .A1(n1), .A2(din[12]), .Y(N36) );
  AND2X1_RVT U18 ( .A1(n1), .A2(din[13]), .Y(N37) );
  AND2X1_RVT U19 ( .A1(n1), .A2(din[14]), .Y(N38) );
  AND2X1_RVT U20 ( .A1(n1), .A2(din[15]), .Y(N39) );
  AND2X1_RVT U21 ( .A1(n1), .A2(din[16]), .Y(N40) );
  AND2X1_RVT U22 ( .A1(n1), .A2(din[17]), .Y(N41) );
  NAND2X0_RVT U24 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dffe_SIZE2_16 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dffe_SIZE2_15 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE10_0 ( din, en, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, net24408, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24408), .TE(1'b0) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24408), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24408), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24408), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24408), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24408), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24408), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24408), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24408), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24408), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24408), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  OR2X1_RVT U14 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module dffe_SIZE2_14 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE9 ( din, rst, en, clk, q, se, si, so );
  input [8:0] din;
  output [8:0] q;
  input [8:0] si;
  output [8:0] so;
  input rst, en, clk, se;
  wire   N15, N16, N17, N18, N19, N20, N21, N22, N23, net24570, n4, n1, n2, n3
;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE9 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24570), .TE(1'b0) );
  DFFX1_RVT \q_reg[8]  ( .D(N23), .CLK(net24570), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N22), .CLK(net24570), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N21), .CLK(net24570), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N20), .CLK(net24570), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N19), .CLK(net24570), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N18), .CLK(net24570), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N17), .CLK(net24570), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N16), .CLK(net24570), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N15), .CLK(net24570), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N15) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N16) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N17) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N18) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N19) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N20) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[6]), .Y(N21) );
  AND2X1_RVT U12 ( .A1(n1), .A2(din[7]), .Y(N22) );
  AND2X1_RVT U13 ( .A1(n1), .A2(din[8]), .Y(N23) );
  NAND2X0_RVT U15 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE10_2 ( din, en, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, net24408, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_2 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24408), .TE(1'b0) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24408), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24408), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24408), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24408), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24408), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24408), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24408), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24408), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24408), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24408), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  OR2X1_RVT U14 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE6_0 ( din, rst, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input rst, en, clk, se;
  wire   N12, N13, N14, N15, N16, N17, net24282, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE6_0 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24282), .TE(1'b0) );
  DFFX1_RVT \q_reg[5]  ( .D(N17), .CLK(net24282), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N16), .CLK(net24282), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N15), .CLK(net24282), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N14), .CLK(net24282), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N13), .CLK(net24282), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N12), .CLK(net24282), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N12) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N13) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N14) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N15) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N16) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N17) );
  NAND2X0_RVT U12 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dff_SIZE10_0 ( din, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, n1;

  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
endmodule


module dffe_SIZE2_13 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dffre_SIZE1_10 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffe_SIZE1_126 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_125 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_124 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_123 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n2, n3, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n2) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n3), .A4(din[0]), .A5(n2), .Y(n5)
         );
endmodule


module dffe_SIZE1_122 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_121 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_120 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_119 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_118 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_117 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_116 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_115 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_114 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_113 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_112 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_111 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE2_12 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dffe_SIZE1_110 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_109 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE2_11 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dffe_SIZE1_108 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE2_10 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dffe_SIZE1_107 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_106 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_105 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_104 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_103 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_102 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_101 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_100 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_99 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_98 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_97 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_96 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_95 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_94 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_93 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_92 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_91 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_90 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_89 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_88 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module fpu_add_ctl ( inq_in1_51, inq_in1_54, inq_in1_63, inq_in1_50_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_51, 
        inq_in2_54, inq_in2_63, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_op, inq_rnd_mode, inq_id, 
        inq_fcc, inq_add, a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, 
        a1stg_in2_eq_in1_exp, a1stg_expadd1, a2stg_expadd, a2stg_frac2hi_neq_0, 
        a2stg_frac2lo_neq_0, a2stg_exp, a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, 
        a2stg_frac2_63, a4stg_exp, add_of_out_cout, a4stg_frac_neq_0, 
        a4stg_shl_data_neq_0, a4stg_frac_dbl_nx, a4stg_frac_sng_nx, 
        a1stg_expadd2, a1stg_expadd4_inv, a3stg_denorm, a3stg_denorm_inv, 
        a4stg_denorm_inv, a3stg_exp, a3stg_lead0, a4stg_rnd_frac_40, 
        a4stg_rnd_frac_39, a4stg_rnd_frac_11, a4stg_rnd_frac_10, 
        a4stg_frac_38_0_nx, a4stg_frac_9_0_nx, arst_l, grst_l, rclk, 
        add_pipe_active, a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1, 
        a1stg_denorm_sng_in2, a1stg_denorm_dbl_in2, a1stg_norm_sng_in1, 
        a1stg_norm_dbl_in1, a1stg_norm_sng_in2, a1stg_norm_dbl_in2, a1stg_step, 
        a1stg_stepa, a1stg_sngop, a1stg_intlngop, a1stg_fsdtoix, a1stg_fstod, 
        a1stg_fstoi, a1stg_fstox, a1stg_fdtoi, a1stg_fdtox, a1stg_faddsubs, 
        a1stg_faddsubd, a1stg_fdtos, a2stg_faddsubop, a2stg_fsdtoix_fdtos, 
        a2stg_fitos, a2stg_fitod, a2stg_fxtos, a2stg_fxtod, a3stg_faddsubop, 
        a3stg_faddsubopa, a4stg_dblop, a6stg_fadd_in, add_id_out_in, 
        add_fcc_out, a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, 
        a6stg_int_dst, a6stg_fcmpop, a6stg_step, a3stg_sub_in, add_sign_out, 
        add_cc_out, a4stg_in_of, add_exc_out, a2stg_frac1_in_frac1, 
        a2stg_frac1_in_frac2, a1stg_2nan_in_inv, a1stg_faddsubop_inv, 
        a2stg_frac1_in_qnan, a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, 
        a2stg_frac2_in_frac1, a2stg_frac2_in_qnan, a2stg_shr_cnt_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int, 
        a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max, 
        a2stg_sub_step, a2stg_fracadd_frac2_inv_in, 
        a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2, 
        a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add, 
        a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, 
        a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv, 
        a4stg_shl_cnt_in, a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0, 
        add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1, 
        add_exp_out_expadd, a4stg_to_0_inv, se, si, so, add_dest_rdy_BAR, 
        a4stg_round_BAR );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [1:0] inq_fcc;
  input [11:0] a1stg_expadd1;
  input [11:0] a2stg_expadd;
  input [11:0] a2stg_exp;
  input [11:0] a4stg_exp;
  input [5:0] a1stg_expadd2;
  input [10:0] a1stg_expadd4_inv;
  input [10:0] a3stg_exp;
  input [5:0] a3stg_lead0;
  output [1:0] a3stg_faddsubopa;
  output [9:0] add_id_out_in;
  output [1:0] add_fcc_out;
  output [1:0] add_cc_out;
  output [4:0] add_exc_out;
  output [5:0] a2stg_shr_cnt_in;
  output [9:0] a4stg_shl_cnt_in;
  input inq_in1_51, inq_in1_54, inq_in1_63, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_63, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add,
         a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, a1stg_in2_eq_in1_exp,
         a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0, a3stg_fsdtoix_nx,
         a3stg_fsdtoi_nx, a2stg_frac2_63, add_of_out_cout, a4stg_frac_neq_0,
         a4stg_shl_data_neq_0, a4stg_frac_dbl_nx, a4stg_frac_sng_nx,
         a3stg_denorm, a3stg_denorm_inv, a4stg_denorm_inv, a4stg_rnd_frac_40,
         a4stg_rnd_frac_39, a4stg_rnd_frac_11, a4stg_rnd_frac_10,
         a4stg_frac_38_0_nx, a4stg_frac_9_0_nx, arst_l, grst_l, rclk, se, si,
         add_dest_rdy_BAR, a4stg_round_BAR;
  output add_pipe_active, a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1,
         a1stg_denorm_sng_in2, a1stg_denorm_dbl_in2, a1stg_norm_sng_in1,
         a1stg_norm_dbl_in1, a1stg_norm_sng_in2, a1stg_norm_dbl_in2,
         a1stg_step, a1stg_stepa, a1stg_sngop, a1stg_intlngop, a1stg_fsdtoix,
         a1stg_fstod, a1stg_fstoi, a1stg_fstox, a1stg_fdtoi, a1stg_fdtox,
         a1stg_faddsubs, a1stg_faddsubd, a1stg_fdtos, a2stg_faddsubop,
         a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod, a2stg_fxtos,
         a2stg_fxtod, a3stg_faddsubop, a4stg_dblop, a6stg_fadd_in,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         a6stg_fcmpop, a6stg_step, a3stg_sub_in, add_sign_out, a4stg_in_of,
         a2stg_frac1_in_frac1, a2stg_frac1_in_frac2, a1stg_2nan_in_inv,
         a1stg_faddsubop_inv, a2stg_frac1_in_qnan, a2stg_frac1_in_nv,
         a2stg_frac1_in_nv_dbl, a2stg_frac2_in_frac1, a2stg_frac2_in_qnan,
         a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add,
         a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0,
         a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1,
         add_exp_out_expadd, a4stg_to_0_inv, so;
  wire   add_dest_rdy, a4stg_round, add_exc_out_0, add_exp_out_expinc,
         add_exp_out_expadd, add_ctl_rst_l, a1stg_in1_51, a1stg_in1_54,
         a1stg_in1_63, a1stg_in1_50_0_neq_0, a1stg_in1_53_32_neq_0,
         a1stg_in1_exp_eq_0, a1stg_in1_exp_neq_ffs, a1stg_in2_51, a1stg_in2_54,
         a1stg_in2_63, a1stg_in2_50_0_neq_0, a1stg_in2_53_32_neq_0,
         a1stg_in2_exp_eq_0, a1stg_in2_exp_neq_ffs, a1stg_snan_in1,
         a1stg_snan_in2, a1stg_qnan_in1, a1stg_qnan_in2, a1stg_nan_in2,
         a1stg_nan_in, a1stg_2inf_in, a1stg_2zero_in, a1stg_dblop,
         a2stg_opdec_36, a2stg_opdec_28, a3stg_opdec_36, a3stg_opdec_24,
         a3stg_fsdtoix, a4stg_faddsub_dtosop, a4stg_fsdtoix, a4stg_fcmpop,
         a5stg_opdec_9, a5stg_fixtos_fxtod, a5stg_fixtos, a5stg_fxtod,
         a6stg_opdec_in_9, \a6stg_opdec[34] , add_pipe_active_in, a1stg_sub,
         a2stg_sign1, a2stg_sign2, a2stg_sub, a2stg_in2_neq_in1_frac,
         a2stg_in2_gt_in1_frac, a2stg_in2_eq_in1_exp, a2stg_in2_gt_in1_exp,
         a2stg_nan_in, a2stg_nan_in2, a2stg_snan_in2, a2stg_qnan_in2,
         a2stg_snan_in1, a2stg_qnan_in1, a2stg_2zero_in, a2stg_2inf_in,
         a3stg_sign_in, a3stg_sign, a4stg_sign2, a4stg_sign_in, a4stg_sign,
         a1stg_nv, a2stg_nv, a2stg_of_mask, a3stg_nv_in, a3stg_nv,
         a3stg_of_mask, a2stg_nx_tmp1, a2stg_nx_tmp2, a2stg_nx_tmp3,
         a3stg_a2_expadd_11, a3stg_nx_tmp1, a3stg_nx_tmp2, a3stg_nx_tmp3,
         a3stg_nx, a4stg_nv2, a4stg_nv_in, a4stg_nv, a4stg_of_mask2,
         a4stg_of_mask_in, a4stg_of_mask, a4stg_nx2, a4stg_nx_in, a4stg_nx,
         add_of_out_tmp1_in, add_of_out_tmp1, add_of_out_tmp2, a4stg_uf,
         add_nx_out_in, add_nx_out, a2stg_fracadd_frac2_in, N27, N1616, n242,
         n244, n256, n257, n258, n259, n260, n261, n262, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n243, n245, n246, n247, n248,
         n249, a1stg_stepa;
  wire   [3:0] a1stg_sngopa;
  wire   [3:0] a1stg_dblopa;
  wire   [7:0] a1stg_op_in;
  wire   [7:0] a1stg_op;
  wire   [1:0] a1stg_rnd_mode;
  wire   [4:0] a1stg_id;
  wire   [1:0] a1stg_fcc;
  wire   [30:0] a2stg_opdec_in;
  wire   [34:30] a2stg_opdec;
  wire   [3:0] a2stg_opdec_24_21;
  wire   [8:4] a2stg_opdec_19_11;
  wire   [9:1] a2stg_opdec_9_0;
  wire   [1:0] a2stg_rnd_mode;
  wire   [4:0] a2stg_id;
  wire   [1:0] a2stg_fcc;
  wire   [34:30] a3stg_opdec;
  wire   [9:0] a3stg_opdec_9_0;
  wire   [1:0] a3stg_rnd_mode;
  wire   [4:0] a3stg_id;
  wire   [1:0] a3stg_fcc;
  wire   [34:29] a4stg_opdec;
  wire   [7:0] a4stg_opdec_7_0;
  wire   [1:0] a4stg_rnd_mode2;
  wire   [1:0] a4stg_rnd_mode_in;
  wire   [1:0] a4stg_rnd_mode;
  wire   [9:0] a4stg_id;
  wire   [1:0] a4stg_fcc;
  wire   [34:30] a5stg_opdec;
  wire   [9:0] a5stg_id;
  wire   [34:30] a6stg_opdec_in;
  wire   [9:0] add_id_out;
  wire   [1:0] add_fcc_out_in;
  wire   [1:0] a2stg_cc;
  wire   [1:0] a3stg_cc;
  wire   [1:0] a4stg_cc;
  wire   [1:0] add_cc_out_in;
  assign add_dest_rdy = add_dest_rdy_BAR;
  assign a4stg_round = a4stg_round_BAR;
  assign add_exc_out[0] = add_exc_out_0;
  assign add_frac_out_rndadd = add_exp_out_expinc;
  assign add_frac_out_shl = add_exp_out_expadd;
  assign a4stg_to_0_inv = N1616;
  assign add_exc_out[1] = 1'b0;
  assign so = 1'b0;
  assign a1stg_step = a1stg_stepa;

  dffrl_async_SIZE1_4 dffrl_add_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(add_ctl_rst_l), .se(se), .si(1'b0) );
  dffe_SIZE1_0 i_a1stg_in1_51 ( .din(inq_in1_51), .en(a1stg_stepa), .clk(rclk), 
        .q(a1stg_in1_51), .se(se), .si(1'b0) );
  dffe_SIZE1_141 i_a1stg_in1_54 ( .din(inq_in1_54), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_in1_54), .se(se), .si(1'b0) );
  dffe_SIZE1_140 i_a1stg_in1_63 ( .din(inq_in1_63), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_in1_63), .se(se), .si(1'b0) );
  dffe_SIZE1_139 i_a1stg_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in1_50_0_neq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_138 i_a1stg_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in1_53_32_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_137 i_a1stg_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in1_exp_eq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_136 i_a1stg_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in1_exp_neq_ffs), .se(se), .si(1'b0) );
  dffe_SIZE1_135 i_a1stg_in2_51 ( .din(inq_in2_51), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_in2_51), .se(se), .si(1'b0) );
  dffe_SIZE1_134 i_a1stg_in2_54 ( .din(inq_in2_54), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_in2_54), .se(se), .si(1'b0) );
  dffe_SIZE1_133 i_a1stg_in2_63 ( .din(inq_in2_63), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_in2_63), .se(se), .si(1'b0) );
  dffe_SIZE1_132 i_a1stg_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in2_50_0_neq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_131 i_a1stg_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in2_53_32_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_130 i_a1stg_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in2_exp_eq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_129 i_a1stg_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_in2_exp_neq_ffs), .se(se), .si(1'b0) );
  dffre_SIZE8 i_a1stg_op ( .din(a1stg_op_in), .rst(n242), .en(a1stg_stepa), 
        .clk(rclk), .q(a1stg_op), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE1_128 i_a1stg_sngop ( .din(inq_op[0]), .en(a1stg_stepa), .clk(rclk), 
        .q(a1stg_sngop), .se(se), .si(1'b0) );
  dffe_SIZE4_0 i_a1stg_sngopa ( .din({1'b0, 1'b0, 1'b0, inq_op[0]}), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_sngopa), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dffe_SIZE1_127 i_a1stg_dblop ( .din(inq_op[1]), .en(a1stg_stepa), .clk(rclk), 
        .q(a1stg_dblop), .se(se), .si(1'b0) );
  dffe_SIZE4_4 i_a1stg_dblopa ( .din({1'b0, 1'b0, 1'b0, inq_op[1]}), .en(
        a1stg_stepa), .clk(rclk), .q(a1stg_dblopa), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dffe_SIZE2_0 i_a1stg_rnd_mode ( .din(inq_rnd_mode), .en(a1stg_stepa), .clk(
        rclk), .q(a1stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_0 i_a1stg_id ( .din(inq_id), .en(a1stg_stepa), .clk(rclk), .q(
        a1stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_21 i_a1stg_fcc ( .din(inq_fcc), .en(a1stg_stepa), .clk(rclk), .q(
        a1stg_fcc), .se(se), .si({1'b0, 1'b0}) );
  dffre_SIZE31 i_a2stg_opdec ( .din(a2stg_opdec_in), .rst(n242), .en(
        a6stg_step), .clk(rclk), .q({a2stg_opdec_36, a2stg_opdec, 
        a2stg_faddsubop, a2stg_opdec_28, a2stg_opdec_24_21, a2stg_opdec_19_11, 
        a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod, a2stg_fxtos, 
        a2stg_opdec_9_0, a2stg_fxtod}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_20 i_a2stg_rnd_mode ( .din(a1stg_rnd_mode), .en(a6stg_step), 
        .clk(rclk), .q(a2stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_12 i_a2stg_id ( .din(a1stg_id), .en(a6stg_step), .clk(rclk), .q(
        a2stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_19 i_a2stg_fcc ( .din(a1stg_fcc), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_fcc), .se(se), .si({1'b0, 1'b0}) );
  dffre_SIZE19 i_a3stg_opdec ( .din({a2stg_opdec_36, a2stg_opdec, 
        a2stg_faddsubop, a2stg_opdec_24_21[3], a2stg_opdec_24_21[0], 
        a2stg_opdec_9_0, a2stg_fxtod}), .rst(n242), .en(a6stg_step), .clk(rclk), .q({a3stg_opdec_36, a3stg_opdec, a3stg_faddsubop, a3stg_opdec_24, 
        a3stg_fsdtoix, a3stg_opdec_9_0}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffre_SIZE2 i_a3stg_faddsubopa ( .din({1'b0, a2stg_faddsubop}), .rst(n242), 
        .en(a6stg_step), .clk(rclk), .q(a3stg_faddsubopa), .se(se), .si({1'b0, 
        1'b0}) );
  dffe_SIZE2_18 i_a3stg_rnd_mode ( .din(a2stg_rnd_mode), .en(a6stg_step), 
        .clk(rclk), .q(a3stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_11 i_a3stg_id ( .din(a2stg_id), .en(a6stg_step), .clk(rclk), .q(
        a3stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_17 i_a3stg_fcc ( .din(a2stg_fcc), .en(a6stg_step), .clk(rclk), 
        .q(a3stg_fcc), .se(se), .si({1'b0, 1'b0}) );
  dffre_SIZE18 i_a4stg_opdec ( .din({a3stg_opdec_36, a3stg_opdec, 
        a3stg_faddsubop, a3stg_opdec_24, a3stg_fsdtoix, a3stg_opdec_9_0[9], 
        a3stg_opdec_9_0[7:0]}), .rst(n242), .en(a6stg_step), .clk(rclk), .se(
        se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\q[17] (a4stg_dblop), .\q[16] (a4stg_opdec[34]), .\q[15] (a4stg_opdec[33]), .\q[14] (
        a4stg_opdec[32]), .\q[13] (a4stg_opdec[31]), .\q[12] (a4stg_opdec[30]), 
        .\q[11] (a4stg_opdec[29]), .\q[10]_BAR (a4stg_faddsub_dtosop), 
        .\q[9] (a4stg_fsdtoix), .\q[8] (a4stg_fcmpop), .\q[7] (
        a4stg_opdec_7_0[7]), .\q[6] (a4stg_opdec_7_0[6]), .\q[5] (
        a4stg_opdec_7_0[5]), .\q[4] (a4stg_opdec_7_0[4]), .\q[3] (
        a4stg_opdec_7_0[3]), .\q[2] (a4stg_opdec_7_0[2]), .\q[1] (
        a4stg_opdec_7_0[1]), .\q[0] (a4stg_opdec_7_0[0]) );
  dffe_SIZE2_16 i_a4stg_rnd_mode ( .din(a4stg_rnd_mode_in), .en(a6stg_step), 
        .clk(rclk), .q(a4stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE2_15 i_a4stg_rnd_mode2 ( .din(a3stg_rnd_mode), .en(a6stg_step), 
        .clk(rclk), .q(a4stg_rnd_mode2), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE10_0 i_a4stg_id ( .din({N27, n262, n256, n261, n257, n260, n258, 
        n259, a3stg_id[1:0]}), .en(a6stg_step), .clk(rclk), .q(a4stg_id), .se(
        se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0})
         );
  dffe_SIZE2_14 i_a4stg_fcc ( .din(a3stg_fcc), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_fcc), .se(se), .si({1'b0, 1'b0}) );
  dffre_SIZE9 i_a5stg_opdec ( .din({a4stg_opdec[34:30], a4stg_fcmpop, 
        a4stg_opdec_7_0[7], a4stg_opdec_7_0[1:0]}), .rst(n242), .en(a6stg_step), .clk(rclk), .q({a5stg_opdec, a5stg_opdec_9, a5stg_fixtos_fxtod, a5stg_fixtos, 
        a5stg_fxtod}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dffe_SIZE10_2 i_a5stg_id ( .din(a4stg_id), .en(a6stg_step), .clk(rclk), .q(
        a5stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffre_SIZE6_0 i_a6stg_opdec ( .din({a6stg_opdec_in, a6stg_opdec_in_9}), 
        .rst(n242), .en(a6stg_step), .clk(rclk), .q({\a6stg_opdec[34] , 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        a6stg_fcmpop}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE10_0 i_add_id_out ( .din(add_id_out_in), .clk(rclk), .q(add_id_out), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE2_13 i_add_fcc_out ( .din(add_fcc_out_in), .en(a6stg_step), .clk(
        rclk), .q(add_fcc_out), .se(se), .si({1'b0, 1'b0}) );
  dffre_SIZE1_10 i_add_pipe_active ( .din(add_pipe_active_in), .rst(n242), 
        .en(1'b1), .clk(rclk), .q(add_pipe_active), .se(se), .si(1'b0) );
  dffe_SIZE1_126 i_a2stg_sign1 ( .din(a1stg_in1_63), .en(a6stg_step), .clk(
        rclk), .q(a2stg_sign1), .se(se), .si(1'b0) );
  dffe_SIZE1_125 i_a2stg_sign2 ( .din(a1stg_in2_63), .en(a6stg_step), .clk(
        rclk), .q(a2stg_sign2), .se(se), .si(1'b0) );
  dffe_SIZE1_124 i_a2stg_sub ( .din(a1stg_sub), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_sub), .se(se), .si(1'b0) );
  dffe_SIZE1_123 i_a2stg_in2_neq_in1_frac ( .din(a1stg_in2_neq_in1_frac), .en(
        a6stg_step), .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (
        a2stg_in2_neq_in1_frac) );
  dffe_SIZE1_122 i_a2stg_in2_gt_in1_frac ( .din(a1stg_in2_gt_in1_frac), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_gt_in1_frac), .se(se), .si(1'b0)
         );
  dffe_SIZE1_121 i_a2stg_in2_eq_in1_exp ( .din(a1stg_in2_eq_in1_exp), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_eq_in1_exp), .se(se), .si(1'b0)
         );
  dffe_SIZE1_120 i_a2stg_in2_gt_in1_exp ( .din(a1stg_expadd1[11]), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_gt_in1_exp), .se(se), .si(1'b0)
         );
  dffe_SIZE1_119 i_a2stg_nan_in ( .din(a1stg_nan_in), .en(a6stg_step), .clk(
        rclk), .q(a2stg_nan_in), .se(se), .si(1'b0) );
  dffe_SIZE1_118 i_a2stg_nan_in2 ( .din(a1stg_nan_in2), .en(a6stg_step), .clk(
        rclk), .q(a2stg_nan_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_117 i_a2stg_snan_in2 ( .din(a1stg_snan_in2), .en(a6stg_step), 
        .clk(rclk), .q(a2stg_snan_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_116 i_a2stg_qnan_in2 ( .din(a1stg_qnan_in2), .en(a6stg_step), 
        .clk(rclk), .q(a2stg_qnan_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_115 i_a2stg_snan_in1 ( .din(a1stg_snan_in1), .en(a6stg_step), 
        .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (a2stg_snan_in1) );
  dffe_SIZE1_114 i_a2stg_qnan_in1 ( .din(a1stg_qnan_in1), .en(a6stg_step), 
        .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (a2stg_qnan_in1) );
  dffe_SIZE1_113 i_a2stg_2zero_in ( .din(a1stg_2zero_in), .en(a6stg_step), 
        .clk(rclk), .q(a2stg_2zero_in), .se(se), .si(1'b0) );
  dffe_SIZE1_112 i_a2stg_2inf_in ( .din(a1stg_2inf_in), .en(a6stg_step), .clk(
        rclk), .q(a2stg_2inf_in), .se(se), .si(1'b0) );
  dffe_SIZE1_111 i_a3stg_sign ( .din(a3stg_sign_in), .en(a6stg_step), .clk(
        rclk), .q(a3stg_sign), .se(se), .si(1'b0) );
  dffe_SIZE2_12 i_a3stg_cc ( .din(a2stg_cc), .en(a6stg_step), .clk(rclk), .q(
        a3stg_cc), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE1_110 i_a4stg_sign ( .din(a4stg_sign_in), .en(a6stg_step), .clk(
        rclk), .q(a4stg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_109 i_a4stg_sign2 ( .din(a3stg_sign), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_sign2), .se(se), .si(1'b0) );
  dffe_SIZE2_11 i_a4stg_cc ( .din(a3stg_cc), .en(a6stg_step), .clk(rclk), .q(
        a4stg_cc), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE1_108 i_add_sign_out ( .din(a4stg_sign), .en(a6stg_step), .clk(rclk), .q(add_sign_out), .se(se), .si(1'b0) );
  dffe_SIZE2_10 i_add_cc_out ( .din(add_cc_out_in), .en(a6stg_step), .clk(rclk), .q(add_cc_out), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE1_107 i_a2stg_nv ( .din(a1stg_nv), .en(a6stg_step), .clk(rclk), .q(
        a2stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_106 i_a2stg_of_mask ( .din(n244), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_105 i_a3stg_nv ( .din(a3stg_nv_in), .en(a6stg_step), .clk(rclk), 
        .q(a3stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_104 i_a3stg_of_mask ( .din(a2stg_of_mask), .en(a6stg_step), .clk(
        rclk), .q(a3stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_103 i_a3stg_a2_expadd_11 ( .din(a2stg_expadd[11]), .en(a6stg_step), .clk(rclk), .q(a3stg_a2_expadd_11), .se(se), .si(1'b0) );
  dffe_SIZE1_102 i_a3stg_nx_tmp1 ( .din(a2stg_nx_tmp1), .en(a6stg_step), .clk(
        rclk), .q(a3stg_nx_tmp1), .se(se), .si(1'b0) );
  dffe_SIZE1_101 i_a3stg_nx_tmp2 ( .din(a2stg_nx_tmp2), .en(a6stg_step), .clk(
        rclk), .q(a3stg_nx_tmp2), .se(se), .si(1'b0) );
  dffe_SIZE1_100 i_a3stg_nx_tmp3 ( .din(a2stg_nx_tmp3), .en(a6stg_step), .clk(
        rclk), .q(a3stg_nx_tmp3), .se(se), .si(1'b0) );
  dffe_SIZE1_99 i_a4stg_nv ( .din(a4stg_nv_in), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_98 i_a4stg_nv2 ( .din(a3stg_nv), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nv2), .se(se), .si(1'b0) );
  dffe_SIZE1_97 i_a4stg_of_mask ( .din(a4stg_of_mask_in), .en(a6stg_step), 
        .clk(rclk), .q(a4stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_96 i_a4stg_of_mask2 ( .din(a3stg_of_mask), .en(a6stg_step), .clk(
        rclk), .q(a4stg_of_mask2), .se(se), .si(1'b0) );
  dffe_SIZE1_95 i_a4stg_nx ( .din(a4stg_nx_in), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_nx), .se(se), .si(1'b0) );
  dffe_SIZE1_94 i_a4stg_nx2 ( .din(a3stg_nx), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nx2), .se(se), .si(1'b0) );
  dffe_SIZE1_93 i_add_nv_out ( .din(a4stg_nv), .en(a6stg_step), .clk(rclk), 
        .q(add_exc_out[4]), .se(se), .si(1'b0) );
  dffe_SIZE1_92 i_add_of_out_tmp1 ( .din(add_of_out_tmp1_in), .en(a6stg_step), 
        .clk(rclk), .q(add_of_out_tmp1), .se(se), .si(1'b0) );
  dffe_SIZE1_91 i_add_of_out_tmp2 ( .din(a4stg_in_of), .en(a6stg_step), .clk(
        rclk), .q(add_of_out_tmp2), .se(se), .si(1'b0) );
  dffe_SIZE1_90 i_add_uf_out ( .din(a4stg_uf), .en(a6stg_step), .clk(rclk), 
        .q(add_exc_out[2]), .se(se), .si(1'b0) );
  dffe_SIZE1_89 i_add_nx_out ( .din(add_nx_out_in), .en(a6stg_step), .clk(rclk), .q(add_nx_out), .se(se), .si(1'b0) );
  dffe_SIZE1_88 i_a2stg_fracadd_frac2 ( .din(a2stg_fracadd_frac2_in), .en(
        a6stg_step), .clk(rclk), .q(a2stg_fracadd_frac2), .se(se), .si(1'b0)
         );
  INVX0_RVT U3 ( .A(n202), .Y(n203) );
  OR3X1_RVT U4 ( .A1(a1stg_expadd1[11]), .A2(a1stg_expadd1[0]), .A3(n198), .Y(
        n201) );
  OR3X1_RVT U5 ( .A1(a1stg_expadd1[8]), .A2(a1stg_expadd1[7]), .A3(n177), .Y(
        n198) );
  OR3X1_RVT U6 ( .A1(a1stg_expadd1[9]), .A2(a1stg_expadd1[6]), .A3(
        a1stg_expadd1[10]), .Y(n177) );
  INVX0_RVT U7 ( .A(a1stg_expadd1[11]), .Y(n178) );
  INVX0_RVT U8 ( .A(a2stg_expadd[11]), .Y(n96) );
  INVX0_RVT U9 ( .A(n222), .Y(n218) );
  INVX0_RVT U10 ( .A(n224), .Y(n219) );
  INVX0_RVT U11 ( .A(a2stg_expadd[9]), .Y(n124) );
  INVX0_RVT U12 ( .A(a3stg_denorm), .Y(n225) );
  INVX0_RVT U13 ( .A(a2stg_expadd[7]), .Y(n123) );
  INVX0_RVT U14 ( .A(n213), .Y(n211) );
  INVX0_RVT U15 ( .A(n208), .Y(n204) );
  INVX0_RVT U16 ( .A(n87), .Y(a2stg_opdec_in[5]) );
  INVX0_RVT U17 ( .A(n194), .Y(n133) );
  OR3X1_RVT U18 ( .A1(a4stg_exp[8]), .A2(a4stg_exp[9]), .A3(a4stg_exp[10]), 
        .Y(n18) );
  INVX0_RVT U19 ( .A(a4stg_exp[1]), .Y(n160) );
  INVX0_RVT U20 ( .A(a4stg_exp[7]), .Y(n159) );
  INVX0_RVT U21 ( .A(n67), .Y(n86) );
  OR3X1_RVT U22 ( .A1(a2stg_exp[9]), .A2(a2stg_exp[7]), .A3(a2stg_exp[8]), .Y(
        n142) );
  INVX0_RVT U23 ( .A(a2stg_exp[5]), .Y(n138) );
  INVX0_RVT U24 ( .A(a2stg_exp[6]), .Y(n139) );
  INVX0_RVT U25 ( .A(a3stg_exp[2]), .Y(n235) );
  INVX0_RVT U26 ( .A(a3stg_exp[1]), .Y(n236) );
  INVX0_RVT U27 ( .A(n73), .Y(n78) );
  INVX0_RVT U28 ( .A(n7), .Y(n80) );
  INVX0_RVT U29 ( .A(n43), .Y(n77) );
  INVX0_RVT U30 ( .A(n68), .Y(n70) );
  INVX0_RVT U31 ( .A(n172), .Y(a1stg_snan_in1) );
  INVX0_RVT U32 ( .A(n35), .Y(n58) );
  INVX1_RVT U33 ( .A(\a6stg_opdec[34] ), .Y(n94) );
  INVX0_RVT U34 ( .A(a4stg_opdec_7_0[6]), .Y(n22) );
  INVX0_RVT U35 ( .A(a2stg_opdec_19_11[5]), .Y(n141) );
  INVX0_RVT U36 ( .A(n115), .Y(n98) );
  INVX0_RVT U37 ( .A(a2stg_opdec_28), .Y(n102) );
  INVX0_RVT U38 ( .A(a1stg_op[3]), .Y(n4) );
  INVX0_RVT U39 ( .A(a4stg_opdec_7_0[3]), .Y(n157) );
  INVX0_RVT U40 ( .A(n33), .Y(n54) );
  INVX0_RVT U41 ( .A(n34), .Y(n56) );
  INVX0_RVT U42 ( .A(n32), .Y(n55) );
  INVX1_RVT U43 ( .A(a2stg_sub), .Y(n114) );
  INVX0_RVT U44 ( .A(a2stg_2inf_in), .Y(n97) );
  INVX0_RVT U45 ( .A(a2stg_nan_in), .Y(n107) );
  INVX0_RVT U46 ( .A(a2stg_snan_in2), .Y(n110) );
  INVX0_RVT U47 ( .A(a4stg_rnd_mode[0]), .Y(n12) );
  INVX0_RVT U48 ( .A(a1stg_in1_51), .Y(n40) );
  INVX0_RVT U49 ( .A(a4stg_sign), .Y(n13) );
  INVX0_RVT U50 ( .A(a1stg_in1_54), .Y(n39) );
  INVX0_RVT U51 ( .A(a1stg_in2_51), .Y(n9) );
  INVX0_RVT U52 ( .A(a1stg_in2_54), .Y(n8) );
  AND2X1_RVT U53 ( .A1(a2stg_sub), .A2(a6stg_step), .Y(a2stg_sub_step) );
  AND2X1_RVT U54 ( .A1(n3), .A2(a6stg_step), .Y(a1stg_stepa) );
  AND2X1_RVT U55 ( .A1(\a6stg_opdec[34] ), .A2(add_dest_rdy), .Y(n92) );
  INVX1_RVT U56 ( .A(n92), .Y(a6stg_step) );
  INVX1_RVT U57 ( .A(a1stg_op[1]), .Y(n44) );
  INVX1_RVT U58 ( .A(a1stg_op[0]), .Y(n82) );
  INVX1_RVT U59 ( .A(a1stg_op[2]), .Y(n60) );
  NAND2X0_RVT U60 ( .A1(a1stg_op[6]), .A2(n60), .Y(n1) );
  NAND4X0_RVT U61 ( .A1(a1stg_op[7]), .A2(n44), .A3(n82), .A4(n1), .Y(n2) );
  NAND2X0_RVT U62 ( .A1(a2stg_opdec_9_0[7]), .A2(n2), .Y(n3) );
  INVX1_RVT U63 ( .A(a1stg_in1_exp_eq_0), .Y(n5) );
  AND2X1_RVT U64 ( .A1(a1stg_dblopa[0]), .A2(n5), .Y(a1stg_norm_dbl_in1) );
  INVX1_RVT U65 ( .A(a1stg_in2_exp_eq_0), .Y(n6) );
  AND2X1_RVT U66 ( .A1(a1stg_dblopa[0]), .A2(n6), .Y(a1stg_norm_dbl_in2) );
  NOR2X0_RVT U67 ( .A1(a1stg_sngopa[3]), .A2(a1stg_dblop), .Y(a1stg_intlngop)
         );
  AND2X1_RVT U68 ( .A1(a1stg_in2_exp_eq_0), .A2(a1stg_dblopa[0]), .Y(
        a1stg_denorm_dbl_in2) );
  AND2X1_RVT U69 ( .A1(a1stg_in1_exp_eq_0), .A2(a1stg_dblopa[0]), .Y(
        a1stg_denorm_dbl_in1) );
  NAND2X0_RVT U70 ( .A1(a1stg_op[0]), .A2(n44), .Y(n43) );
  NAND2X0_RVT U71 ( .A1(a1stg_op[1]), .A2(n82), .Y(n7) );
  NAND2X0_RVT U72 ( .A1(n43), .A2(n7), .Y(n74) );
  INVX1_RVT U73 ( .A(a1stg_op[7]), .Y(n48) );
  NOR3X0_RVT U74 ( .A1(a1stg_op[5]), .A2(a1stg_op[2]), .A3(n48), .Y(n45) );
  INVX1_RVT U75 ( .A(a1stg_op[6]), .Y(n85) );
  INVX1_RVT U76 ( .A(a1stg_op[4]), .Y(n46) );
  NAND4X0_RVT U77 ( .A1(n45), .A2(n4), .A3(n85), .A4(n46), .Y(n61) );
  NAND4X0_RVT U78 ( .A1(a1stg_op[6]), .A2(a1stg_op[4]), .A3(n45), .A4(n4), .Y(
        n73) );
  NAND2X0_RVT U79 ( .A1(n61), .A2(n73), .Y(n76) );
  NAND2X0_RVT U80 ( .A1(n74), .A2(n76), .Y(n190) );
  INVX1_RVT U81 ( .A(n190), .Y(a1stg_fsdtoix) );
  AND2X1_RVT U82 ( .A1(a1stg_in1_exp_eq_0), .A2(a1stg_sngopa[0]), .Y(
        a1stg_denorm_sng_in1) );
  AND2X1_RVT U83 ( .A1(a1stg_sngopa[0]), .A2(n5), .Y(a1stg_norm_sng_in1) );
  AND2X1_RVT U84 ( .A1(a1stg_sngopa[0]), .A2(n6), .Y(a1stg_norm_sng_in2) );
  AND2X1_RVT U85 ( .A1(a1stg_in2_exp_eq_0), .A2(a1stg_sngopa[0]), .Y(
        a1stg_denorm_sng_in2) );
  NOR3X0_RVT U86 ( .A1(a1stg_op[3]), .A2(a1stg_op[5]), .A3(n85), .Y(n69) );
  NAND4X0_RVT U87 ( .A1(n69), .A2(n80), .A3(a1stg_op[2]), .A4(n46), .Y(n84) );
  OR2X1_RVT U88 ( .A1(n48), .A2(n84), .Y(n30) );
  INVX1_RVT U89 ( .A(n30), .Y(a1stg_fdtos) );
  INVX1_RVT U90 ( .A(add_ctl_rst_l), .Y(n242) );
  NAND3X0_RVT U91 ( .A1(a1stg_in2_53_32_neq_0), .A2(a1stg_sngopa[1]), .A3(n8), 
        .Y(n11) );
  NAND3X0_RVT U92 ( .A1(a1stg_in2_50_0_neq_0), .A2(a1stg_dblopa[1]), .A3(n9), 
        .Y(n10) );
  AOI21X1_RVT U93 ( .A1(n11), .A2(n10), .A3(a1stg_in2_exp_neq_ffs), .Y(
        a1stg_snan_in2) );
  OR2X1_RVT U94 ( .A1(a5stg_fxtod), .A2(a4stg_opdec_7_0[4]), .Y(a4stg_rnd_dbl)
         );
  NOR2X0_RVT U95 ( .A1(a4stg_rnd_mode[0]), .A2(a4stg_rnd_mode[1]), .Y(n17) );
  OA21X1_RVT U96 ( .A1(a4stg_frac_9_0_nx), .A2(a4stg_rnd_frac_11), .A3(
        a4stg_rnd_frac_10), .Y(n14) );
  OA221X1_RVT U97 ( .A1(a4stg_rnd_mode[0]), .A2(n13), .A3(n12), .A4(a4stg_sign), .A5(a4stg_rnd_mode[1]), .Y(n15) );
  AO22X1_RVT U98 ( .A1(n17), .A2(n14), .A3(n15), .A4(a4stg_frac_dbl_nx), .Y(
        n27) );
  OA21X1_RVT U99 ( .A1(a4stg_frac_38_0_nx), .A2(a4stg_rnd_frac_40), .A3(
        a4stg_rnd_frac_39), .Y(n16) );
  AO22X1_RVT U100 ( .A1(n17), .A2(n16), .A3(n15), .A4(a4stg_frac_sng_nx), .Y(
        n26) );
  AOI22X1_RVT U101 ( .A1(a5stg_fxtod), .A2(n27), .A3(a5stg_fixtos), .A4(n26), 
        .Y(n228) );
  INVX1_RVT U102 ( .A(a4stg_round), .Y(n149) );
  AO222X1_RVT U103 ( .A1(a4stg_opdec_7_0[6]), .A2(a4stg_exp[11]), .A3(
        a4stg_opdec_7_0[6]), .A4(n18), .A5(a4stg_exp[11]), .A6(
        a4stg_opdec_7_0[4]), .Y(n24) );
  NAND4X0_RVT U104 ( .A1(a4stg_exp[5]), .A2(a4stg_exp[6]), .A3(a4stg_exp[3]), 
        .A4(a4stg_exp[4]), .Y(n20) );
  NAND4X0_RVT U105 ( .A1(a4stg_exp[7]), .A2(a4stg_of_mask), .A3(a4stg_exp[1]), 
        .A4(a4stg_exp[2]), .Y(n19) );
  NOR2X0_RVT U106 ( .A1(n20), .A2(n19), .Y(n153) );
  NAND4X0_RVT U107 ( .A1(a4stg_exp[8]), .A2(a4stg_opdec_7_0[4]), .A3(
        a4stg_exp[9]), .A4(a4stg_exp[10]), .Y(n21) );
  NAND2X0_RVT U108 ( .A1(n22), .A2(n21), .Y(n150) );
  AND2X1_RVT U109 ( .A1(a4stg_exp[0]), .A2(n150), .Y(n23) );
  AO22X1_RVT U110 ( .A1(a4stg_of_mask), .A2(n24), .A3(n153), .A4(n23), .Y(
        a4stg_in_of) );
  INVX1_RVT U111 ( .A(a4stg_in_of), .Y(n231) );
  OA221X1_RVT U112 ( .A1(a4stg_opdec_7_0[3]), .A2(a4stg_opdec[29]), .A3(
        a4stg_opdec_7_0[3]), .A4(n149), .A5(n231), .Y(n226) );
  AO21X1_RVT U113 ( .A1(a4stg_opdec_7_0[3]), .A2(a4stg_of_mask), .A3(
        a4stg_opdec_7_0[5]), .Y(n25) );
  AO22X1_RVT U114 ( .A1(a4stg_opdec_7_0[4]), .A2(n27), .A3(n26), .A4(n25), .Y(
        n152) );
  INVX1_RVT U115 ( .A(n152), .Y(n227) );
  AO22X1_RVT U116 ( .A1(a5stg_fixtos_fxtod), .A2(n228), .A3(n226), .A4(n227), 
        .Y(add_exp_out_exp1) );
  OR2X1_RVT U117 ( .A1(a5stg_fixtos), .A2(a4stg_opdec_7_0[6]), .Y(
        a4stg_rnd_sng) );
  AND3X1_RVT U118 ( .A1(n69), .A2(n46), .A3(n48), .Y(n66) );
  NAND2X0_RVT U119 ( .A1(n66), .A2(n74), .Y(a1stg_faddsubop_inv) );
  INVX1_RVT U120 ( .A(a1stg_faddsubop_inv), .Y(n197) );
  AND2X1_RVT U121 ( .A1(n197), .A2(a1stg_op[2]), .Y(n75) );
  FADDX1_RVT U122 ( .A(a1stg_in1_63), .B(a1stg_in2_63), .CI(n75), .S(n31) );
  INVX1_RVT U123 ( .A(a1stg_in2_exp_neq_ffs), .Y(n171) );
  OR2X1_RVT U124 ( .A1(a1stg_in2_50_0_neq_0), .A2(a1stg_in2_51), .Y(n35) );
  OR2X1_RVT U125 ( .A1(a1stg_in2_53_32_neq_0), .A2(a1stg_in2_54), .Y(n34) );
  AO22X1_RVT U126 ( .A1(a1stg_dblopa[2]), .A2(n35), .A3(a1stg_sngopa[2]), .A4(
        n34), .Y(n28) );
  NAND2X0_RVT U127 ( .A1(n171), .A2(n28), .Y(n47) );
  INVX1_RVT U128 ( .A(a1stg_in1_exp_neq_ffs), .Y(n174) );
  OR2X1_RVT U129 ( .A1(a1stg_in1_53_32_neq_0), .A2(a1stg_in1_54), .Y(n32) );
  OR2X1_RVT U130 ( .A1(a1stg_in1_50_0_neq_0), .A2(a1stg_in1_51), .Y(n33) );
  AO22X1_RVT U131 ( .A1(a1stg_sngopa[2]), .A2(n32), .A3(a1stg_dblopa[2]), .A4(
        n33), .Y(n173) );
  NAND2X0_RVT U132 ( .A1(n174), .A2(n173), .Y(n29) );
  NAND2X0_RVT U133 ( .A1(n47), .A2(n29), .Y(a1stg_nan_in) );
  NAND2X0_RVT U134 ( .A1(n197), .A2(a1stg_nan_in), .Y(n176) );
  AND3X1_RVT U135 ( .A1(n31), .A2(n30), .A3(n176), .Y(a1stg_sub) );
  AO22X1_RVT U136 ( .A1(a1stg_sngopa[2]), .A2(n55), .A3(a1stg_dblopa[2]), .A4(
        n54), .Y(n37) );
  AO22X1_RVT U137 ( .A1(n56), .A2(a1stg_sngopa[2]), .A3(n58), .A4(
        a1stg_dblopa[2]), .Y(n36) );
  AND4X1_RVT U138 ( .A1(n171), .A2(n174), .A3(n37), .A4(n36), .Y(a1stg_2inf_in) );
  NAND3X0_RVT U139 ( .A1(n197), .A2(a1stg_sub), .A3(a1stg_2inf_in), .Y(n175)
         );
  INVX1_RVT U140 ( .A(n175), .Y(a2stg_frac1_in_nv) );
  OA22X1_RVT U141 ( .A1(a1stg_sngopa[3]), .A2(a1stg_dblopa[3]), .A3(n171), 
        .A4(n174), .Y(n249) );
  NOR2X0_RVT U142 ( .A1(n249), .A2(a1stg_faddsubop_inv), .Y(
        a2stg_frac2_in_frac1) );
  NAND2X0_RVT U143 ( .A1(a4stg_sign), .A2(a4stg_rnd_mode[1]), .Y(n38) );
  HADDX1_RVT U144 ( .A0(a4stg_rnd_mode[0]), .B0(n38), .SO(N1616) );
  INVX1_RVT U145 ( .A(N1616), .Y(a4stg_to_0) );
  NAND3X0_RVT U146 ( .A1(a1stg_in1_53_32_neq_0), .A2(a1stg_sngopa[1]), .A3(n39), .Y(n42) );
  NAND3X0_RVT U147 ( .A1(a1stg_in1_50_0_neq_0), .A2(a1stg_dblopa[1]), .A3(n40), 
        .Y(n41) );
  AO21X1_RVT U148 ( .A1(n42), .A2(n41), .A3(a1stg_in1_exp_neq_ffs), .Y(n172)
         );
  NAND2X0_RVT U149 ( .A1(a1stg_fdtos), .A2(n3), .Y(n88) );
  INVX1_RVT U150 ( .A(n88), .Y(a2stg_opdec_in[3]) );
  AND2X1_RVT U151 ( .A1(n77), .A2(n66), .Y(a1stg_faddsubs) );
  NAND2X0_RVT U152 ( .A1(a1stg_faddsubs), .A2(n3), .Y(n87) );
  AND4X1_RVT U153 ( .A1(a1stg_op[3]), .A2(n45), .A3(n44), .A4(n46), .Y(n59) );
  NAND2X0_RVT U154 ( .A1(a1stg_op[6]), .A2(n59), .Y(n64) );
  INVX1_RVT U155 ( .A(n64), .Y(n81) );
  NAND2X0_RVT U156 ( .A1(a1stg_op[0]), .A2(n81), .Y(n205) );
  INVX1_RVT U157 ( .A(n205), .Y(a1stg_fstod) );
  NAND4X0_RVT U158 ( .A1(a1stg_op[7]), .A2(a1stg_op[2]), .A3(n82), .A4(n46), 
        .Y(n68) );
  NOR4X1_RVT U159 ( .A1(a1stg_op[1]), .A2(a1stg_op[3]), .A3(a1stg_op[5]), .A4(
        n68), .Y(a2stg_opdec_in[1]) );
  INVX1_RVT U160 ( .A(n47), .Y(a1stg_nan_in2) );
  INVX0_RVT U161 ( .A(a3stg_opdec_9_0[3]), .Y(a3stg_fdtos_inv) );
  INVX0_RVT U162 ( .A(a4stg_opdec_7_0[7]), .Y(a4stg_fixtos_fxtod_inv) );
  OR2X1_RVT U170 ( .A1(a1stg_snan_in2), .A2(a1stg_snan_in1), .Y(n50) );
  AND4X1_RVT U171 ( .A1(n69), .A2(a1stg_op[4]), .A3(n74), .A4(n48), .Y(n83) );
  OA221X1_RVT U172 ( .A1(a1stg_op[2]), .A2(n50), .A3(n60), .A4(a1stg_nan_in), 
        .A5(n83), .Y(n49) );
  AOI221X1_RVT U173 ( .A1(a1stg_snan_in2), .A2(a1stg_fdtos), .A3(
        a1stg_snan_in2), .A4(a1stg_fstod), .A5(n49), .Y(n52) );
  NAND2X0_RVT U174 ( .A1(n197), .A2(n50), .Y(n51) );
  NAND3X0_RVT U175 ( .A1(n52), .A2(n175), .A3(n51), .Y(a1stg_nv) );
  AND3X1_RVT U177 ( .A1(a3stg_id[4]), .A2(a3stg_id[3]), .A3(a3stg_id[2]), .Y(
        N27) );
  AO22X1_RVT U178 ( .A1(a1stg_in1_54), .A2(a1stg_sngopa[1]), .A3(a1stg_in1_51), 
        .A4(a1stg_dblopa[1]), .Y(n53) );
  AND2X1_RVT U179 ( .A1(n174), .A2(n53), .Y(a1stg_qnan_in1) );
  OA221X1_RVT U180 ( .A1(a1stg_dblopa[3]), .A2(n56), .A3(a1stg_dblopa[3]), 
        .A4(n55), .A5(n54), .Y(n57) );
  AND4X1_RVT U181 ( .A1(n58), .A2(a1stg_in1_exp_eq_0), .A3(a1stg_in2_exp_eq_0), 
        .A4(n57), .Y(a1stg_2zero_in) );
  AND2X1_RVT U182 ( .A1(inq_add), .A2(inq_op[7]), .Y(a1stg_op_in[7]) );
  AND2X1_RVT U183 ( .A1(inq_add), .A2(inq_op[6]), .Y(a1stg_op_in[6]) );
  AND2X1_RVT U184 ( .A1(inq_add), .A2(inq_op[5]), .Y(a1stg_op_in[5]) );
  AND2X1_RVT U185 ( .A1(inq_add), .A2(inq_op[4]), .Y(a1stg_op_in[4]) );
  AND2X1_RVT U186 ( .A1(inq_add), .A2(inq_op[3]), .Y(a1stg_op_in[3]) );
  AND2X1_RVT U187 ( .A1(inq_add), .A2(inq_op[2]), .Y(a1stg_op_in[2]) );
  AND2X1_RVT U188 ( .A1(inq_add), .A2(inq_op[1]), .Y(a1stg_op_in[1]) );
  AND2X1_RVT U189 ( .A1(inq_add), .A2(inq_op[0]), .Y(a1stg_op_in[0]) );
  AND2X1_RVT U190 ( .A1(a1stg_dblop), .A2(n3), .Y(a2stg_opdec_in[30]) );
  INVX1_RVT U191 ( .A(a2stg_opdec_in[1]), .Y(n72) );
  NAND2X0_RVT U192 ( .A1(n59), .A2(n82), .Y(n67) );
  NAND2X0_RVT U193 ( .A1(n72), .A2(n67), .Y(n208) );
  NAND2X0_RVT U194 ( .A1(n69), .A2(n74), .Y(n63) );
  NAND2X0_RVT U195 ( .A1(a1stg_op[4]), .A2(n60), .Y(n62) );
  INVX1_RVT U196 ( .A(n61), .Y(n79) );
  NAND2X0_RVT U197 ( .A1(n79), .A2(n74), .Y(n243) );
  OA221X1_RVT U198 ( .A1(n63), .A2(a1stg_op[7]), .A3(n63), .A4(n62), .A5(n243), 
        .Y(n65) );
  NAND4X0_RVT U199 ( .A1(n204), .A2(n65), .A3(n84), .A4(n64), .Y(n93) );
  AND2X1_RVT U200 ( .A1(n93), .A2(n3), .Y(a2stg_opdec_in[29]) );
  AND2X1_RVT U201 ( .A1(n80), .A2(n66), .Y(a1stg_faddsubd) );
  AND2X1_RVT U202 ( .A1(a1stg_faddsubd), .A2(n3), .Y(a2stg_opdec_in[4]) );
  AO221X1_RVT U203 ( .A1(n3), .A2(n81), .A3(n3), .A4(n86), .A5(
        a2stg_opdec_in[4]), .Y(a2stg_opdec_in[28]) );
  NAND3X0_RVT U204 ( .A1(n70), .A2(n69), .A3(n3), .Y(n71) );
  NAND3X0_RVT U205 ( .A1(n72), .A2(n87), .A3(n71), .Y(a2stg_opdec_in[27]) );
  AND3X1_RVT U206 ( .A1(n79), .A2(n74), .A3(n3), .Y(a2stg_opdec_in[26]) );
  AND3X1_RVT U207 ( .A1(n78), .A2(n74), .A3(n3), .Y(a2stg_opdec_in[25]) );
  AND2X1_RVT U208 ( .A1(n197), .A2(n3), .Y(a2stg_opdec_in[24]) );
  AND2X1_RVT U209 ( .A1(n75), .A2(n3), .Y(a2stg_opdec_in[23]) );
  AND3X1_RVT U210 ( .A1(n80), .A2(n76), .A3(n3), .Y(a2stg_opdec_in[21]) );
  AND3X1_RVT U211 ( .A1(n77), .A2(n76), .A3(n3), .Y(a2stg_opdec_in[20]) );
  AND2X1_RVT U212 ( .A1(a1stg_fstod), .A2(n3), .Y(a2stg_opdec_in[18]) );
  AND2X1_RVT U213 ( .A1(n77), .A2(n78), .Y(a1stg_fstoi) );
  AND2X1_RVT U214 ( .A1(a1stg_fstoi), .A2(n3), .Y(a2stg_opdec_in[17]) );
  AND2X1_RVT U215 ( .A1(n77), .A2(n79), .Y(a1stg_fstox) );
  AND2X1_RVT U216 ( .A1(a1stg_fstox), .A2(n3), .Y(a2stg_opdec_in[16]) );
  AND2X1_RVT U217 ( .A1(n80), .A2(n78), .Y(a1stg_fdtoi) );
  AND2X1_RVT U218 ( .A1(a1stg_fdtoi), .A2(n3), .Y(a2stg_opdec_in[15]) );
  AND2X1_RVT U219 ( .A1(n80), .A2(n79), .Y(a1stg_fdtox) );
  AND2X1_RVT U220 ( .A1(a1stg_fdtox), .A2(n3), .Y(a2stg_opdec_in[14]) );
  AND2X1_RVT U221 ( .A1(a1stg_fsdtoix), .A2(n3), .Y(a2stg_opdec_in[19]) );
  OR2X1_RVT U222 ( .A1(a2stg_opdec_in[3]), .A2(a2stg_opdec_in[19]), .Y(
        a2stg_opdec_in[13]) );
  AND2X1_RVT U223 ( .A1(a1stg_op[6]), .A2(a2stg_opdec_in[1]), .Y(
        a2stg_opdec_in[12]) );
  AND2X1_RVT U224 ( .A1(n81), .A2(n3), .Y(a2stg_opdec_in[2]) );
  AND2X1_RVT U225 ( .A1(a2stg_opdec_in[2]), .A2(n82), .Y(a2stg_opdec_in[11])
         );
  AND2X1_RVT U226 ( .A1(a2stg_opdec_in[1]), .A2(n85), .Y(a2stg_opdec_in[10])
         );
  AND2X1_RVT U227 ( .A1(n83), .A2(n3), .Y(a2stg_opdec_in[9]) );
  NAND2X0_RVT U228 ( .A1(a1stg_faddsubop_inv), .A2(n84), .Y(n248) );
  AND2X1_RVT U229 ( .A1(n248), .A2(n3), .Y(a2stg_opdec_in[22]) );
  OR2X1_RVT U230 ( .A1(a2stg_opdec_in[2]), .A2(a2stg_opdec_in[22]), .Y(
        a2stg_opdec_in[8]) );
  AND2X1_RVT U231 ( .A1(n86), .A2(n85), .Y(a2stg_opdec_in[0]) );
  OR2X1_RVT U232 ( .A1(a2stg_opdec_in[1]), .A2(a2stg_opdec_in[0]), .Y(
        a2stg_opdec_in[7]) );
  NAND2X0_RVT U233 ( .A1(n88), .A2(n87), .Y(a2stg_opdec_in[6]) );
  INVX1_RVT U234 ( .A(a3stg_opdec_9_0[8]), .Y(n121) );
  AO22X1_RVT U235 ( .A1(a3stg_opdec_9_0[8]), .A2(a3stg_rnd_mode[1]), .A3(n121), 
        .A4(a4stg_rnd_mode2[1]), .Y(a4stg_rnd_mode_in[1]) );
  AO22X1_RVT U236 ( .A1(a3stg_opdec_9_0[8]), .A2(a3stg_rnd_mode[0]), .A3(n121), 
        .A4(a4stg_rnd_mode2[0]), .Y(a4stg_rnd_mode_in[0]) );
  INVX1_RVT U237 ( .A(a5stg_fixtos_fxtod), .Y(n230) );
  AND2X1_RVT U238 ( .A1(n230), .A2(a4stg_fixtos_fxtod_inv), .Y(n89) );
  AO22X1_RVT U239 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec[33]), .A3(n89), 
        .A4(a4stg_opdec[33]), .Y(a6stg_opdec_in[33]) );
  AO22X1_RVT U240 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec[32]), .A3(n89), 
        .A4(a4stg_opdec[32]), .Y(a6stg_opdec_in[32]) );
  AO22X1_RVT U241 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec[31]), .A3(n89), 
        .A4(a4stg_opdec[31]), .Y(a6stg_opdec_in[31]) );
  AO22X1_RVT U242 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec[30]), .A3(n89), 
        .A4(a4stg_opdec[30]), .Y(a6stg_opdec_in[30]) );
  AO22X1_RVT U243 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec_9), .A3(n89), 
        .A4(a4stg_fcmpop), .Y(a6stg_opdec_in_9) );
  AO22X1_RVT U244 ( .A1(a5stg_fixtos_fxtod), .A2(a5stg_opdec[34]), .A3(
        a4stg_opdec[34]), .A4(n89), .Y(a6stg_opdec_in[34]) );
  OA21X1_RVT U245 ( .A1(n92), .A2(a6stg_opdec_in[34]), .A3(add_ctl_rst_l), .Y(
        a6stg_fadd_in) );
  AND2X1_RVT U246 ( .A1(n230), .A2(a6stg_step), .Y(n90) );
  AND2X1_RVT U247 ( .A1(a5stg_fixtos_fxtod), .A2(a6stg_step), .Y(n91) );
  AO222X1_RVT U248 ( .A1(n92), .A2(add_id_out[9]), .A3(n90), .A4(a4stg_id[9]), 
        .A5(n91), .A6(a5stg_id[9]), .Y(add_id_out_in[9]) );
  AO222X1_RVT U249 ( .A1(n92), .A2(add_id_out[8]), .A3(n91), .A4(a5stg_id[8]), 
        .A5(a4stg_id[8]), .A6(n90), .Y(add_id_out_in[8]) );
  AO222X1_RVT U250 ( .A1(n92), .A2(add_id_out[7]), .A3(n91), .A4(a5stg_id[7]), 
        .A5(a4stg_id[7]), .A6(n90), .Y(add_id_out_in[7]) );
  AO222X1_RVT U251 ( .A1(n92), .A2(add_id_out[6]), .A3(n91), .A4(a5stg_id[6]), 
        .A5(a4stg_id[6]), .A6(n90), .Y(add_id_out_in[6]) );
  AO222X1_RVT U252 ( .A1(n92), .A2(add_id_out[5]), .A3(n91), .A4(a5stg_id[5]), 
        .A5(a4stg_id[5]), .A6(n90), .Y(add_id_out_in[5]) );
  AO222X1_RVT U253 ( .A1(n92), .A2(add_id_out[4]), .A3(n91), .A4(a5stg_id[4]), 
        .A5(a4stg_id[4]), .A6(n90), .Y(add_id_out_in[4]) );
  AO222X1_RVT U254 ( .A1(n92), .A2(add_id_out[3]), .A3(n91), .A4(a5stg_id[3]), 
        .A5(a4stg_id[3]), .A6(n90), .Y(add_id_out_in[3]) );
  AO222X1_RVT U255 ( .A1(n92), .A2(add_id_out[2]), .A3(n91), .A4(a5stg_id[2]), 
        .A5(a4stg_id[2]), .A6(n90), .Y(add_id_out_in[2]) );
  AO222X1_RVT U256 ( .A1(n92), .A2(add_id_out[1]), .A3(n91), .A4(a5stg_id[1]), 
        .A5(a4stg_id[1]), .A6(n90), .Y(add_id_out_in[1]) );
  AO222X1_RVT U257 ( .A1(n92), .A2(add_id_out[0]), .A3(n91), .A4(a5stg_id[0]), 
        .A5(a4stg_id[0]), .A6(n90), .Y(add_id_out_in[0]) );
  AND2X1_RVT U258 ( .A1(a4stg_fcmpop), .A2(a4stg_fcc[1]), .Y(add_fcc_out_in[1]) );
  AND2X1_RVT U259 ( .A1(a4stg_fcmpop), .A2(a4stg_fcc[0]), .Y(add_fcc_out_in[0]) );
  NOR4X1_RVT U260 ( .A1(a2stg_opdec[34]), .A2(a5stg_opdec[34]), .A3(
        a4stg_opdec[34]), .A4(n93), .Y(n95) );
  INVX1_RVT U261 ( .A(a3stg_opdec[34]), .Y(n145) );
  NAND3X0_RVT U262 ( .A1(n95), .A2(n94), .A3(n145), .Y(add_pipe_active_in) );
  AND2X1_RVT U263 ( .A1(a2stg_opdec_24_21[0]), .A2(n96), .Y(n131) );
  NOR3X0_RVT U264 ( .A1(a2stg_nan_in), .A2(n131), .A3(n114), .Y(a3stg_sub_in)
         );
  OAI22X1_RVT U265 ( .A1(a2stg_snan_in2), .A2(a2stg_snan_in1), .A3(
        a2stg_nan_in2), .A4(a2stg_qnan_in1), .Y(n108) );
  NAND2X0_RVT U266 ( .A1(a2stg_in2_neq_in1_frac), .A2(a2stg_in2_eq_in1_exp), 
        .Y(n115) );
  AND4X1_RVT U267 ( .A1(a2stg_rnd_mode[1]), .A2(n98), .A3(a2stg_rnd_mode[0]), 
        .A4(n97), .Y(n105) );
  AO21X1_RVT U268 ( .A1(a2stg_in2_eq_in1_exp), .A2(a2stg_in2_gt_in1_frac), 
        .A3(a2stg_in2_gt_in1_exp), .Y(n100) );
  INVX1_RVT U269 ( .A(n100), .Y(n116) );
  NAND2X0_RVT U270 ( .A1(a2stg_2inf_in), .A2(a2stg_sub), .Y(n99) );
  AND3X1_RVT U271 ( .A1(n116), .A2(n115), .A3(n99), .Y(n104) );
  INVX1_RVT U272 ( .A(a2stg_sign2), .Y(n126) );
  OA221X1_RVT U273 ( .A1(a2stg_sign1), .A2(n115), .A3(a2stg_sign1), .A4(n100), 
        .A5(n99), .Y(n101) );
  OA222X1_RVT U274 ( .A1(a2stg_opdec_28), .A2(a2stg_sign2), .A3(n102), .A4(
        n126), .A5(n105), .A6(n101), .Y(n103) );
  AO221X1_RVT U275 ( .A1(a2stg_sign1), .A2(n105), .A3(a2stg_sign1), .A4(n104), 
        .A5(n103), .Y(n106) );
  AO22X1_RVT U276 ( .A1(a2stg_sign1), .A2(n108), .A3(n107), .A4(n106), .Y(n112) );
  NAND2X0_RVT U277 ( .A1(a2stg_snan_in1), .A2(a2stg_qnan_in2), .Y(n109) );
  NAND3X0_RVT U278 ( .A1(a2stg_faddsubop), .A2(n110), .A3(n109), .Y(n111) );
  AO22X1_RVT U279 ( .A1(a2stg_faddsubop), .A2(n112), .A3(a2stg_sign2), .A4(
        n111), .Y(a3stg_sign_in) );
  NAND2X0_RVT U280 ( .A1(n115), .A2(n114), .Y(n113) );
  OAI22X1_RVT U281 ( .A1(n116), .A2(n113), .A3(a2stg_2zero_in), .A4(n114), .Y(
        n118) );
  AND3X1_RVT U282 ( .A1(n116), .A2(n115), .A3(n114), .Y(n119) );
  AO221X1_RVT U283 ( .A1(a2stg_sign2), .A2(n118), .A3(n126), .A4(n119), .A5(
        a2stg_nan_in), .Y(n117) );
  AND2X1_RVT U284 ( .A1(a2stg_opdec_9_0[9]), .A2(n117), .Y(a2stg_cc[1]) );
  AO221X1_RVT U285 ( .A1(a2stg_sign2), .A2(n119), .A3(n126), .A4(n118), .A5(
        a2stg_nan_in), .Y(n120) );
  AND2X1_RVT U286 ( .A1(a2stg_opdec_9_0[9]), .A2(n120), .Y(a2stg_cc[0]) );
  AO22X1_RVT U287 ( .A1(a3stg_opdec_9_0[8]), .A2(a3stg_sign), .A3(n121), .A4(
        a4stg_sign2), .Y(a4stg_sign_in) );
  AND2X1_RVT U288 ( .A1(a4stg_fcmpop), .A2(a4stg_cc[1]), .Y(add_cc_out_in[1])
         );
  AND2X1_RVT U289 ( .A1(a4stg_fcmpop), .A2(a4stg_cc[0]), .Y(add_cc_out_in[0])
         );
  NOR4X1_RVT U290 ( .A1(a2stg_expadd[8]), .A2(a2stg_expadd[10]), .A3(
        a2stg_expadd[2]), .A4(a2stg_expadd[0]), .Y(n129) );
  NOR4X1_RVT U291 ( .A1(a2stg_expadd[1]), .A2(a2stg_expadd[5]), .A3(
        a2stg_expadd[3]), .A4(a2stg_expadd[4]), .Y(n128) );
  NAND2X0_RVT U292 ( .A1(a2stg_frac2lo_neq_0), .A2(a2stg_opdec[31]), .Y(n122)
         );
  NAND3X0_RVT U293 ( .A1(n124), .A2(n123), .A3(n122), .Y(n125) );
  NOR4X1_RVT U294 ( .A1(a2stg_expadd[6]), .A2(a2stg_frac2hi_neq_0), .A3(n126), 
        .A4(n125), .Y(n127) );
  NAND3X0_RVT U295 ( .A1(n129), .A2(n128), .A3(n127), .Y(n130) );
  AO21X1_RVT U296 ( .A1(n131), .A2(n130), .A3(a2stg_nv), .Y(a3stg_nv_in) );
  OR2X1_RVT U297 ( .A1(a2stg_exp[10]), .A2(a2stg_exp[11]), .Y(n194) );
  NOR4X1_RVT U298 ( .A1(a2stg_exp[9]), .A2(a2stg_exp[7]), .A3(a2stg_exp[8]), 
        .A4(n194), .Y(n132) );
  INVX1_RVT U299 ( .A(n132), .Y(n195) );
  AO22X1_RVT U300 ( .A1(a2stg_opdec_24_21[1]), .A2(n195), .A3(
        a2stg_opdec_24_21[2]), .A4(n194), .Y(a2stg_nx_tmp1) );
  AO22X1_RVT U301 ( .A1(n133), .A2(a2stg_opdec_24_21[2]), .A3(n132), .A4(
        a2stg_opdec_24_21[1]), .Y(n136) );
  NOR3X0_RVT U302 ( .A1(a2stg_exp[6]), .A2(a2stg_exp[10]), .A3(n142), .Y(n217)
         );
  NOR4X1_RVT U303 ( .A1(a2stg_exp[3]), .A2(a2stg_exp[1]), .A3(a2stg_exp[2]), 
        .A4(a2stg_exp[4]), .Y(n134) );
  INVX1_RVT U304 ( .A(a2stg_frac2hi_neq_0), .Y(n137) );
  NAND4X0_RVT U305 ( .A1(n217), .A2(n134), .A3(n137), .A4(n138), .Y(n135) );
  AO222X1_RVT U306 ( .A1(n136), .A2(a2stg_frac2lo_neq_0), .A3(n136), .A4(
        a2stg_frac2_63), .A5(n136), .A6(n135), .Y(a2stg_nx_tmp2) );
  AND2X1_RVT U307 ( .A1(a2stg_exp[1]), .A2(a2stg_exp[2]), .Y(n214) );
  AND4X1_RVT U308 ( .A1(a2stg_sign2), .A2(a2stg_exp[3]), .A3(a2stg_exp[0]), 
        .A4(n137), .Y(n144) );
  NAND4X0_RVT U309 ( .A1(a2stg_exp[10]), .A2(a2stg_exp[4]), .A3(n139), .A4(
        n138), .Y(n140) );
  NOR4X1_RVT U310 ( .A1(a2stg_exp[11]), .A2(n142), .A3(n141), .A4(n140), .Y(
        n143) );
  AND4X1_RVT U311 ( .A1(a2stg_frac2lo_neq_0), .A2(n214), .A3(n144), .A4(n143), 
        .Y(a2stg_nx_tmp3) );
  OR2X1_RVT U312 ( .A1(a3stg_opdec_9_0[7]), .A2(n145), .Y(n147) );
  INVX1_RVT U313 ( .A(n147), .Y(n148) );
  AO22X1_RVT U314 ( .A1(n148), .A2(a3stg_nv), .A3(n147), .A4(a4stg_nv2), .Y(
        a4stg_nv_in) );
  AO22X1_RVT U315 ( .A1(n148), .A2(a3stg_of_mask), .A3(n147), .A4(
        a4stg_of_mask2), .Y(a4stg_of_mask_in) );
  OA221X1_RVT U316 ( .A1(a3stg_fsdtoix_nx), .A2(a3stg_opdec[30]), .A3(
        a3stg_fsdtoix_nx), .A4(a3stg_fsdtoi_nx), .A5(a3stg_nx_tmp1), .Y(n146)
         );
  AO221X1_RVT U317 ( .A1(a3stg_a2_expadd_11), .A2(a3stg_nx_tmp2), .A3(
        a3stg_a2_expadd_11), .A4(n146), .A5(a3stg_nx_tmp3), .Y(a3stg_nx) );
  AO22X1_RVT U318 ( .A1(n148), .A2(a3stg_nx), .A3(n147), .A4(a4stg_nx2), .Y(
        a4stg_nx_in) );
  AO22X1_RVT U319 ( .A1(a4stg_opdec_7_0[6]), .A2(a4stg_opdec_7_0[3]), .A3(n150), .A4(n149), .Y(n151) );
  AND3X1_RVT U320 ( .A1(n153), .A2(n152), .A3(n151), .Y(add_of_out_tmp1_in) );
  NAND4X0_RVT U321 ( .A1(a4stg_opdec[29]), .A2(a4stg_round), .A3(
        a4stg_shl_data_neq_0), .A4(n157), .Y(n163) );
  NOR2X0_RVT U322 ( .A1(a4stg_exp[9]), .A2(a4stg_exp[10]), .Y(n156) );
  NOR4X1_RVT U323 ( .A1(a4stg_exp[2]), .A2(a4stg_exp[5]), .A3(a4stg_exp[6]), 
        .A4(a4stg_exp[3]), .Y(n155) );
  NOR4X1_RVT U324 ( .A1(a4stg_exp[4]), .A2(a4stg_exp[8]), .A3(a4stg_exp[0]), 
        .A4(a4stg_faddsub_dtosop), .Y(n154) );
  NAND4X0_RVT U325 ( .A1(n156), .A2(a4stg_frac_neq_0), .A3(n155), .A4(n154), 
        .Y(n162) );
  NAND2X0_RVT U326 ( .A1(a4stg_round), .A2(n157), .Y(n158) );
  NAND3X0_RVT U327 ( .A1(n160), .A2(n159), .A3(n158), .Y(n161) );
  OAI22X1_RVT U328 ( .A1(a4stg_denorm_inv), .A2(n163), .A3(n162), .A4(n161), 
        .Y(a4stg_uf) );
  AND2X1_RVT U330 ( .A1(a4stg_rnd_sng), .A2(a4stg_frac_sng_nx), .Y(n165) );
  NAND2X0_RVT U331 ( .A1(a4stg_round), .A2(a4stg_opdec_7_0[5]), .Y(n164) );
  AND2X1_RVT U332 ( .A1(n165), .A2(n164), .Y(n169) );
  AND2X1_RVT U333 ( .A1(a4stg_rnd_dbl), .A2(a4stg_frac_dbl_nx), .Y(n167) );
  NAND2X0_RVT U334 ( .A1(a4stg_opdec_7_0[4]), .A2(a4stg_round), .Y(n166) );
  AND2X1_RVT U335 ( .A1(n167), .A2(n166), .Y(n168) );
  AO221X1_RVT U336 ( .A1(a4stg_of_mask), .A2(n169), .A3(a4stg_of_mask), .A4(
        n168), .A5(a4stg_nx), .Y(add_nx_out_in) );
  AO21X1_RVT U337 ( .A1(add_of_out_cout), .A2(add_of_out_tmp1), .A3(
        add_of_out_tmp2), .Y(add_exc_out[3]) );
  OR2X1_RVT U338 ( .A1(add_nx_out), .A2(add_exc_out[3]), .Y(add_exc_out_0) );
  AO22X1_RVT U339 ( .A1(a1stg_in2_54), .A2(a1stg_sngopa[1]), .A3(a1stg_in2_51), 
        .A4(a1stg_dblopa[1]), .Y(n170) );
  AND2X1_RVT U340 ( .A1(n171), .A2(n170), .Y(a1stg_qnan_in2) );
  AO21X1_RVT U341 ( .A1(a1stg_qnan_in2), .A2(n172), .A3(a1stg_snan_in2), .Y(
        a2stg_frac1_in_frac1) );
  NAND3X0_RVT U342 ( .A1(a1stg_nan_in2), .A2(n174), .A3(n173), .Y(
        a1stg_2nan_in_inv) );
  OA21X1_RVT U343 ( .A1(a1stg_2nan_in_inv), .A2(a2stg_frac1_in_frac1), .A3(
        n197), .Y(a2stg_frac1_in_frac2) );
  NAND2X0_RVT U344 ( .A1(n176), .A2(n175), .Y(a2stg_frac1_in_qnan) );
  AND3X1_RVT U345 ( .A1(a1stg_sub), .A2(a1stg_2inf_in), .A3(a1stg_faddsubd), 
        .Y(a2stg_frac1_in_nv_dbl) );
  AND2X1_RVT U346 ( .A1(a1stg_snan_in2), .A2(a1stg_faddsubop_inv), .Y(
        a2stg_frac2_in_qnan) );
  INVX1_RVT U347 ( .A(n198), .Y(n180) );
  NAND2X0_RVT U348 ( .A1(n178), .A2(n248), .Y(n181) );
  AND4X1_RVT U349 ( .A1(a1stg_expadd4_inv[7]), .A2(a1stg_expadd4_inv[8]), .A3(
        a1stg_expadd4_inv[9]), .A4(a1stg_expadd4_inv[10]), .Y(n179) );
  AND2X1_RVT U350 ( .A1(a1stg_expadd4_inv[6]), .A2(n179), .Y(n199) );
  NAND2X0_RVT U351 ( .A1(n197), .A2(a1stg_expadd1[11]), .Y(n241) );
  OA22X1_RVT U352 ( .A1(n180), .A2(n181), .A3(n199), .A4(n241), .Y(n245) );
  OA22X1_RVT U353 ( .A1(a1stg_expadd4_inv[4]), .A2(n241), .A3(a1stg_expadd2[4]), .A4(n190), .Y(n183) );
  INVX1_RVT U354 ( .A(n181), .Y(n240) );
  NAND2X0_RVT U355 ( .A1(n240), .A2(a1stg_expadd1[4]), .Y(n182) );
  NAND3X0_RVT U356 ( .A1(n245), .A2(n183), .A3(n182), .Y(a2stg_shr_cnt_in[4])
         );
  NAND2X0_RVT U357 ( .A1(a1stg_expadd1[3]), .A2(n240), .Y(n185) );
  OA22X1_RVT U358 ( .A1(a1stg_expadd4_inv[3]), .A2(n241), .A3(a1stg_expadd2[3]), .A4(n190), .Y(n184) );
  NAND3X0_RVT U359 ( .A1(n185), .A2(n184), .A3(n245), .Y(a2stg_shr_cnt_in[3])
         );
  NAND2X0_RVT U360 ( .A1(a1stg_expadd1[2]), .A2(n240), .Y(n187) );
  OA22X1_RVT U361 ( .A1(a1stg_expadd4_inv[2]), .A2(n241), .A3(a1stg_expadd2[2]), .A4(n190), .Y(n186) );
  NAND3X0_RVT U362 ( .A1(n187), .A2(n186), .A3(n245), .Y(a2stg_shr_cnt_in[2])
         );
  NAND2X0_RVT U363 ( .A1(a1stg_expadd1[1]), .A2(n240), .Y(n189) );
  OA22X1_RVT U364 ( .A1(a1stg_expadd4_inv[1]), .A2(n241), .A3(a1stg_expadd2[1]), .A4(n190), .Y(n188) );
  NAND3X0_RVT U365 ( .A1(n189), .A2(n188), .A3(n245), .Y(a2stg_shr_cnt_in[1])
         );
  NAND2X0_RVT U366 ( .A1(n240), .A2(a1stg_expadd1[0]), .Y(n192) );
  OA22X1_RVT U367 ( .A1(a1stg_expadd4_inv[0]), .A2(n241), .A3(a1stg_expadd2[0]), .A4(n190), .Y(n191) );
  NAND3X0_RVT U368 ( .A1(n192), .A2(n191), .A3(n245), .Y(a2stg_shr_cnt_in[0])
         );
  AND2X1_RVT U369 ( .A1(a2stg_opdec_24_21[3]), .A2(a6stg_step), .Y(
        a2stg_shr_frac2_shr_int) );
  AO22X1_RVT U370 ( .A1(a2stg_opdec_19_11[6]), .A2(n195), .A3(
        a2stg_opdec_19_11[4]), .A4(n194), .Y(n193) );
  AND2X1_RVT U371 ( .A1(a6stg_step), .A2(n193), .Y(a2stg_shr_frac2_shr_dbl) );
  AO22X1_RVT U372 ( .A1(a2stg_opdec_19_11[7]), .A2(n195), .A3(
        a2stg_opdec_19_11[5]), .A4(n194), .Y(n196) );
  AND2X1_RVT U373 ( .A1(a6stg_step), .A2(n196), .Y(a2stg_shr_frac2_shr_sng) );
  AND2X1_RVT U374 ( .A1(a2stg_opdec_24_21[0]), .A2(a6stg_step), .Y(
        a2stg_shr_frac2_max) );
  AND2X1_RVT U375 ( .A1(n197), .A2(a1stg_sub), .Y(n207) );
  NAND3X0_RVT U376 ( .A1(a1stg_expadd1[11]), .A2(a1stg_expadd4_inv[0]), .A3(
        n199), .Y(n200) );
  NAND2X0_RVT U377 ( .A1(n201), .A2(n200), .Y(n202) );
  AO22X1_RVT U378 ( .A1(a1stg_in2_63), .A2(n208), .A3(n207), .A4(n202), .Y(
        a2stg_fracadd_frac2_inv_in) );
  AND2X1_RVT U379 ( .A1(n207), .A2(n203), .Y(a2stg_fracadd_frac2_inv_shr1_in)
         );
  OA22X1_RVT U380 ( .A1(a1stg_in2_63), .A2(n204), .A3(a1stg_sub), .A4(
        a1stg_faddsubop_inv), .Y(n206) );
  NAND2X0_RVT U381 ( .A1(n206), .A2(n205), .Y(a2stg_fracadd_frac2_in) );
  AO21X1_RVT U382 ( .A1(a1stg_in2_63), .A2(n208), .A3(n207), .Y(
        a2stg_fracadd_cin_in) );
  AND4X1_RVT U383 ( .A1(a2stg_exp[5]), .A2(a2stg_exp[3]), .A3(a2stg_exp[4]), 
        .A4(a2stg_exp[0]), .Y(n209) );
  NAND4X0_RVT U384 ( .A1(a2stg_exp[7]), .A2(a2stg_exp[6]), .A3(n214), .A4(n209), .Y(n212) );
  INVX1_RVT U385 ( .A(n212), .Y(n210) );
  AND2X1_RVT U386 ( .A1(n210), .A2(a2stg_opdec_19_11[8]), .Y(a3stg_exp_7ff) );
  NAND4X0_RVT U387 ( .A1(a2stg_exp[9]), .A2(a2stg_exp[8]), .A3(a2stg_exp[10]), 
        .A4(n210), .Y(n213) );
  AND2X1_RVT U388 ( .A1(n211), .A2(a2stg_opdec_9_0[3]), .Y(a3stg_exp_ff) );
  AO22X1_RVT U389 ( .A1(a2stg_opdec_9_0[3]), .A2(n213), .A3(
        a2stg_opdec_19_11[8]), .A4(n212), .Y(a3stg_exp_add) );
  OR2X1_RVT U390 ( .A1(a2stg_exp[3]), .A2(n214), .Y(n215) );
  NAND3X0_RVT U391 ( .A1(n215), .A2(a2stg_exp[4]), .A3(a2stg_exp[5]), .Y(n216)
         );
  AND3X1_RVT U392 ( .A1(n217), .A2(a2stg_faddsubop), .A3(n216), .Y(
        a2stg_expdec_neq_0) );
  NAND2X0_RVT U393 ( .A1(a3stg_exp[4]), .A2(a3stg_denorm), .Y(n224) );
  NAND2X0_RVT U394 ( .A1(a3stg_lead0[5]), .A2(n225), .Y(n222) );
  AO22X1_RVT U395 ( .A1(a3stg_exp[5]), .A2(n219), .A3(a3stg_lead0[4]), .A4(
        n218), .Y(a4stg_shl_cnt_in[9]) );
  NAND2X0_RVT U396 ( .A1(a3stg_exp[5]), .A2(a3stg_denorm), .Y(n221) );
  OAI22X1_RVT U397 ( .A1(a3stg_lead0[4]), .A2(n222), .A3(a3stg_exp[4]), .A4(
        n221), .Y(a4stg_shl_cnt_in[8]) );
  NAND2X0_RVT U398 ( .A1(a3stg_lead0[4]), .A2(n225), .Y(n223) );
  OAI22X1_RVT U399 ( .A1(a3stg_lead0[5]), .A2(n223), .A3(a3stg_exp[5]), .A4(
        n224), .Y(a4stg_shl_cnt_in[7]) );
  OR2X1_RVT U400 ( .A1(a3stg_exp[4]), .A2(a3stg_exp[5]), .Y(n220) );
  AOI222X1_RVT U401 ( .A1(n225), .A2(a3stg_lead0[4]), .A3(n225), .A4(
        a3stg_lead0[5]), .A5(n220), .A6(a3stg_denorm), .Y(a4stg_shl_cnt_in[6])
         );
  NAND2X0_RVT U402 ( .A1(n222), .A2(n221), .Y(a4stg_shl_cnt_in[5]) );
  NAND2X0_RVT U403 ( .A1(n224), .A2(n223), .Y(a4stg_shl_cnt_in[4]) );
  AO22X1_RVT U404 ( .A1(a3stg_denorm), .A2(a3stg_exp[3]), .A3(n225), .A4(
        a3stg_lead0[3]), .Y(a4stg_shl_cnt_in[3]) );
  AO22X1_RVT U405 ( .A1(a3stg_denorm), .A2(a3stg_exp[2]), .A3(n225), .A4(
        a3stg_lead0[2]), .Y(a4stg_shl_cnt_in[2]) );
  AO22X1_RVT U406 ( .A1(a3stg_denorm), .A2(a3stg_exp[1]), .A3(n225), .A4(
        a3stg_lead0[1]), .Y(a4stg_shl_cnt_in[1]) );
  AO22X1_RVT U407 ( .A1(a3stg_denorm), .A2(a3stg_exp[0]), .A3(n225), .A4(
        a3stg_lead0[0]), .Y(a4stg_shl_cnt_in[0]) );
  OR2X1_RVT U408 ( .A1(a4stg_fsdtoix), .A2(add_exp_out_exp1), .Y(
        add_frac_out_rnd_frac) );
  INVX1_RVT U409 ( .A(n226), .Y(n229) );
  OAI22X1_RVT U410 ( .A1(n228), .A2(n230), .A3(n227), .A4(n229), .Y(
        add_exp_out_expinc) );
  NAND2X0_RVT U411 ( .A1(n230), .A2(n229), .Y(add_exp_out_exp) );
  OA222X1_RVT U412 ( .A1(a4stg_opdec_7_0[2]), .A2(a4stg_opdec[29]), .A3(
        a4stg_opdec_7_0[2]), .A4(n231), .A5(a4stg_opdec_7_0[2]), .A6(
        a4stg_round), .Y(add_exp_out_expadd) );
  INVX1_RVT U413 ( .A(a3stg_id[2]), .Y(n232) );
  AND3X1_RVT U414 ( .A1(a3stg_id[3]), .A2(a3stg_id[4]), .A3(n232), .Y(n262) );
  INVX1_RVT U415 ( .A(a3stg_id[3]), .Y(n234) );
  AND3X1_RVT U416 ( .A1(a3stg_id[4]), .A2(n234), .A3(n232), .Y(n261) );
  INVX1_RVT U417 ( .A(a3stg_id[4]), .Y(n233) );
  AND3X1_RVT U418 ( .A1(a3stg_id[3]), .A2(n233), .A3(n232), .Y(n260) );
  AND3X1_RVT U419 ( .A1(n233), .A2(n234), .A3(n232), .Y(n259) );
  AND3X1_RVT U420 ( .A1(a3stg_id[2]), .A2(n233), .A3(n234), .Y(n258) );
  AND3X1_RVT U421 ( .A1(a3stg_id[3]), .A2(a3stg_id[2]), .A3(n233), .Y(n257) );
  AND3X1_RVT U422 ( .A1(a3stg_id[4]), .A2(a3stg_id[2]), .A3(n234), .Y(n256) );
  NOR4X1_RVT U423 ( .A1(a3stg_exp[9]), .A2(a3stg_exp[6]), .A3(a3stg_exp[4]), 
        .A4(a3stg_exp[5]), .Y(n238) );
  NOR4X1_RVT U424 ( .A1(a3stg_exp[7]), .A2(a3stg_exp[10]), .A3(a3stg_exp[8]), 
        .A4(a3stg_exp[3]), .Y(n237) );
  AND4X1_RVT U425 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .Y(
        a3stg_exp10_1_eq0) );
  INVX1_RVT U426 ( .A(a3stg_exp[0]), .Y(n239) );
  AND2X1_RVT U427 ( .A1(a3stg_exp10_1_eq0), .A2(n239), .Y(a3stg_exp10_0_eq0)
         );
  AOI21X1_RVT U428 ( .A1(a3stg_exp10_0_eq0), .A2(a3stg_faddsubop), .A3(
        a3stg_fsdtoix), .Y(a4stg_rnd_frac_add_inv) );
  NAND2X0_RVT U429 ( .A1(a1stg_expadd1[5]), .A2(n240), .Y(n247) );
  OA22X1_RVT U430 ( .A1(a1stg_expadd2[5]), .A2(n243), .A3(a1stg_expadd4_inv[5]), .A4(n241), .Y(n246) );
  NAND3X0_RVT U431 ( .A1(n247), .A2(n246), .A3(n245), .Y(a2stg_shr_cnt_in[5])
         );
  INVX0_RVT U432 ( .A(a2stg_shr_cnt_in[5]), .Y(a2stg_shr_cnt_5_inv_in) );
  NAND2X0_RVT U433 ( .A1(n249), .A2(n248), .Y(n244) );
endmodule


module clken_buf_11 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_0 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_14 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_14 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_13 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_13 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_12 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_12 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_0 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, net24246, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N4), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N4), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_15 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, net24246, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_15 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N4), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N4), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_14 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, net24246, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_14 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N4), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N4), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N4), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N4), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N4), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_13 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, net24246, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_13 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N4), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N4), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N4), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N4), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N4), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE4_3 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N4, net24462, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_3 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24462), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24462), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24462), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24462), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24462), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_11 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_11 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_10 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_10 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE12 ( din, en, clk, q, se, si, so );
  input [11:0] din;
  output [11:0] q;
  input [11:0] si;
  output [11:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, net24552, n3,
         n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE12 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24552), .TE(1'b0) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24552), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24552), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24552), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24552), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24552), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24552), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24552), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24552), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24552), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24552), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24552), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24552), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  OR2X1_RVT U16 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_12 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, net24246, n1,
         n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_12 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  OR2X1_RVT U16 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_11 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N9, N10, N11, N12, N14, net24246, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_11 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N10), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N10), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U5 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U6 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U7 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U8 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U10 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_10 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, net24246, n1,
         n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_10 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  OR2X1_RVT U16 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dff_SIZE13_0 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1, n2;

  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[11]), .A2(n2), .Y(N14) );
endmodule


module dff_SIZE13_6 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1;

  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
endmodule


module dff_SIZE13_5 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1;

  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
endmodule


module dff_SIZE13_4 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1;

  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_9 ( din, en, clk, se, si, so, \q[12] , \q[11] , \q[10] , 
        \q[9] , \q[8] , \q[7] , \q[6]_BAR , \q[0] , \q[5]_BAR , \q[4]_BAR , 
        \q[3]_BAR , \q[2]_BAR , \q[1]_BAR  );
  input [12:0] din;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  output \q[12] , \q[11] , \q[10] , \q[9] , \q[8] , \q[7] , \q[6]_BAR , \q[0] ,
         \q[5]_BAR , \q[4]_BAR , \q[3]_BAR , \q[2]_BAR , \q[1]_BAR ;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, net24246, n8,
         n9;
  wire   [12:0] q;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_9 clk_gate_q_reg ( .CLK(clk), .EN(n9), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .QN(\q[6]_BAR ) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .QN(\q[5]_BAR ) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .QN(\q[4]_BAR ) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .QN(\q[3]_BAR ) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .QN(\q[2]_BAR ) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .QN(\q[1]_BAR ) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n8) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n8), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n8), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n8), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n8), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n8), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n8), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n8), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n8), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n8), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n8), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n8), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n8), .Y(N15) );
  OR2X1_RVT U16 ( .A1(se), .A2(en), .Y(n9) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_9 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_9 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_8 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_8 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_7 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_7 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_6 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_6 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N4), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N4), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N4), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N4), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N4), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module fpu_add_exp_dp ( inq_in1, inq_in2, inq_op, inq_op_7, a1stg_step, 
        a1stg_faddsubd, a1stg_faddsubs, a1stg_fsdtoix, a6stg_step, a1stg_fstod, 
        a1stg_fdtos, a1stg_fstoi, a1stg_fstox, a1stg_fdtoi, a1stg_fdtox, 
        a2stg_fsdtoix_fdtos, a2stg_faddsubop, a2stg_fitos, a2stg_fitod, 
        a2stg_fxtos, a2stg_fxtod, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add, 
        a3stg_inc_exp_inv, a3stg_same_exp_inv, a3stg_dec_exp_inv, 
        a3stg_faddsubop, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, 
        a4stg_shl_cnt, a4stg_denorm_inv, a4stg_rndadd_cout, add_exp_out_expinc, 
        add_exp_out_exp, add_exp_out_exp1, a4stg_in_of, add_exp_out_expadd, 
        a4stg_dblop, a4stg_to_0_inv, fadd_clken_l, rclk, a1stg_expadd3_11, 
        a1stg_expadd1_11_0, a1stg_expadd4_inv, a1stg_expadd2_5_0, a2stg_exp, 
        a2stg_expadd, a3stg_exp_10_0, a4stg_exp_11_0, add_exp_out, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [1:0] inq_op;
  input [5:0] a4stg_shl_cnt;
  output [11:0] a1stg_expadd1_11_0;
  output [10:0] a1stg_expadd4_inv;
  output [5:0] a1stg_expadd2_5_0;
  output [11:0] a2stg_exp;
  output [12:0] a2stg_expadd;
  output [10:0] a3stg_exp_10_0;
  output [11:0] a4stg_exp_11_0;
  output [10:0] add_exp_out;
  input inq_op_7, a1stg_step, a1stg_faddsubd, a1stg_faddsubs, a1stg_fsdtoix,
         a6stg_step, a1stg_fstod, a1stg_fdtos, a1stg_fstoi, a1stg_fstox,
         a1stg_fdtoi, a1stg_fdtox, a2stg_fsdtoix_fdtos, a2stg_faddsubop,
         a2stg_fitos, a2stg_fitod, a2stg_fxtos, a2stg_fxtod, a3stg_exp_7ff,
         a3stg_exp_ff, a3stg_exp_add, a3stg_inc_exp_inv, a3stg_same_exp_inv,
         a3stg_dec_exp_inv, a3stg_faddsubop, a3stg_fdtos_inv,
         a4stg_fixtos_fxtod_inv, a4stg_denorm_inv, a4stg_rndadd_cout,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1, a4stg_in_of,
         add_exp_out_expadd, a4stg_dblop, a4stg_to_0_inv, fadd_clken_l, rclk,
         se, si;
  output a1stg_expadd3_11, so;
  wire   clk, a1stg_op_7_0, \a3stg_exp[11] , N346, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, \intadd_3/CI ,
         \intadd_3/SUM[4] , \intadd_3/SUM[3] , \intadd_3/SUM[2] ,
         \intadd_3/SUM[1] , \intadd_3/SUM[0] , \intadd_3/n5 , \intadd_3/n4 ,
         \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 , \intadd_0/n12 ,
         \intadd_0/n11 , \intadd_0/n10 , \intadd_0/n9 , \intadd_0/n8 ,
         \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/A[8] ,
         \intadd_1/A[7] , \intadd_1/A[6] , \intadd_1/A[5] , \intadd_1/A[4] ,
         \intadd_1/A[3] , \intadd_1/A[2] , \intadd_1/A[1] , \intadd_1/A[0] ,
         \intadd_1/B[8] , \intadd_1/B[7] , \intadd_1/B[6] , \intadd_1/B[5] ,
         \intadd_1/B[4] , \intadd_1/B[3] , \intadd_1/B[2] , \intadd_1/B[1] ,
         \intadd_1/B[0] , \intadd_1/CI , \intadd_1/SUM[9] , \intadd_1/SUM[8] ,
         \intadd_1/SUM[7] , \intadd_1/SUM[6] , \intadd_1/SUM[5] ,
         \intadd_1/SUM[4] , \intadd_1/SUM[3] , \intadd_1/SUM[2] ,
         \intadd_1/SUM[1] , \intadd_1/SUM[0] , \intadd_1/n10 , \intadd_1/n9 ,
         \intadd_1/n8 , \intadd_1/n7 , \intadd_1/n6 , \intadd_1/n5 ,
         \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 , \intadd_2/A[9] ,
         \intadd_2/A[8] , \intadd_2/A[7] , \intadd_2/A[6] , \intadd_2/A[5] ,
         \intadd_2/A[4] , \intadd_2/A[3] , \intadd_2/A[2] , \intadd_2/A[1] ,
         \intadd_2/A[0] , \intadd_2/B[9] , \intadd_2/B[8] , \intadd_2/B[7] ,
         \intadd_2/B[6] , \intadd_2/B[5] , \intadd_2/B[4] , \intadd_2/B[3] ,
         \intadd_2/B[2] , \intadd_2/B[1] , \intadd_2/B[0] , \intadd_2/CI ,
         \intadd_2/SUM[9] , \intadd_2/SUM[8] , \intadd_2/SUM[7] ,
         \intadd_2/SUM[6] , \intadd_2/SUM[5] , \intadd_2/SUM[4] ,
         \intadd_2/SUM[3] , \intadd_2/SUM[2] , \intadd_2/SUM[1] ,
         \intadd_2/SUM[0] , \intadd_2/n10 , \intadd_2/n9 , \intadd_2/n8 ,
         \intadd_2/n7 , \intadd_2/n6 , \intadd_2/n5 , \intadd_2/n4 ,
         \intadd_2/n3 , \intadd_2/n2 , \intadd_2/n1 , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n334;
  wire   [62:52] a1stg_in1;
  wire   [62:52] a1stg_in1a;
  wire   [62:52] a1stg_in2;
  wire   [62:52] a1stg_in2a;
  wire   [12:0] a1stg_dp_sngop;
  wire   [12:0] a1stg_dp_sngopa;
  wire   [12:0] a1stg_dp_dblop;
  wire   [12:0] a1stg_dp_dblopa;
  wire   [9:7] a1stg_op_7;
  wire   [10:0] a1stg_expadd3_in1;
  wire   [10:0] a1stg_expadd3_in2;
  wire   [12:0] a2stg_exp_in;
  wire   [12:0] a2stg_expa;
  wire   [12:5] a2stg_expadd_in2_in;
  wire   [12:0] a2stg_expadd_in2;
  wire   [12:0] a3stg_exp_in;
  wire   [12:0] a4stg_exp_pre1_in;
  wire   [12:0] a4stg_exp_pre1;
  wire   [12:0] a4stg_exp_pre3_in;
  wire   [12:0] a4stg_exp_pre3;
  wire   [12:0] a4stg_exp_pre2_in;
  wire   [12:0] a4stg_exp_pre2;
  wire   [12:0] a4stg_exp_pre4_in;
  wire   [12:0] a4stg_exp_pre4;
  wire   [12:0] a4stg_exp2;
  wire   [10:0] add_exp_out1;
  wire   [10:0] add_exp_out2;
  wire   [10:0] add_exp_out3;
  wire   [10:0] add_exp_out4;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19;
  assign a1stg_expadd4_inv[10] = \intadd_1/SUM[9] ;
  assign a1stg_expadd4_inv[9] = \intadd_1/SUM[8] ;
  assign a1stg_expadd4_inv[8] = \intadd_1/SUM[7] ;
  assign a1stg_expadd4_inv[7] = \intadd_1/SUM[6] ;
  assign a1stg_expadd4_inv[6] = \intadd_1/SUM[5] ;
  assign a1stg_expadd4_inv[5] = \intadd_1/SUM[4] ;
  assign a1stg_expadd4_inv[4] = \intadd_1/SUM[3] ;
  assign a1stg_expadd4_inv[3] = \intadd_1/SUM[2] ;
  assign a1stg_expadd4_inv[2] = \intadd_1/SUM[1] ;
  assign a1stg_expadd4_inv[1] = \intadd_1/SUM[0] ;
  assign a1stg_expadd1_11_0[11] = \intadd_2/n1 ;
  assign so = 1'b0;

  clken_buf_11 ckbuf_add_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fadd_clken_l), 
        .tmb_l(n334) );
  dffe_SIZE11_0 i_a1stg_in1 ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_14 i_a1stg_in1a ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1a), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_13 i_a1stg_in2 ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_12 i_a1stg_in2a ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2a), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_0 i_a1stg_dp_sngop ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0]}), .en(a1stg_step), .clk(clk), .q({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, a1stg_dp_sngop[7:0]}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_15 i_a1stg_dp_sngopa ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0]}), .en(a1stg_step), .clk(clk), .q({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, a1stg_dp_sngopa[7:0]}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_14 i_a1stg_dp_dblop ( .din({1'b0, 1'b0, inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1]}), .en(a1stg_step), .clk(clk), .q({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        a1stg_dp_dblop[10:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_13 i_a1stg_dp_dblopa ( .din({1'b0, 1'b0, inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1]}), .en(a1stg_step), .clk(clk), .q({
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        a1stg_dp_dblopa[10:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE4_3 i_a1stg_op_7 ( .din({1'b0, 1'b0, 1'b0, inq_op_7}), .en(
        a1stg_step), .clk(clk), .q({a1stg_op_7, a1stg_op_7_0}), .se(se), .si({
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_11 i_a1stg_expadd3_in1 ( .din(inq_in1), .en(a1stg_step), .clk(
        clk), .q(a1stg_expadd3_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_10 i_a1stg_expadd3_in2 ( .din({n157, n158, n159, n160, n161, 
        n162, n163, n164, n165, n166, n167}), .en(a1stg_step), .clk(clk), .q(
        a1stg_expadd3_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE12 i_a2stg_exp ( .din(a2stg_exp_in[11:0]), .en(a6stg_step), .clk(
        clk), .q(a2stg_exp), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_12 i_a2stg_expa ( .din({1'b0, a2stg_exp_in[11:0]}), .en(
        a6stg_step), .clk(clk), .q({SYNOPSYS_UNCONNECTED__14, a2stg_expa[11:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_11 i_a2stg_expadd2_in2 ( .din({1'b0, 1'b0, 
        a2stg_expadd_in2_in[10], 1'b0, a2stg_expadd_in2_in[8:5], 1'b0, 1'b0, 
        1'b0, 1'b0, a1stg_fdtos}), .en(a6stg_step), .clk(clk), .q(
        a2stg_expadd_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_10 i_a3stg_exp ( .din({1'b0, N346, a3stg_exp_in[10:0]}), .en(
        a6stg_step), .clk(clk), .q({SYNOPSYS_UNCONNECTED__15, \a3stg_exp[11] , 
        a3stg_exp_10_0}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE13_0 i_a4stg_exp_pre1 ( .din({1'b0, a4stg_exp_pre1_in[11:0]}), .clk(
        clk), .q({SYNOPSYS_UNCONNECTED__16, a4stg_exp_pre1[11:0]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dff_SIZE13_6 i_a4stg_exp_pre3 ( .din({1'b0, a4stg_exp_pre3_in[11:0]}), .clk(
        clk), .q({SYNOPSYS_UNCONNECTED__17, a4stg_exp_pre3[11:0]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dff_SIZE13_5 i_a4stg_exp_pre2 ( .din({1'b0, a4stg_exp_pre2_in[11:0]}), .clk(
        clk), .q({SYNOPSYS_UNCONNECTED__18, a4stg_exp_pre2[11:0]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dff_SIZE13_4 i_a4stg_exp_pre4 ( .din({1'b0, a4stg_exp_pre4_in[11:0]}), .clk(
        clk), .q({SYNOPSYS_UNCONNECTED__19, a4stg_exp_pre4[11:0]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dffe_SIZE13_9 i_a4stg_exp2 ( .din({1'b0, \a3stg_exp[11] , a3stg_exp_10_0}), 
        .en(a6stg_step), .clk(clk), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\q[11] (
        a4stg_exp2[11]), .\q[10] (a4stg_exp2[10]), .\q[9] (a4stg_exp2[9]), 
        .\q[8] (a4stg_exp2[8]), .\q[7] (a4stg_exp2[7]), .\q[6]_BAR (
        a4stg_exp2[6]), .\q[0] (a4stg_exp2[0]), .\q[5]_BAR (a4stg_exp2[5]), 
        .\q[4]_BAR (a4stg_exp2[4]), .\q[3]_BAR (a4stg_exp2[3]), .\q[2]_BAR (
        a4stg_exp2[2]), .\q[1]_BAR (a4stg_exp2[1]) );
  dffe_SIZE11_9 i_add_exp_out1 ( .din({n145, n143, n141, n139, n137, n135, 
        n133, n131, n129, n127, n125}), .en(a6stg_step), .clk(clk), .q(
        add_exp_out1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_8 i_add_exp_out2 ( .din({n113, n114, n115, n116, n117, n118, 
        n119, n120, n121, n122, n123}), .en(a6stg_step), .clk(clk), .q(
        add_exp_out2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_7 i_add_exp_out3 ( .din({n144, n142, n140, n138, n136, n134, 
        n132, n130, n128, n126, n124}), .en(a6stg_step), .clk(clk), .q(
        add_exp_out3), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_6 i_add_exp_out4 ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, a4stg_rndadd_cout}), .en(a6stg_step), .clk(clk), .q(add_exp_out4), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  FADDX1_RVT \intadd_3/U6  ( .A(a4stg_exp2[1]), .B(a4stg_shl_cnt[1]), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n5 ), .S(\intadd_3/SUM[0] ) );
  FADDX1_RVT \intadd_3/U5  ( .A(a4stg_exp2[2]), .B(a4stg_shl_cnt[2]), .CI(
        \intadd_3/n5 ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[1] ) );
  FADDX1_RVT \intadd_3/U4  ( .A(a4stg_exp2[3]), .B(a4stg_shl_cnt[3]), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[2] ) );
  FADDX1_RVT \intadd_3/U3  ( .A(a4stg_exp2[4]), .B(a4stg_shl_cnt[4]), .CI(
        \intadd_3/n3 ), .CO(\intadd_3/n2 ), .S(\intadd_3/SUM[3] ) );
  FADDX1_RVT \intadd_3/U2  ( .A(a4stg_exp2[5]), .B(a4stg_shl_cnt[5]), .CI(
        \intadd_3/n2 ), .CO(\intadd_3/n1 ), .S(\intadd_3/SUM[4] ) );
  FADDX1_RVT \intadd_0/U13  ( .A(a2stg_expadd_in2[0]), .B(a2stg_fsdtoix_fdtos), 
        .CI(a2stg_expa[0]), .CO(\intadd_0/n12 ), .S(a2stg_expadd[0]) );
  FADDX1_RVT \intadd_0/U12  ( .A(a2stg_expa[1]), .B(a2stg_expadd_in2[1]), .CI(
        \intadd_0/n12 ), .CO(\intadd_0/n11 ), .S(a2stg_expadd[1]) );
  FADDX1_RVT \intadd_0/U11  ( .A(a2stg_expa[2]), .B(a2stg_expadd_in2[2]), .CI(
        \intadd_0/n11 ), .CO(\intadd_0/n10 ), .S(a2stg_expadd[2]) );
  FADDX1_RVT \intadd_0/U10  ( .A(a2stg_expa[3]), .B(a2stg_expadd_in2[3]), .CI(
        \intadd_0/n10 ), .CO(\intadd_0/n9 ), .S(a2stg_expadd[3]) );
  FADDX1_RVT \intadd_0/U9  ( .A(a2stg_expa[4]), .B(a2stg_expadd_in2[4]), .CI(
        \intadd_0/n9 ), .CO(\intadd_0/n8 ), .S(a2stg_expadd[4]) );
  FADDX1_RVT \intadd_0/U8  ( .A(a2stg_expa[5]), .B(a2stg_expadd_in2[5]), .CI(
        \intadd_0/n8 ), .CO(\intadd_0/n7 ), .S(a2stg_expadd[5]) );
  FADDX1_RVT \intadd_0/U7  ( .A(a2stg_expa[6]), .B(a2stg_expadd_in2[6]), .CI(
        \intadd_0/n7 ), .CO(\intadd_0/n6 ), .S(a2stg_expadd[6]) );
  FADDX1_RVT \intadd_0/U6  ( .A(a2stg_expa[7]), .B(a2stg_expadd_in2[7]), .CI(
        \intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(a2stg_expadd[7]) );
  FADDX1_RVT \intadd_0/U5  ( .A(a2stg_expa[8]), .B(a2stg_expadd_in2[8]), .CI(
        \intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(a2stg_expadd[8]) );
  FADDX1_RVT \intadd_0/U4  ( .A(a2stg_expa[9]), .B(a2stg_expadd_in2[9]), .CI(
        \intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(a2stg_expadd[9]) );
  FADDX1_RVT \intadd_0/U3  ( .A(a2stg_expa[10]), .B(a2stg_expadd_in2[10]), 
        .CI(\intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(a2stg_expadd[10]) );
  FADDX1_RVT \intadd_0/U2  ( .A(a2stg_expa[11]), .B(a2stg_expadd_in2[11]), 
        .CI(\intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(a2stg_expadd[11]) );
  FADDX1_RVT \intadd_1/U11  ( .A(\intadd_1/B[0] ), .B(\intadd_1/A[0] ), .CI(
        \intadd_1/CI ), .CO(\intadd_1/n10 ), .S(\intadd_1/SUM[0] ) );
  FADDX1_RVT \intadd_1/U10  ( .A(\intadd_1/B[1] ), .B(\intadd_1/A[1] ), .CI(
        \intadd_1/n10 ), .CO(\intadd_1/n9 ), .S(\intadd_1/SUM[1] ) );
  FADDX1_RVT \intadd_1/U9  ( .A(\intadd_1/B[2] ), .B(\intadd_1/A[2] ), .CI(
        \intadd_1/n9 ), .CO(\intadd_1/n8 ), .S(\intadd_1/SUM[2] ) );
  FADDX1_RVT \intadd_1/U8  ( .A(\intadd_1/B[3] ), .B(\intadd_1/A[3] ), .CI(
        \intadd_1/n8 ), .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[3] ) );
  FADDX1_RVT \intadd_1/U7  ( .A(\intadd_1/B[4] ), .B(\intadd_1/A[4] ), .CI(
        \intadd_1/n7 ), .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[4] ) );
  FADDX1_RVT \intadd_1/U6  ( .A(\intadd_1/B[5] ), .B(\intadd_1/A[5] ), .CI(
        \intadd_1/n6 ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[5] ) );
  FADDX1_RVT \intadd_1/U5  ( .A(\intadd_1/B[6] ), .B(\intadd_1/A[6] ), .CI(
        \intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[6] ) );
  FADDX1_RVT \intadd_1/U4  ( .A(\intadd_1/B[7] ), .B(\intadd_1/A[7] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[7] ) );
  FADDX1_RVT \intadd_1/U3  ( .A(\intadd_1/B[8] ), .B(\intadd_1/A[8] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[8] ) );
  FADDX1_RVT \intadd_2/U11  ( .A(\intadd_2/B[0] ), .B(\intadd_2/A[0] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n10 ), .S(\intadd_2/SUM[0] ) );
  FADDX1_RVT \intadd_2/U10  ( .A(\intadd_2/B[1] ), .B(\intadd_2/A[1] ), .CI(
        \intadd_2/n10 ), .CO(\intadd_2/n9 ), .S(\intadd_2/SUM[1] ) );
  FADDX1_RVT \intadd_2/U9  ( .A(\intadd_2/B[2] ), .B(\intadd_2/A[2] ), .CI(
        \intadd_2/n9 ), .CO(\intadd_2/n8 ), .S(\intadd_2/SUM[2] ) );
  FADDX1_RVT \intadd_2/U8  ( .A(\intadd_2/B[3] ), .B(\intadd_2/A[3] ), .CI(
        \intadd_2/n8 ), .CO(\intadd_2/n7 ), .S(\intadd_2/SUM[3] ) );
  FADDX1_RVT \intadd_2/U7  ( .A(\intadd_2/B[4] ), .B(\intadd_2/A[4] ), .CI(
        \intadd_2/n7 ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[4] ) );
  FADDX1_RVT \intadd_2/U6  ( .A(\intadd_2/B[5] ), .B(\intadd_2/A[5] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[5] ) );
  FADDX1_RVT \intadd_2/U5  ( .A(\intadd_2/B[6] ), .B(\intadd_2/A[6] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[6] ) );
  FADDX1_RVT \intadd_2/U4  ( .A(\intadd_2/B[7] ), .B(\intadd_2/A[7] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[7] ) );
  FADDX1_RVT \intadd_2/U3  ( .A(\intadd_2/B[8] ), .B(\intadd_2/A[8] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[8] ) );
  FADDX1_RVT \intadd_2/U2  ( .A(\intadd_2/B[9] ), .B(\intadd_2/A[9] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[9] ) );
  INVX0_RVT U3 ( .A(n238), .Y(n239) );
  INVX0_RVT U4 ( .A(n308), .Y(n307) );
  INVX0_RVT U5 ( .A(\intadd_2/n1 ), .Y(n29) );
  INVX0_RVT U6 ( .A(n147), .Y(n146) );
  INVX0_RVT U7 ( .A(n13), .Y(n8) );
  INVX0_RVT U8 ( .A(n109), .Y(n108) );
  INVX0_RVT U9 ( .A(n172), .Y(n156) );
  INVX0_RVT U10 ( .A(n168), .Y(n151) );
  INVX0_RVT U11 ( .A(n16), .Y(n7) );
  INVX0_RVT U12 ( .A(n152), .Y(n70) );
  INVX0_RVT U13 ( .A(n220), .Y(n208) );
  INVX0_RVT U14 ( .A(n104), .Y(n103) );
  INVX0_RVT U15 ( .A(inq_in2[55]), .Y(n164) );
  INVX0_RVT U16 ( .A(inq_in2[56]), .Y(n163) );
  INVX0_RVT U17 ( .A(inq_in2[58]), .Y(n161) );
  INVX0_RVT U18 ( .A(inq_in2[61]), .Y(n158) );
  INVX0_RVT U19 ( .A(inq_in2[57]), .Y(n162) );
  INVX0_RVT U20 ( .A(inq_in2[59]), .Y(n160) );
  INVX0_RVT U21 ( .A(inq_in2[60]), .Y(n159) );
  INVX0_RVT U22 ( .A(inq_in2[62]), .Y(n157) );
  INVX0_RVT U23 ( .A(n19), .Y(n6) );
  OR3X1_RVT U24 ( .A1(a2stg_fxtod), .A2(a2stg_fxtos), .A3(n237), .Y(n229) );
  INVX0_RVT U25 ( .A(n99), .Y(n98) );
  INVX0_RVT U26 ( .A(n22), .Y(n5) );
  INVX0_RVT U27 ( .A(n250), .Y(n251) );
  INVX0_RVT U28 ( .A(n94), .Y(n93) );
  OR3X1_RVT U29 ( .A1(a1stg_fstoi), .A2(a1stg_fstox), .A3(
        a2stg_expadd_in2_in[7]), .Y(a2stg_expadd_in2_in[8]) );
  INVX0_RVT U30 ( .A(n25), .Y(n4) );
  OR3X1_RVT U31 ( .A1(a1stg_fdtoi), .A2(a1stg_fdtox), .A3(
        a2stg_expadd_in2_in[10]), .Y(a2stg_expadd_in2_in[6]) );
  OR3X1_RVT U32 ( .A1(a1stg_fstod), .A2(a1stg_fdtoi), .A3(a1stg_fdtox), .Y(
        a2stg_expadd_in2_in[7]) );
  INVX0_RVT U33 ( .A(n89), .Y(n88) );
  INVX0_RVT U34 ( .A(a1stg_fsdtoix), .Y(n209) );
  OR3X1_RVT U35 ( .A1(a1stg_fdtos), .A2(a1stg_fstoi), .A3(a1stg_fstox), .Y(
        a2stg_expadd_in2_in[10]) );
  OR3X1_RVT U36 ( .A1(a1stg_fdtos), .A2(a1stg_fstoi), .A3(a1stg_fdtoi), .Y(
        a2stg_expadd_in2_in[5]) );
  OR3X1_RVT U37 ( .A1(\intadd_1/A[1] ), .A2(a1stg_expadd2_5_0[0]), .A3(
        \intadd_1/A[0] ), .Y(n40) );
  INVX0_RVT U38 ( .A(n28), .Y(n3) );
  INVX0_RVT U39 ( .A(n261), .Y(n262) );
  INVX0_RVT U40 ( .A(n260), .Y(n263) );
  INVX0_RVT U41 ( .A(n84), .Y(n83) );
  INVX0_RVT U42 ( .A(n210), .Y(n178) );
  INVX0_RVT U43 ( .A(a4stg_shl_cnt[0]), .Y(n280) );
  INVX0_RVT U44 ( .A(\a3stg_exp[11] ), .Y(n242) );
  INVX0_RVT U45 ( .A(a3stg_exp_10_0[2]), .Y(n76) );
  INVX0_RVT U46 ( .A(a3stg_exp_10_0[3]), .Y(n80) );
  INVX0_RVT U47 ( .A(a3stg_exp_10_0[4]), .Y(n85) );
  INVX0_RVT U48 ( .A(a3stg_exp_10_0[5]), .Y(n90) );
  INVX0_RVT U49 ( .A(a3stg_exp_10_0[6]), .Y(n95) );
  INVX0_RVT U50 ( .A(a3stg_exp_10_0[7]), .Y(n100) );
  INVX0_RVT U51 ( .A(a3stg_exp_10_0[8]), .Y(n105) );
  INVX0_RVT U52 ( .A(a3stg_exp_10_0[9]), .Y(n110) );
  INVX0_RVT U53 ( .A(a3stg_exp_10_0[10]), .Y(n148) );
  INVX1_RVT U54 ( .A(a4stg_fixtos_fxtod_inv), .Y(n266) );
  AOI22X1_RVT U55 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[0]), .A3(
        a1stg_in2[55]), .A4(n200), .Y(n1) );
  XOR2X1_RVT U56 ( .A1(\intadd_0/n1 ), .A2(a2stg_expadd_in2[12]), .Y(
        a2stg_expadd[12]) );
  INVX1_RVT U57 ( .A(a6stg_step), .Y(n282) );
  NOR4X1_RVT U58 ( .A1(a4stg_exp_pre1[0]), .A2(a4stg_exp_pre2[0]), .A3(
        a4stg_exp_pre3[0]), .A4(a4stg_exp_pre4[0]), .Y(n300) );
  INVX1_RVT U59 ( .A(n300), .Y(a4stg_exp_11_0[0]) );
  NOR4X1_RVT U60 ( .A1(a4stg_exp_pre1[1]), .A2(a4stg_exp_pre2[1]), .A3(
        a4stg_exp_pre3[1]), .A4(a4stg_exp_pre4[1]), .Y(n299) );
  INVX1_RVT U61 ( .A(n299), .Y(a4stg_exp_11_0[1]) );
  AOI22X1_RVT U62 ( .A1(a1stg_in2a[55]), .A2(a1stg_dp_sngopa[0]), .A3(
        a1stg_dp_dblopa[0]), .A4(a1stg_in2a[52]), .Y(a1stg_expadd2_5_0[0]) );
  NOR4X1_RVT U63 ( .A1(a4stg_exp_pre1[2]), .A2(a4stg_exp_pre2[2]), .A3(
        a4stg_exp_pre3[2]), .A4(a4stg_exp_pre4[2]), .Y(n302) );
  INVX1_RVT U64 ( .A(n302), .Y(a4stg_exp_11_0[2]) );
  NOR4X1_RVT U65 ( .A1(a4stg_exp_pre1[7]), .A2(a4stg_exp_pre2[7]), .A3(
        a4stg_exp_pre3[7]), .A4(a4stg_exp_pre4[7]), .Y(n14) );
  INVX1_RVT U66 ( .A(n14), .Y(a4stg_exp_11_0[7]) );
  NOR4X1_RVT U67 ( .A1(a4stg_exp_pre1[4]), .A2(a4stg_exp_pre2[4]), .A3(
        a4stg_exp_pre3[4]), .A4(a4stg_exp_pre4[4]), .Y(n23) );
  INVX1_RVT U68 ( .A(n23), .Y(a4stg_exp_11_0[4]) );
  NOR4X1_RVT U69 ( .A1(a4stg_exp_pre1[3]), .A2(a4stg_exp_pre2[3]), .A3(
        a4stg_exp_pre3[3]), .A4(a4stg_exp_pre4[3]), .Y(n26) );
  INVX1_RVT U70 ( .A(n26), .Y(a4stg_exp_11_0[3]) );
  NOR4X1_RVT U71 ( .A1(a4stg_exp_pre1[6]), .A2(a4stg_exp_pre2[6]), .A3(
        a4stg_exp_pre3[6]), .A4(a4stg_exp_pre4[6]), .Y(n17) );
  INVX1_RVT U72 ( .A(n17), .Y(a4stg_exp_11_0[6]) );
  NOR4X1_RVT U73 ( .A1(a4stg_exp_pre1[5]), .A2(a4stg_exp_pre2[5]), .A3(
        a4stg_exp_pre3[5]), .A4(a4stg_exp_pre4[5]), .Y(n20) );
  INVX1_RVT U74 ( .A(n20), .Y(a4stg_exp_11_0[5]) );
  NOR4X1_RVT U75 ( .A1(a4stg_exp_pre1[10]), .A2(a4stg_exp_pre2[10]), .A3(
        a4stg_exp_pre3[10]), .A4(a4stg_exp_pre4[10]), .Y(n309) );
  INVX1_RVT U76 ( .A(n309), .Y(a4stg_exp_11_0[10]) );
  NOR4X1_RVT U77 ( .A1(a4stg_exp_pre1[9]), .A2(a4stg_exp_pre2[9]), .A3(
        a4stg_exp_pre3[9]), .A4(a4stg_exp_pre4[9]), .Y(n9) );
  INVX1_RVT U78 ( .A(n9), .Y(a4stg_exp_11_0[9]) );
  NOR4X1_RVT U79 ( .A1(a4stg_exp_pre1[8]), .A2(a4stg_exp_pre2[8]), .A3(
        a4stg_exp_pre3[8]), .A4(a4stg_exp_pre4[8]), .Y(n11) );
  INVX1_RVT U80 ( .A(n11), .Y(a4stg_exp_11_0[8]) );
  AOI22X1_RVT U81 ( .A1(a1stg_in2a[56]), .A2(a1stg_dp_sngopa[1]), .A3(
        a1stg_dp_dblopa[1]), .A4(a1stg_in2a[53]), .Y(\intadd_1/A[0] ) );
  AOI22X1_RVT U82 ( .A1(a1stg_in2a[60]), .A2(a1stg_dp_sngopa[5]), .A3(
        a1stg_dp_dblopa[5]), .A4(a1stg_in2a[57]), .Y(\intadd_1/A[4] ) );
  INVX1_RVT U83 ( .A(se), .Y(n334) );
  NOR2X0_RVT U84 ( .A1(a1stg_expadd2_5_0[0]), .A2(\intadd_1/A[0] ), .Y(n36) );
  AOI21X1_RVT U85 ( .A1(\intadd_1/A[0] ), .A2(a1stg_expadd2_5_0[0]), .A3(n36), 
        .Y(a1stg_expadd2_5_0[1]) );
  INVX1_RVT U86 ( .A(\intadd_2/SUM[0] ), .Y(a1stg_expadd1_11_0[1]) );
  INVX1_RVT U87 ( .A(\intadd_2/SUM[1] ), .Y(a1stg_expadd1_11_0[2]) );
  INVX1_RVT U88 ( .A(\intadd_2/SUM[3] ), .Y(a1stg_expadd1_11_0[4]) );
  AO22X1_RVT U89 ( .A1(a1stg_in2a[57]), .A2(a1stg_dp_sngopa[2]), .A3(
        a1stg_dp_dblopa[2]), .A4(a1stg_in2a[54]), .Y(n35) );
  INVX1_RVT U90 ( .A(n35), .Y(\intadd_1/A[1] ) );
  INVX1_RVT U91 ( .A(\intadd_2/SUM[2] ), .Y(a1stg_expadd1_11_0[3]) );
  INVX1_RVT U92 ( .A(\intadd_2/SUM[9] ), .Y(a1stg_expadd1_11_0[10]) );
  INVX1_RVT U93 ( .A(\intadd_2/SUM[5] ), .Y(a1stg_expadd1_11_0[6]) );
  INVX1_RVT U94 ( .A(\intadd_2/SUM[8] ), .Y(a1stg_expadd1_11_0[9]) );
  INVX1_RVT U95 ( .A(\intadd_2/SUM[6] ), .Y(a1stg_expadd1_11_0[7]) );
  INVX1_RVT U96 ( .A(\intadd_2/SUM[7] ), .Y(a1stg_expadd1_11_0[8]) );
  AO22X1_RVT U97 ( .A1(a1stg_in1a[55]), .A2(a1stg_dp_sngop[0]), .A3(
        a1stg_dp_dblop[0]), .A4(a1stg_in1a[52]), .Y(n311) );
  NAND2X0_RVT U98 ( .A1(a1stg_expadd2_5_0[0]), .A2(n311), .Y(n310) );
  INVX1_RVT U99 ( .A(n310), .Y(\intadd_1/B[0] ) );
  AO22X1_RVT U100 ( .A1(a1stg_in2a[59]), .A2(a1stg_dp_sngopa[4]), .A3(
        a1stg_dp_dblopa[4]), .A4(a1stg_in2a[56]), .Y(n44) );
  INVX1_RVT U101 ( .A(n44), .Y(\intadd_1/A[3] ) );
  INVX1_RVT U102 ( .A(\intadd_2/SUM[4] ), .Y(a1stg_expadd1_11_0[5]) );
  AO22X1_RVT U103 ( .A1(a1stg_dp_sngopa[0]), .A2(a1stg_in1[55]), .A3(
        a1stg_dp_dblopa[0]), .A4(a1stg_in1[52]), .Y(n2) );
  NOR2X0_RVT U104 ( .A1(a1stg_op_7_0), .A2(n2), .Y(n193) );
  AO22X1_RVT U105 ( .A1(a1stg_in2[55]), .A2(a1stg_dp_sngop[0]), .A3(
        a1stg_dp_dblop[0]), .A4(a1stg_in2[52]), .Y(n192) );
  NAND2X0_RVT U106 ( .A1(n193), .A2(n192), .Y(n191) );
  INVX1_RVT U107 ( .A(n191), .Y(\intadd_2/B[0] ) );
  NAND2X0_RVT U130 ( .A1(a4stg_rndadd_cout), .A2(add_exp_out_expinc), .Y(n306)
         );
  NAND4X0_RVT U131 ( .A1(a4stg_exp_11_0[3]), .A2(a4stg_exp_11_0[2]), .A3(
        a4stg_exp_11_0[0]), .A4(a4stg_exp_11_0[1]), .Y(n28) );
  NAND2X0_RVT U132 ( .A1(n3), .A2(a4stg_exp_11_0[4]), .Y(n25) );
  NAND2X0_RVT U133 ( .A1(n4), .A2(a4stg_exp_11_0[5]), .Y(n22) );
  NAND2X0_RVT U134 ( .A1(n5), .A2(a4stg_exp_11_0[6]), .Y(n19) );
  NAND2X0_RVT U135 ( .A1(n6), .A2(a4stg_exp_11_0[7]), .Y(n16) );
  NAND2X0_RVT U136 ( .A1(n7), .A2(a4stg_exp_11_0[8]), .Y(n13) );
  NAND2X0_RVT U137 ( .A1(n8), .A2(a4stg_exp_11_0[9]), .Y(n308) );
  NAND2X0_RVT U138 ( .A1(n9), .A2(n13), .Y(n10) );
  NAND3X0_RVT U139 ( .A1(n303), .A2(n308), .A3(n10), .Y(n114) );
  NAND2X0_RVT U140 ( .A1(n11), .A2(n16), .Y(n12) );
  NAND3X0_RVT U141 ( .A1(n303), .A2(n13), .A3(n12), .Y(n115) );
  NAND2X0_RVT U142 ( .A1(n14), .A2(n19), .Y(n15) );
  NAND3X0_RVT U143 ( .A1(n303), .A2(n16), .A3(n15), .Y(n116) );
  INVX1_RVT U144 ( .A(n306), .Y(n303) );
  NAND2X0_RVT U145 ( .A1(n17), .A2(n22), .Y(n18) );
  NAND3X0_RVT U146 ( .A1(n303), .A2(n19), .A3(n18), .Y(n117) );
  NAND2X0_RVT U147 ( .A1(n20), .A2(n25), .Y(n21) );
  NAND3X0_RVT U148 ( .A1(n303), .A2(n22), .A3(n21), .Y(n118) );
  NAND2X0_RVT U149 ( .A1(n23), .A2(n28), .Y(n24) );
  NAND3X0_RVT U150 ( .A1(n303), .A2(n25), .A3(n24), .Y(n119) );
  NAND3X0_RVT U151 ( .A1(a4stg_exp_11_0[2]), .A2(a4stg_exp_11_0[0]), .A3(
        a4stg_exp_11_0[1]), .Y(n304) );
  NAND2X0_RVT U152 ( .A1(n26), .A2(n304), .Y(n27) );
  NAND3X0_RVT U153 ( .A1(n303), .A2(n28), .A3(n27), .Y(n120) );
  AO21X1_RVT U154 ( .A1(\intadd_2/n1 ), .A2(a1stg_faddsubs), .A3(a1stg_fstod), 
        .Y(n200) );
  AND2X1_RVT U155 ( .A1(a1stg_faddsubd), .A2(n29), .Y(n217) );
  AND2X1_RVT U156 ( .A1(a1stg_faddsubs), .A2(n29), .Y(n199) );
  AOI22X1_RVT U157 ( .A1(n217), .A2(a1stg_in1a[52]), .A3(n199), .A4(
        a1stg_in1a[55]), .Y(n31) );
  AO21X1_RVT U158 ( .A1(a1stg_faddsubd), .A2(\intadd_2/n1 ), .A3(a1stg_fdtos), 
        .Y(n216) );
  NAND2X0_RVT U159 ( .A1(a1stg_in2[52]), .A2(n216), .Y(n30) );
  NAND3X0_RVT U160 ( .A1(n1), .A2(n31), .A3(n30), .Y(a2stg_exp_in[0]) );
  AOI22X1_RVT U161 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[1]), .A3(
        a1stg_in2[56]), .A4(n200), .Y(n34) );
  AOI22X1_RVT U162 ( .A1(n217), .A2(a1stg_in1a[53]), .A3(n199), .A4(
        a1stg_in1a[56]), .Y(n33) );
  NAND2X0_RVT U163 ( .A1(a1stg_in2[53]), .A2(n216), .Y(n32) );
  NAND3X0_RVT U164 ( .A1(n34), .A2(n33), .A3(n32), .Y(a2stg_exp_in[1]) );
  OA21X1_RVT U165 ( .A1(n36), .A2(n35), .A3(n40), .Y(a1stg_expadd2_5_0[2]) );
  AOI22X1_RVT U166 ( .A1(a1stg_in2[57]), .A2(n200), .A3(a1stg_in2[54]), .A4(
        n216), .Y(n39) );
  AOI22X1_RVT U167 ( .A1(n217), .A2(a1stg_in1a[54]), .A3(n199), .A4(
        a1stg_in1a[57]), .Y(n38) );
  NAND2X0_RVT U168 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[2]), .Y(n37) );
  NAND3X0_RVT U169 ( .A1(n39), .A2(n38), .A3(n37), .Y(a2stg_exp_in[2]) );
  AOI22X1_RVT U170 ( .A1(a1stg_in2a[58]), .A2(a1stg_dp_sngopa[3]), .A3(
        a1stg_in2a[55]), .A4(a1stg_dp_dblopa[3]), .Y(\intadd_1/A[2] ) );
  NOR4X1_RVT U171 ( .A1(\intadd_1/A[2] ), .A2(\intadd_1/A[1] ), .A3(
        a1stg_expadd2_5_0[0]), .A4(\intadd_1/A[0] ), .Y(n45) );
  AOI21X1_RVT U172 ( .A1(\intadd_1/A[2] ), .A2(n40), .A3(n45), .Y(
        a1stg_expadd2_5_0[3]) );
  AOI22X1_RVT U173 ( .A1(a1stg_in2[58]), .A2(n200), .A3(a1stg_in2[55]), .A4(
        n216), .Y(n43) );
  AOI22X1_RVT U174 ( .A1(n217), .A2(a1stg_in1a[55]), .A3(n199), .A4(
        a1stg_in1a[58]), .Y(n42) );
  NAND2X0_RVT U175 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[3]), .Y(n41) );
  NAND3X0_RVT U176 ( .A1(n43), .A2(n42), .A3(n41), .Y(a2stg_exp_in[3]) );
  NAND2X0_RVT U177 ( .A1(n45), .A2(n44), .Y(n194) );
  OA21X1_RVT U178 ( .A1(n45), .A2(n44), .A3(n194), .Y(a1stg_expadd2_5_0[4]) );
  AOI22X1_RVT U179 ( .A1(a1stg_in2[59]), .A2(n200), .A3(a1stg_in2[56]), .A4(
        n216), .Y(n48) );
  AOI22X1_RVT U180 ( .A1(n217), .A2(a1stg_in1a[56]), .A3(a1stg_in1a[59]), .A4(
        n199), .Y(n47) );
  NAND2X0_RVT U181 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[4]), .Y(n46) );
  NAND3X0_RVT U182 ( .A1(n48), .A2(n47), .A3(n46), .Y(a2stg_exp_in[4]) );
  HADDX1_RVT U183 ( .A0(\intadd_1/A[4] ), .B0(n194), .SO(a1stg_expadd2_5_0[5])
         );
  AOI22X1_RVT U184 ( .A1(a1stg_in2[60]), .A2(n200), .A3(a1stg_in2[57]), .A4(
        n216), .Y(n51) );
  AOI22X1_RVT U185 ( .A1(n217), .A2(a1stg_in1a[57]), .A3(a1stg_in1a[60]), .A4(
        n199), .Y(n50) );
  NAND2X0_RVT U186 ( .A1(a1stg_fsdtoix), .A2(a1stg_expadd2_5_0[5]), .Y(n49) );
  NAND3X0_RVT U187 ( .A1(n51), .A2(n50), .A3(n49), .Y(a2stg_exp_in[5]) );
  AOI22X1_RVT U188 ( .A1(a1stg_in2a[62]), .A2(a1stg_dp_sngopa[7]), .A3(
        a1stg_dp_dblopa[7]), .A4(a1stg_in2a[59]), .Y(\intadd_1/A[6] ) );
  INVX1_RVT U189 ( .A(a4stg_in_of), .Y(n73) );
  AND2X1_RVT U190 ( .A1(a4stg_denorm_inv), .A2(add_exp_out_expadd), .Y(n297)
         );
  INVX1_RVT U191 ( .A(\intadd_3/SUM[0] ), .Y(n279) );
  NAND2X0_RVT U192 ( .A1(n297), .A2(n279), .Y(n52) );
  AND2X1_RVT U193 ( .A1(n73), .A2(n52), .Y(n54) );
  NAND2X0_RVT U194 ( .A1(a4stg_exp_11_0[1]), .A2(add_exp_out_exp1), .Y(n53) );
  AND2X1_RVT U195 ( .A1(n54), .A2(n53), .Y(n127) );
  INVX1_RVT U196 ( .A(\intadd_3/SUM[1] ), .Y(n278) );
  NAND2X0_RVT U197 ( .A1(n297), .A2(n278), .Y(n55) );
  AND2X1_RVT U198 ( .A1(n73), .A2(n55), .Y(n57) );
  NAND2X0_RVT U199 ( .A1(a4stg_exp_11_0[2]), .A2(add_exp_out_exp1), .Y(n56) );
  AND2X1_RVT U200 ( .A1(n57), .A2(n56), .Y(n129) );
  INVX1_RVT U201 ( .A(\intadd_3/SUM[2] ), .Y(n277) );
  NAND2X0_RVT U202 ( .A1(n297), .A2(n277), .Y(n58) );
  AND2X1_RVT U203 ( .A1(n73), .A2(n58), .Y(n60) );
  NAND2X0_RVT U204 ( .A1(a4stg_exp_11_0[3]), .A2(add_exp_out_exp1), .Y(n59) );
  AND2X1_RVT U205 ( .A1(n60), .A2(n59), .Y(n131) );
  INVX1_RVT U206 ( .A(\intadd_3/SUM[3] ), .Y(n276) );
  NAND2X0_RVT U207 ( .A1(n297), .A2(n276), .Y(n61) );
  AND2X1_RVT U208 ( .A1(n73), .A2(n61), .Y(n63) );
  NAND2X0_RVT U209 ( .A1(a4stg_exp_11_0[4]), .A2(add_exp_out_exp1), .Y(n62) );
  AND2X1_RVT U210 ( .A1(n63), .A2(n62), .Y(n133) );
  INVX1_RVT U211 ( .A(\intadd_3/SUM[4] ), .Y(n275) );
  NAND2X0_RVT U212 ( .A1(n297), .A2(n275), .Y(n64) );
  AND2X1_RVT U213 ( .A1(n73), .A2(n64), .Y(n66) );
  NAND2X0_RVT U214 ( .A1(a4stg_exp_11_0[5]), .A2(add_exp_out_exp1), .Y(n65) );
  AND2X1_RVT U215 ( .A1(n66), .A2(n65), .Y(n135) );
  NAND2X0_RVT U216 ( .A1(\intadd_3/n1 ), .A2(a4stg_exp2[6]), .Y(n71) );
  OAI21X1_RVT U217 ( .A1(\intadd_3/n1 ), .A2(a4stg_exp2[6]), .A3(n71), .Y(n274) );
  NAND2X0_RVT U218 ( .A1(n297), .A2(n274), .Y(n67) );
  AND2X1_RVT U219 ( .A1(n73), .A2(n67), .Y(n69) );
  NAND2X0_RVT U220 ( .A1(a4stg_exp_11_0[6]), .A2(add_exp_out_exp1), .Y(n68) );
  AND2X1_RVT U221 ( .A1(n69), .A2(n68), .Y(n137) );
  OR2X1_RVT U222 ( .A1(a4stg_exp2[7]), .A2(n71), .Y(n152) );
  AO21X1_RVT U223 ( .A1(a4stg_exp2[7]), .A2(n71), .A3(n70), .Y(n273) );
  NAND2X0_RVT U224 ( .A1(n297), .A2(n273), .Y(n72) );
  AND2X1_RVT U225 ( .A1(n73), .A2(n72), .Y(n75) );
  NAND2X0_RVT U226 ( .A1(a4stg_exp_11_0[7]), .A2(add_exp_out_exp1), .Y(n74) );
  AND2X1_RVT U227 ( .A1(n75), .A2(n74), .Y(n139) );
  NAND3X0_RVT U228 ( .A1(a3stg_exp_10_0[2]), .A2(a3stg_exp_10_0[0]), .A3(
        a3stg_exp_10_0[1]), .Y(n79) );
  NAND2X0_RVT U229 ( .A1(a6stg_step), .A2(a3stg_faddsubop), .Y(n284) );
  NOR2X0_RVT U230 ( .A1(a3stg_inc_exp_inv), .A2(n284), .Y(n240) );
  AND2X1_RVT U231 ( .A1(n79), .A2(n240), .Y(n78) );
  NAND2X0_RVT U232 ( .A1(a3stg_exp_10_0[0]), .A2(a3stg_exp_10_0[1]), .Y(n260)
         );
  NAND2X0_RVT U233 ( .A1(n76), .A2(n260), .Y(n77) );
  AND2X1_RVT U234 ( .A1(n78), .A2(n77), .Y(a4stg_exp_pre1_in[2]) );
  NAND4X0_RVT U235 ( .A1(a3stg_exp_10_0[3]), .A2(a3stg_exp_10_0[2]), .A3(
        a3stg_exp_10_0[0]), .A4(a3stg_exp_10_0[1]), .Y(n84) );
  AND2X1_RVT U236 ( .A1(n84), .A2(n240), .Y(n82) );
  NAND2X0_RVT U237 ( .A1(n80), .A2(n79), .Y(n81) );
  AND2X1_RVT U238 ( .A1(n82), .A2(n81), .Y(a4stg_exp_pre1_in[3]) );
  NAND2X0_RVT U239 ( .A1(a3stg_exp_10_0[4]), .A2(n83), .Y(n89) );
  AND2X1_RVT U240 ( .A1(n89), .A2(n240), .Y(n87) );
  NAND2X0_RVT U241 ( .A1(n85), .A2(n84), .Y(n86) );
  AND2X1_RVT U242 ( .A1(n87), .A2(n86), .Y(a4stg_exp_pre1_in[4]) );
  NAND2X0_RVT U243 ( .A1(a3stg_exp_10_0[5]), .A2(n88), .Y(n94) );
  AND2X1_RVT U244 ( .A1(n94), .A2(n240), .Y(n92) );
  NAND2X0_RVT U245 ( .A1(n90), .A2(n89), .Y(n91) );
  AND2X1_RVT U246 ( .A1(n92), .A2(n91), .Y(a4stg_exp_pre1_in[5]) );
  NAND2X0_RVT U247 ( .A1(a3stg_exp_10_0[6]), .A2(n93), .Y(n99) );
  AND2X1_RVT U248 ( .A1(n99), .A2(n240), .Y(n97) );
  NAND2X0_RVT U249 ( .A1(n95), .A2(n94), .Y(n96) );
  AND2X1_RVT U250 ( .A1(n97), .A2(n96), .Y(a4stg_exp_pre1_in[6]) );
  NAND2X0_RVT U251 ( .A1(a3stg_exp_10_0[7]), .A2(n98), .Y(n104) );
  AND2X1_RVT U252 ( .A1(n104), .A2(n240), .Y(n102) );
  NAND2X0_RVT U253 ( .A1(n100), .A2(n99), .Y(n101) );
  AND2X1_RVT U254 ( .A1(n102), .A2(n101), .Y(a4stg_exp_pre1_in[7]) );
  NAND2X0_RVT U255 ( .A1(a3stg_exp_10_0[8]), .A2(n103), .Y(n109) );
  AND2X1_RVT U256 ( .A1(n109), .A2(n240), .Y(n107) );
  NAND2X0_RVT U257 ( .A1(n105), .A2(n104), .Y(n106) );
  AND2X1_RVT U258 ( .A1(n107), .A2(n106), .Y(a4stg_exp_pre1_in[8]) );
  NAND2X0_RVT U259 ( .A1(a3stg_exp_10_0[9]), .A2(n108), .Y(n147) );
  AND2X1_RVT U260 ( .A1(n147), .A2(n240), .Y(n112) );
  NAND2X0_RVT U261 ( .A1(n110), .A2(n109), .Y(n111) );
  AND2X1_RVT U262 ( .A1(n112), .A2(n111), .Y(a4stg_exp_pre1_in[9]) );
  NAND2X0_RVT U263 ( .A1(a3stg_exp_10_0[10]), .A2(n146), .Y(n238) );
  AND2X1_RVT U264 ( .A1(n238), .A2(n240), .Y(n150) );
  NAND2X0_RVT U265 ( .A1(n148), .A2(n147), .Y(n149) );
  AND2X1_RVT U266 ( .A1(n150), .A2(n149), .Y(a4stg_exp_pre1_in[10]) );
  NAND2X0_RVT U267 ( .A1(a4stg_in_of), .A2(a4stg_dblop), .Y(n174) );
  OR2X1_RVT U268 ( .A1(a4stg_exp2[8]), .A2(n152), .Y(n168) );
  AO21X1_RVT U269 ( .A1(a4stg_exp2[8]), .A2(n152), .A3(n151), .Y(n272) );
  NAND2X0_RVT U270 ( .A1(n297), .A2(n272), .Y(n153) );
  AND2X1_RVT U271 ( .A1(n174), .A2(n153), .Y(n155) );
  NAND2X0_RVT U272 ( .A1(a4stg_exp_11_0[8]), .A2(add_exp_out_exp1), .Y(n154)
         );
  AND2X1_RVT U273 ( .A1(n155), .A2(n154), .Y(n141) );
  OR2X1_RVT U274 ( .A1(a4stg_exp2[9]), .A2(n168), .Y(n172) );
  AO21X1_RVT U275 ( .A1(a4stg_exp2[9]), .A2(n168), .A3(n156), .Y(n271) );
  NAND2X0_RVT U276 ( .A1(n297), .A2(n271), .Y(n169) );
  AND2X1_RVT U277 ( .A1(n174), .A2(n169), .Y(n171) );
  NAND2X0_RVT U278 ( .A1(a4stg_exp_11_0[9]), .A2(add_exp_out_exp1), .Y(n170)
         );
  AND2X1_RVT U279 ( .A1(n171), .A2(n170), .Y(n143) );
  NOR2X0_RVT U280 ( .A1(a4stg_exp2[10]), .A2(n172), .Y(n267) );
  AO21X1_RVT U281 ( .A1(a4stg_exp2[10]), .A2(n172), .A3(n267), .Y(n270) );
  NAND2X0_RVT U282 ( .A1(n297), .A2(n270), .Y(n173) );
  AND2X1_RVT U283 ( .A1(n174), .A2(n173), .Y(n176) );
  NAND2X0_RVT U284 ( .A1(a4stg_exp_11_0[10]), .A2(add_exp_out_exp1), .Y(n175)
         );
  AND2X1_RVT U285 ( .A1(n176), .A2(n175), .Y(n145) );
  NAND2X0_RVT U286 ( .A1(a1stg_dp_dblopa[10]), .A2(a1stg_in2a[62]), .Y(n210)
         );
  NAND2X0_RVT U287 ( .A1(a1stg_in1a[62]), .A2(a1stg_dp_dblop[10]), .Y(n177) );
  XOR2X1_RVT U288 ( .A1(n178), .A2(n177), .Y(n179) );
  XOR2X1_RVT U289 ( .A1(\intadd_1/n2 ), .A2(n179), .Y(\intadd_1/SUM[9] ) );
  OA22X1_RVT U290 ( .A1(a1stg_expadd3_in1[0]), .A2(a1stg_expadd3_in2[0]), .A3(
        a1stg_expadd3_in1[1]), .A4(a1stg_expadd3_in2[1]), .Y(n180) );
  AO21X1_RVT U291 ( .A1(a1stg_expadd3_in2[1]), .A2(a1stg_expadd3_in1[1]), .A3(
        n180), .Y(n181) );
  AO222X1_RVT U292 ( .A1(a1stg_expadd3_in2[2]), .A2(a1stg_expadd3_in1[2]), 
        .A3(a1stg_expadd3_in2[2]), .A4(n181), .A5(a1stg_expadd3_in1[2]), .A6(
        n181), .Y(n182) );
  AO222X1_RVT U293 ( .A1(a1stg_expadd3_in2[3]), .A2(a1stg_expadd3_in1[3]), 
        .A3(a1stg_expadd3_in2[3]), .A4(n182), .A5(a1stg_expadd3_in1[3]), .A6(
        n182), .Y(n183) );
  AO222X1_RVT U294 ( .A1(a1stg_expadd3_in2[4]), .A2(a1stg_expadd3_in1[4]), 
        .A3(a1stg_expadd3_in2[4]), .A4(n183), .A5(a1stg_expadd3_in1[4]), .A6(
        n183), .Y(n184) );
  AO222X1_RVT U295 ( .A1(a1stg_expadd3_in2[5]), .A2(a1stg_expadd3_in1[5]), 
        .A3(a1stg_expadd3_in2[5]), .A4(n184), .A5(a1stg_expadd3_in1[5]), .A6(
        n184), .Y(n185) );
  AO222X1_RVT U296 ( .A1(a1stg_expadd3_in2[6]), .A2(a1stg_expadd3_in1[6]), 
        .A3(a1stg_expadd3_in2[6]), .A4(n185), .A5(a1stg_expadd3_in1[6]), .A6(
        n185), .Y(n186) );
  AO222X1_RVT U297 ( .A1(a1stg_expadd3_in2[7]), .A2(a1stg_expadd3_in1[7]), 
        .A3(a1stg_expadd3_in2[7]), .A4(n186), .A5(a1stg_expadd3_in1[7]), .A6(
        n186), .Y(n187) );
  AO222X1_RVT U298 ( .A1(a1stg_expadd3_in2[8]), .A2(a1stg_expadd3_in1[8]), 
        .A3(a1stg_expadd3_in2[8]), .A4(n187), .A5(a1stg_expadd3_in1[8]), .A6(
        n187), .Y(n188) );
  AO222X1_RVT U299 ( .A1(a1stg_expadd3_in2[9]), .A2(a1stg_expadd3_in1[9]), 
        .A3(a1stg_expadd3_in2[9]), .A4(n188), .A5(a1stg_expadd3_in1[9]), .A6(
        n188), .Y(n189) );
  AOI222X1_RVT U300 ( .A1(a1stg_expadd3_in1[10]), .A2(a1stg_expadd3_in2[10]), 
        .A3(a1stg_expadd3_in1[10]), .A4(n189), .A5(a1stg_expadd3_in2[10]), 
        .A6(n189), .Y(a1stg_expadd3_11) );
  NAND2X0_RVT U301 ( .A1(a1stg_dp_dblopa[10]), .A2(a1stg_in1[62]), .Y(
        \intadd_2/A[9] ) );
  AND2X1_RVT U302 ( .A1(a1stg_in2[62]), .A2(a1stg_dp_dblop[10]), .Y(
        \intadd_2/B[9] ) );
  AOI21X1_RVT U303 ( .A1(a1stg_dp_dblopa[9]), .A2(a1stg_in1[61]), .A3(
        a1stg_op_7[9]), .Y(\intadd_2/A[8] ) );
  AND2X1_RVT U304 ( .A1(a1stg_in2[61]), .A2(a1stg_dp_dblop[9]), .Y(
        \intadd_2/B[8] ) );
  AOI21X1_RVT U305 ( .A1(a1stg_dp_dblopa[8]), .A2(a1stg_in1[60]), .A3(
        a1stg_op_7[8]), .Y(\intadd_2/A[7] ) );
  AND2X1_RVT U306 ( .A1(a1stg_in2[60]), .A2(a1stg_dp_dblop[8]), .Y(
        \intadd_2/B[7] ) );
  AO22X1_RVT U307 ( .A1(a1stg_dp_dblopa[7]), .A2(a1stg_in1[59]), .A3(
        a1stg_dp_sngopa[7]), .A4(a1stg_in1[62]), .Y(n190) );
  NOR2X0_RVT U308 ( .A1(a1stg_op_7[7]), .A2(n190), .Y(\intadd_2/A[6] ) );
  AOI22X1_RVT U309 ( .A1(a1stg_dp_dblopa[6]), .A2(a1stg_in1[58]), .A3(
        a1stg_dp_sngopa[6]), .A4(a1stg_in1[61]), .Y(\intadd_2/A[5] ) );
  AOI22X1_RVT U310 ( .A1(a1stg_dp_dblopa[5]), .A2(a1stg_in1[57]), .A3(
        a1stg_dp_sngopa[5]), .A4(a1stg_in1[60]), .Y(\intadd_2/A[4] ) );
  AOI22X1_RVT U311 ( .A1(a1stg_dp_sngopa[4]), .A2(a1stg_in1[59]), .A3(
        a1stg_dp_dblopa[4]), .A4(a1stg_in1[56]), .Y(\intadd_2/A[3] ) );
  AOI22X1_RVT U312 ( .A1(a1stg_dp_dblopa[3]), .A2(a1stg_in1[55]), .A3(
        a1stg_dp_sngopa[3]), .A4(a1stg_in1[58]), .Y(\intadd_2/A[2] ) );
  AOI22X1_RVT U313 ( .A1(a1stg_dp_sngopa[2]), .A2(a1stg_in1[57]), .A3(
        a1stg_dp_dblopa[2]), .A4(a1stg_in1[54]), .Y(\intadd_2/A[1] ) );
  AOI22X1_RVT U314 ( .A1(a1stg_dp_sngopa[1]), .A2(a1stg_in1[56]), .A3(
        a1stg_dp_dblopa[1]), .A4(a1stg_in1[53]), .Y(\intadd_2/A[0] ) );
  AO22X1_RVT U315 ( .A1(a1stg_in2[56]), .A2(a1stg_dp_sngop[1]), .A3(
        a1stg_in2[53]), .A4(a1stg_dp_dblop[1]), .Y(\intadd_2/CI ) );
  AO22X1_RVT U316 ( .A1(a1stg_in2[57]), .A2(a1stg_dp_sngop[2]), .A3(
        a1stg_in2[54]), .A4(a1stg_dp_dblop[2]), .Y(\intadd_2/B[1] ) );
  AO22X1_RVT U317 ( .A1(a1stg_in2[58]), .A2(a1stg_dp_sngop[3]), .A3(
        a1stg_in2[55]), .A4(a1stg_dp_dblop[3]), .Y(\intadd_2/B[2] ) );
  AO22X1_RVT U318 ( .A1(a1stg_in2[59]), .A2(a1stg_dp_sngop[4]), .A3(
        a1stg_in2[56]), .A4(a1stg_dp_dblop[4]), .Y(\intadd_2/B[3] ) );
  AO22X1_RVT U319 ( .A1(a1stg_in2[60]), .A2(a1stg_dp_sngop[5]), .A3(
        a1stg_in2[57]), .A4(a1stg_dp_dblop[5]), .Y(\intadd_2/B[4] ) );
  AO22X1_RVT U320 ( .A1(a1stg_in2[61]), .A2(a1stg_dp_sngop[6]), .A3(
        a1stg_in2[58]), .A4(a1stg_dp_dblop[6]), .Y(\intadd_2/B[5] ) );
  AO22X1_RVT U321 ( .A1(a1stg_in2[62]), .A2(a1stg_dp_sngop[7]), .A3(
        a1stg_in2[59]), .A4(a1stg_dp_dblop[7]), .Y(\intadd_2/B[6] ) );
  OAI21X1_RVT U322 ( .A1(n193), .A2(n192), .A3(n191), .Y(a1stg_expadd1_11_0[0]) );
  AOI22X1_RVT U324 ( .A1(a1stg_dp_dblopa[6]), .A2(a1stg_in2a[58]), .A3(
        a1stg_dp_sngopa[6]), .A4(a1stg_in2a[61]), .Y(\intadd_1/A[5] ) );
  AOI22X1_RVT U325 ( .A1(a1stg_in1a[62]), .A2(n199), .A3(n217), .A4(
        a1stg_in1a[59]), .Y(n198) );
  AOI22X1_RVT U326 ( .A1(a1stg_in2[62]), .A2(n200), .A3(a1stg_in2[59]), .A4(
        n216), .Y(n197) );
  OR2X1_RVT U327 ( .A1(\intadd_1/A[4] ), .A2(n194), .Y(n201) );
  OR2X1_RVT U328 ( .A1(\intadd_1/A[5] ), .A2(n201), .Y(n202) );
  OR2X1_RVT U329 ( .A1(\intadd_1/A[6] ), .A2(n202), .Y(n218) );
  NAND2X0_RVT U330 ( .A1(\intadd_1/A[6] ), .A2(n202), .Y(n195) );
  NAND3X0_RVT U331 ( .A1(a1stg_fsdtoix), .A2(n218), .A3(n195), .Y(n196) );
  NAND3X0_RVT U332 ( .A1(n198), .A2(n197), .A3(n196), .Y(a2stg_exp_in[7]) );
  AOI22X1_RVT U333 ( .A1(n217), .A2(a1stg_in1a[58]), .A3(a1stg_in1a[61]), .A4(
        n199), .Y(n206) );
  AOI22X1_RVT U334 ( .A1(a1stg_in2[61]), .A2(n200), .A3(a1stg_in2[58]), .A4(
        n216), .Y(n205) );
  NAND2X0_RVT U335 ( .A1(\intadd_1/A[5] ), .A2(n201), .Y(n203) );
  NAND3X0_RVT U336 ( .A1(n203), .A2(n202), .A3(a1stg_fsdtoix), .Y(n204) );
  NAND3X0_RVT U337 ( .A1(n206), .A2(n205), .A3(n204), .Y(a2stg_exp_in[6]) );
  NOR2X0_RVT U338 ( .A1(n280), .A2(a4stg_exp2[0]), .Y(\intadd_3/CI ) );
  INVX1_RVT U339 ( .A(n218), .Y(n207) );
  NAND3X0_RVT U340 ( .A1(a1stg_dp_dblopa[8]), .A2(a1stg_in2a[60]), .A3(n207), 
        .Y(n220) );
  NAND3X0_RVT U341 ( .A1(a1stg_in2a[61]), .A2(n208), .A3(a1stg_dp_dblopa[9]), 
        .Y(n214) );
  NOR3X0_RVT U342 ( .A1(n209), .A2(n210), .A3(n214), .Y(a2stg_exp_in[11]) );
  HADDX1_RVT U343 ( .A0(n210), .B0(n214), .SO(n212) );
  AO22X1_RVT U344 ( .A1(a1stg_in1a[62]), .A2(n217), .A3(a1stg_in2[62]), .A4(
        n216), .Y(n211) );
  AO21X1_RVT U345 ( .A1(a1stg_fsdtoix), .A2(n212), .A3(n211), .Y(
        a2stg_exp_in[10]) );
  NAND2X0_RVT U346 ( .A1(a1stg_in2a[61]), .A2(a1stg_dp_dblopa[9]), .Y(
        \intadd_1/A[8] ) );
  AO22X1_RVT U347 ( .A1(n217), .A2(a1stg_in1a[61]), .A3(a1stg_in2[61]), .A4(
        n216), .Y(n215) );
  NAND2X0_RVT U348 ( .A1(n220), .A2(\intadd_1/A[8] ), .Y(n213) );
  OA222X1_RVT U349 ( .A1(n215), .A2(a1stg_fsdtoix), .A3(n215), .A4(n214), .A5(
        n215), .A6(n213), .Y(a2stg_exp_in[9]) );
  NAND2X0_RVT U350 ( .A1(a1stg_dp_dblopa[8]), .A2(a1stg_in2a[60]), .Y(
        \intadd_1/A[7] ) );
  AO22X1_RVT U351 ( .A1(n217), .A2(a1stg_in1a[60]), .A3(a1stg_in2[60]), .A4(
        n216), .Y(n221) );
  NAND2X0_RVT U352 ( .A1(\intadd_1/A[7] ), .A2(n218), .Y(n219) );
  OA222X1_RVT U353 ( .A1(n221), .A2(a1stg_fsdtoix), .A3(n221), .A4(n220), .A5(
        n221), .A6(n219), .Y(a2stg_exp_in[8]) );
  AND2X1_RVT U354 ( .A1(a2stg_faddsubop), .A2(a2stg_expa[11]), .Y(N346) );
  INVX1_RVT U355 ( .A(a2stg_expadd[11]), .Y(n222) );
  AND2X1_RVT U356 ( .A1(a3stg_exp_add), .A2(n222), .Y(n235) );
  AO22X1_RVT U357 ( .A1(n235), .A2(a2stg_expadd[10]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[10]), .Y(n223) );
  OR4X1_RVT U358 ( .A1(a2stg_fxtod), .A2(a3stg_exp_7ff), .A3(a2stg_fitod), 
        .A4(n223), .Y(a3stg_exp_in[10]) );
  AO22X1_RVT U359 ( .A1(n235), .A2(a2stg_expadd[9]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[9]), .Y(n224) );
  OR2X1_RVT U360 ( .A1(a3stg_exp_7ff), .A2(n224), .Y(a3stg_exp_in[9]) );
  AO22X1_RVT U361 ( .A1(n235), .A2(a2stg_expadd[8]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[8]), .Y(n225) );
  OR2X1_RVT U362 ( .A1(a3stg_exp_7ff), .A2(n225), .Y(a3stg_exp_in[8]) );
  OR2X1_RVT U363 ( .A1(a3stg_exp_ff), .A2(a3stg_exp_7ff), .Y(n237) );
  AO22X1_RVT U364 ( .A1(n235), .A2(a2stg_expadd[7]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[7]), .Y(n226) );
  OR4X1_RVT U365 ( .A1(a2stg_fitos), .A2(a2stg_fxtos), .A3(n237), .A4(n226), 
        .Y(a3stg_exp_in[7]) );
  AO22X1_RVT U366 ( .A1(n235), .A2(a2stg_expadd[6]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[6]), .Y(n227) );
  OR2X1_RVT U367 ( .A1(n237), .A2(n227), .Y(a3stg_exp_in[6]) );
  AO22X1_RVT U368 ( .A1(n235), .A2(a2stg_expadd[5]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[5]), .Y(n228) );
  OR2X1_RVT U369 ( .A1(n229), .A2(n228), .Y(a3stg_exp_in[5]) );
  OR3X2_RVT U370 ( .A1(a2stg_fitos), .A2(a2stg_fitod), .A3(n229), .Y(n234) );
  AO22X1_RVT U371 ( .A1(n235), .A2(a2stg_expadd[4]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[4]), .Y(n230) );
  OR2X1_RVT U372 ( .A1(n234), .A2(n230), .Y(a3stg_exp_in[4]) );
  AO22X1_RVT U373 ( .A1(n235), .A2(a2stg_expadd[3]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[3]), .Y(n231) );
  OR2X1_RVT U374 ( .A1(n234), .A2(n231), .Y(a3stg_exp_in[3]) );
  AO22X1_RVT U375 ( .A1(n235), .A2(a2stg_expadd[2]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[2]), .Y(n232) );
  OR2X1_RVT U376 ( .A1(n234), .A2(n232), .Y(a3stg_exp_in[2]) );
  AO22X1_RVT U377 ( .A1(n235), .A2(a2stg_expadd[1]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[1]), .Y(n233) );
  OR2X1_RVT U378 ( .A1(n234), .A2(n233), .Y(a3stg_exp_in[1]) );
  AO22X1_RVT U379 ( .A1(n235), .A2(a2stg_expadd[0]), .A3(a2stg_faddsubop), 
        .A4(a2stg_expa[0]), .Y(n236) );
  OR2X1_RVT U380 ( .A1(n237), .A2(n236), .Y(a3stg_exp_in[0]) );
  OA221X1_RVT U381 ( .A1(\a3stg_exp[11] ), .A2(n239), .A3(n242), .A4(n238), 
        .A5(n240), .Y(a4stg_exp_pre1_in[11]) );
  OR2X1_RVT U382 ( .A1(a3stg_exp_10_0[0]), .A2(a3stg_exp_10_0[1]), .Y(n261) );
  AND3X1_RVT U383 ( .A1(n240), .A2(n260), .A3(n261), .Y(a4stg_exp_pre1_in[1])
         );
  INVX1_RVT U384 ( .A(a3stg_exp_10_0[0]), .Y(n264) );
  AND2X1_RVT U385 ( .A1(n240), .A2(n264), .Y(a4stg_exp_pre1_in[0]) );
  NOR4X1_RVT U386 ( .A1(a3stg_exp_10_0[3]), .A2(a3stg_exp_10_0[2]), .A3(
        a3stg_exp_10_0[0]), .A4(a3stg_exp_10_0[1]), .Y(n257) );
  INVX1_RVT U387 ( .A(n257), .Y(n255) );
  OR2X1_RVT U388 ( .A1(n255), .A2(a3stg_exp_10_0[4]), .Y(n254) );
  OR2X1_RVT U389 ( .A1(n254), .A2(a3stg_exp_10_0[5]), .Y(n252) );
  OR2X1_RVT U390 ( .A1(n252), .A2(a3stg_exp_10_0[6]), .Y(n250) );
  OR2X1_RVT U391 ( .A1(n250), .A2(a3stg_exp_10_0[7]), .Y(n248) );
  OR2X1_RVT U392 ( .A1(n248), .A2(a3stg_exp_10_0[8]), .Y(n246) );
  OR2X1_RVT U393 ( .A1(n246), .A2(a3stg_exp_10_0[9]), .Y(n244) );
  OR2X1_RVT U394 ( .A1(n244), .A2(a3stg_exp_10_0[10]), .Y(n241) );
  INVX1_RVT U395 ( .A(n241), .Y(n243) );
  NOR2X0_RVT U396 ( .A1(a3stg_dec_exp_inv), .A2(n284), .Y(n265) );
  OA221X1_RVT U397 ( .A1(\a3stg_exp[11] ), .A2(n243), .A3(n242), .A4(n241), 
        .A5(n265), .Y(a4stg_exp_pre3_in[11]) );
  OA221X1_RVT U398 ( .A1(n243), .A2(a3stg_exp_10_0[10]), .A3(n243), .A4(n244), 
        .A5(n265), .Y(a4stg_exp_pre3_in[10]) );
  INVX1_RVT U399 ( .A(n244), .Y(n245) );
  OA221X1_RVT U400 ( .A1(n245), .A2(a3stg_exp_10_0[9]), .A3(n245), .A4(n246), 
        .A5(n265), .Y(a4stg_exp_pre3_in[9]) );
  INVX1_RVT U401 ( .A(n246), .Y(n247) );
  OA221X1_RVT U402 ( .A1(n247), .A2(a3stg_exp_10_0[8]), .A3(n247), .A4(n248), 
        .A5(n265), .Y(a4stg_exp_pre3_in[8]) );
  INVX1_RVT U403 ( .A(n248), .Y(n249) );
  OA221X1_RVT U404 ( .A1(n249), .A2(a3stg_exp_10_0[7]), .A3(n249), .A4(n250), 
        .A5(n265), .Y(a4stg_exp_pre3_in[7]) );
  OA221X1_RVT U405 ( .A1(n251), .A2(a3stg_exp_10_0[6]), .A3(n251), .A4(n252), 
        .A5(n265), .Y(a4stg_exp_pre3_in[6]) );
  INVX1_RVT U406 ( .A(n252), .Y(n253) );
  OA221X1_RVT U407 ( .A1(n253), .A2(a3stg_exp_10_0[5]), .A3(n253), .A4(n254), 
        .A5(n265), .Y(a4stg_exp_pre3_in[5]) );
  INVX1_RVT U408 ( .A(n254), .Y(n256) );
  OA221X1_RVT U409 ( .A1(n256), .A2(a3stg_exp_10_0[4]), .A3(n256), .A4(n255), 
        .A5(n265), .Y(a4stg_exp_pre3_in[4]) );
  OR3X1_RVT U410 ( .A1(a3stg_exp_10_0[2]), .A2(a3stg_exp_10_0[0]), .A3(
        a3stg_exp_10_0[1]), .Y(n258) );
  OA221X1_RVT U411 ( .A1(n257), .A2(a3stg_exp_10_0[3]), .A3(n257), .A4(n258), 
        .A5(n265), .Y(a4stg_exp_pre3_in[3]) );
  INVX1_RVT U412 ( .A(n258), .Y(n259) );
  OA221X1_RVT U413 ( .A1(n259), .A2(a3stg_exp_10_0[2]), .A3(n259), .A4(n261), 
        .A5(n265), .Y(a4stg_exp_pre3_in[2]) );
  OA21X1_RVT U414 ( .A1(n263), .A2(n262), .A3(n265), .Y(a4stg_exp_pre3_in[1])
         );
  AND2X1_RVT U415 ( .A1(n265), .A2(n264), .Y(a4stg_exp_pre3_in[0]) );
  OR4X1_RVT U416 ( .A1(a4stg_exp_pre1[11]), .A2(a4stg_exp_pre2[11]), .A3(
        a4stg_exp_pre3[11]), .A4(a4stg_exp_pre4[11]), .Y(a4stg_exp_11_0[11])
         );
  AND3X1_RVT U417 ( .A1(n266), .A2(a4stg_denorm_inv), .A3(a6stg_step), .Y(n283) );
  HADDX1_RVT U418 ( .A0(a4stg_exp2[11]), .B0(n267), .SO(n269) );
  NOR2X0_RVT U419 ( .A1(a3stg_fdtos_inv), .A2(n282), .Y(n281) );
  AO22X1_RVT U420 ( .A1(n281), .A2(\a3stg_exp[11] ), .A3(n282), .A4(
        a4stg_exp_11_0[11]), .Y(n268) );
  AO21X1_RVT U421 ( .A1(n283), .A2(n269), .A3(n268), .Y(a4stg_exp_pre2_in[11])
         );
  AO222X1_RVT U422 ( .A1(n270), .A2(n283), .A3(a4stg_exp_11_0[10]), .A4(n282), 
        .A5(a3stg_exp_10_0[10]), .A6(n281), .Y(a4stg_exp_pre2_in[10]) );
  AO222X1_RVT U423 ( .A1(n271), .A2(n283), .A3(a4stg_exp_11_0[9]), .A4(n282), 
        .A5(a3stg_exp_10_0[9]), .A6(n281), .Y(a4stg_exp_pre2_in[9]) );
  AO222X1_RVT U424 ( .A1(n272), .A2(n283), .A3(a4stg_exp_11_0[8]), .A4(n282), 
        .A5(a3stg_exp_10_0[8]), .A6(n281), .Y(a4stg_exp_pre2_in[8]) );
  AO222X1_RVT U425 ( .A1(n273), .A2(n283), .A3(a4stg_exp_11_0[7]), .A4(n282), 
        .A5(a3stg_exp_10_0[7]), .A6(n281), .Y(a4stg_exp_pre2_in[7]) );
  AO222X1_RVT U426 ( .A1(n274), .A2(n283), .A3(a4stg_exp_11_0[6]), .A4(n282), 
        .A5(a3stg_exp_10_0[6]), .A6(n281), .Y(a4stg_exp_pre2_in[6]) );
  AO222X1_RVT U427 ( .A1(n275), .A2(n283), .A3(a4stg_exp_11_0[5]), .A4(n282), 
        .A5(a3stg_exp_10_0[5]), .A6(n281), .Y(a4stg_exp_pre2_in[5]) );
  AO222X1_RVT U428 ( .A1(n276), .A2(n283), .A3(a4stg_exp_11_0[4]), .A4(n282), 
        .A5(a3stg_exp_10_0[4]), .A6(n281), .Y(a4stg_exp_pre2_in[4]) );
  AO222X1_RVT U429 ( .A1(n277), .A2(n283), .A3(a4stg_exp_11_0[3]), .A4(n282), 
        .A5(a3stg_exp_10_0[3]), .A6(n281), .Y(a4stg_exp_pre2_in[3]) );
  AO222X1_RVT U430 ( .A1(n278), .A2(n283), .A3(a4stg_exp_11_0[2]), .A4(n282), 
        .A5(a3stg_exp_10_0[2]), .A6(n281), .Y(a4stg_exp_pre2_in[2]) );
  AO222X1_RVT U431 ( .A1(n279), .A2(n283), .A3(a4stg_exp_11_0[1]), .A4(n282), 
        .A5(a3stg_exp_10_0[1]), .A6(n281), .Y(a4stg_exp_pre2_in[1]) );
  AO21X1_RVT U432 ( .A1(a4stg_exp2[0]), .A2(n280), .A3(\intadd_3/CI ), .Y(n298) );
  AO222X1_RVT U433 ( .A1(n298), .A2(n283), .A3(a4stg_exp_11_0[0]), .A4(n282), 
        .A5(a3stg_exp_10_0[0]), .A6(n281), .Y(a4stg_exp_pre2_in[0]) );
  NOR2X0_RVT U434 ( .A1(a3stg_same_exp_inv), .A2(n284), .Y(n285) );
  AND2X1_RVT U435 ( .A1(\a3stg_exp[11] ), .A2(n285), .Y(a4stg_exp_pre4_in[11])
         );
  AND2X1_RVT U436 ( .A1(a3stg_exp_10_0[10]), .A2(n285), .Y(
        a4stg_exp_pre4_in[10]) );
  AND2X1_RVT U437 ( .A1(a3stg_exp_10_0[9]), .A2(n285), .Y(a4stg_exp_pre4_in[9]) );
  AND2X1_RVT U438 ( .A1(a3stg_exp_10_0[8]), .A2(n285), .Y(a4stg_exp_pre4_in[8]) );
  AND2X1_RVT U439 ( .A1(a3stg_exp_10_0[7]), .A2(n285), .Y(a4stg_exp_pre4_in[7]) );
  AND2X1_RVT U440 ( .A1(a3stg_exp_10_0[6]), .A2(n285), .Y(a4stg_exp_pre4_in[6]) );
  AND2X1_RVT U441 ( .A1(a3stg_exp_10_0[5]), .A2(n285), .Y(a4stg_exp_pre4_in[5]) );
  AND2X1_RVT U442 ( .A1(a3stg_exp_10_0[4]), .A2(n285), .Y(a4stg_exp_pre4_in[4]) );
  AND2X1_RVT U443 ( .A1(a3stg_exp_10_0[3]), .A2(n285), .Y(a4stg_exp_pre4_in[3]) );
  AND2X1_RVT U444 ( .A1(a3stg_exp_10_0[2]), .A2(n285), .Y(a4stg_exp_pre4_in[2]) );
  AND2X1_RVT U445 ( .A1(a3stg_exp_10_0[1]), .A2(n285), .Y(a4stg_exp_pre4_in[1]) );
  AND2X1_RVT U446 ( .A1(a3stg_exp_10_0[0]), .A2(n285), .Y(a4stg_exp_pre4_in[0]) );
  NAND2X0_RVT U447 ( .A1(inq_op[1]), .A2(inq_in2[52]), .Y(n167) );
  NAND2X0_RVT U448 ( .A1(inq_op[1]), .A2(inq_in2[53]), .Y(n166) );
  NAND2X0_RVT U449 ( .A1(inq_op[1]), .A2(inq_in2[54]), .Y(n165) );
  OR2X1_RVT U450 ( .A1(add_exp_out3[10]), .A2(add_exp_out4[10]), .Y(n286) );
  NAND3X0_RVT U451 ( .A1(n286), .A2(add_exp_out1[10]), .A3(add_exp_out2[10]), 
        .Y(add_exp_out[10]) );
  OR2X1_RVT U452 ( .A1(add_exp_out3[9]), .A2(add_exp_out4[9]), .Y(n287) );
  NAND3X0_RVT U453 ( .A1(n287), .A2(add_exp_out1[9]), .A3(add_exp_out2[9]), 
        .Y(add_exp_out[9]) );
  OR2X1_RVT U454 ( .A1(add_exp_out3[8]), .A2(add_exp_out4[8]), .Y(n288) );
  NAND3X0_RVT U455 ( .A1(n288), .A2(add_exp_out1[8]), .A3(add_exp_out2[8]), 
        .Y(add_exp_out[8]) );
  OR2X1_RVT U456 ( .A1(add_exp_out3[7]), .A2(add_exp_out4[7]), .Y(n289) );
  NAND3X0_RVT U457 ( .A1(n289), .A2(add_exp_out1[7]), .A3(add_exp_out2[7]), 
        .Y(add_exp_out[7]) );
  OR2X1_RVT U458 ( .A1(add_exp_out3[6]), .A2(add_exp_out4[6]), .Y(n290) );
  NAND3X0_RVT U459 ( .A1(n290), .A2(add_exp_out1[6]), .A3(add_exp_out2[6]), 
        .Y(add_exp_out[6]) );
  OR2X1_RVT U460 ( .A1(add_exp_out3[5]), .A2(add_exp_out4[5]), .Y(n291) );
  NAND3X0_RVT U461 ( .A1(n291), .A2(add_exp_out1[5]), .A3(add_exp_out2[5]), 
        .Y(add_exp_out[5]) );
  OR2X1_RVT U462 ( .A1(add_exp_out3[4]), .A2(add_exp_out4[4]), .Y(n292) );
  NAND3X0_RVT U463 ( .A1(n292), .A2(add_exp_out1[4]), .A3(add_exp_out2[4]), 
        .Y(add_exp_out[4]) );
  OR2X1_RVT U464 ( .A1(add_exp_out3[3]), .A2(add_exp_out4[3]), .Y(n293) );
  NAND3X0_RVT U465 ( .A1(n293), .A2(add_exp_out1[3]), .A3(add_exp_out2[3]), 
        .Y(add_exp_out[3]) );
  OR2X1_RVT U466 ( .A1(add_exp_out3[2]), .A2(add_exp_out4[2]), .Y(n294) );
  NAND3X0_RVT U467 ( .A1(n294), .A2(add_exp_out1[2]), .A3(add_exp_out2[2]), 
        .Y(add_exp_out[2]) );
  OR2X1_RVT U468 ( .A1(add_exp_out3[1]), .A2(add_exp_out4[1]), .Y(n295) );
  NAND3X0_RVT U469 ( .A1(n295), .A2(add_exp_out1[1]), .A3(add_exp_out2[1]), 
        .Y(add_exp_out[1]) );
  OR2X1_RVT U470 ( .A1(add_exp_out3[0]), .A2(add_exp_out4[0]), .Y(n296) );
  NAND3X0_RVT U471 ( .A1(n296), .A2(add_exp_out1[0]), .A3(add_exp_out2[0]), 
        .Y(add_exp_out[0]) );
  NAND2X0_RVT U472 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[10]), .Y(n144)
         );
  NAND2X0_RVT U473 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[9]), .Y(n142) );
  NAND2X0_RVT U474 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[8]), .Y(n140) );
  NAND2X0_RVT U475 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[7]), .Y(n138) );
  NAND2X0_RVT U476 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[6]), .Y(n136) );
  NAND2X0_RVT U477 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[5]), .Y(n134) );
  NAND2X0_RVT U478 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[4]), .Y(n132) );
  NAND2X0_RVT U479 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[3]), .Y(n130) );
  NAND2X0_RVT U480 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[2]), .Y(n128) );
  NAND2X0_RVT U481 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[1]), .Y(n126) );
  AOI222X1_RVT U482 ( .A1(n298), .A2(n297), .A3(a4stg_in_of), .A4(
        a4stg_to_0_inv), .A5(a4stg_exp_11_0[0]), .A6(add_exp_out_exp1), .Y(
        n125) );
  NAND2X0_RVT U483 ( .A1(add_exp_out_exp), .A2(a4stg_exp_11_0[0]), .Y(n124) );
  NAND2X0_RVT U484 ( .A1(n303), .A2(n300), .Y(n123) );
  AO221X1_RVT U485 ( .A1(n300), .A2(n299), .A3(a4stg_exp_11_0[0]), .A4(
        a4stg_exp_11_0[1]), .A5(n306), .Y(n122) );
  NAND2X0_RVT U486 ( .A1(a4stg_exp_11_0[0]), .A2(a4stg_exp_11_0[1]), .Y(n301)
         );
  NAND2X0_RVT U487 ( .A1(n302), .A2(n301), .Y(n305) );
  NAND3X0_RVT U488 ( .A1(n305), .A2(n304), .A3(n303), .Y(n121) );
  AO221X1_RVT U489 ( .A1(n309), .A2(n308), .A3(a4stg_exp_11_0[10]), .A4(n307), 
        .A5(n306), .Y(n113) );
  OA21X1_RVT U490 ( .A1(a1stg_expadd2_5_0[0]), .A2(n311), .A3(n310), .Y(
        a1stg_expadd4_inv[0]) );
  AO22X1_RVT U491 ( .A1(a1stg_in1a[56]), .A2(a1stg_dp_sngop[1]), .A3(
        a1stg_in1a[53]), .A4(a1stg_dp_dblop[1]), .Y(\intadd_1/CI ) );
  AO22X1_RVT U492 ( .A1(a1stg_in1a[57]), .A2(a1stg_dp_sngop[2]), .A3(
        a1stg_in1a[54]), .A4(a1stg_dp_dblop[2]), .Y(\intadd_1/B[1] ) );
  AO22X1_RVT U493 ( .A1(a1stg_in1a[58]), .A2(a1stg_dp_sngop[3]), .A3(
        a1stg_in1a[55]), .A4(a1stg_dp_dblop[3]), .Y(\intadd_1/B[2] ) );
  AO22X1_RVT U494 ( .A1(a1stg_in1a[59]), .A2(a1stg_dp_sngop[4]), .A3(
        a1stg_in1a[56]), .A4(a1stg_dp_dblop[4]), .Y(\intadd_1/B[3] ) );
  AO22X1_RVT U495 ( .A1(a1stg_in1a[60]), .A2(a1stg_dp_sngop[5]), .A3(
        a1stg_in1a[57]), .A4(a1stg_dp_dblop[5]), .Y(\intadd_1/B[4] ) );
  AO22X1_RVT U496 ( .A1(a1stg_in1a[61]), .A2(a1stg_dp_sngop[6]), .A3(
        a1stg_in1a[58]), .A4(a1stg_dp_dblop[6]), .Y(\intadd_1/B[5] ) );
  AO22X1_RVT U497 ( .A1(a1stg_in1a[62]), .A2(a1stg_dp_sngop[7]), .A3(
        a1stg_in1a[59]), .A4(a1stg_dp_dblop[7]), .Y(\intadd_1/B[6] ) );
  AND2X1_RVT U498 ( .A1(a1stg_in1a[60]), .A2(a1stg_dp_dblop[8]), .Y(
        \intadd_1/B[7] ) );
  AND2X1_RVT U499 ( .A1(a1stg_in1a[61]), .A2(a1stg_dp_dblop[9]), .Y(
        \intadd_1/B[8] ) );
endmodule


module fpu_in2_gt_in1_3b_0 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_2b_0 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [1:0] din1;
  input [1:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6;

  INVX0_RVT U1 ( .A(n4), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[0]), .Y(n2) );
  NAND2X0_RVT U3 ( .A1(din2[0]), .A2(n2), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[1]), .Y(n3) );
  AO222X1_RVT U5 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n3), .A5(n1), .A6(
        n3), .Y(din2_gt_din1) );
  OA22X1_RVT U6 ( .A1(din2[1]), .A2(n3), .A3(din2[0]), .A4(n2), .Y(n6) );
  NAND2X0_RVT U7 ( .A1(din2[1]), .A2(n3), .Y(n5) );
  NAND3X0_RVT U8 ( .A1(n6), .A2(n5), .A3(n4), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3to1_0 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U2 ( .A(din2_neq_din1_mid), .Y(n1) );
  INVX0_RVT U3 ( .A(din2_neq_din1_hi), .Y(n3) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_1 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX1_RVT U2 ( .A(din2_neq_din1_hi), .Y(n3) );
  INVX1_RVT U3 ( .A(din2_neq_din1_mid), .Y(n1) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_2 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U2 ( .A(din2_neq_din1_hi), .Y(n3) );
  INVX0_RVT U3 ( .A(din2_neq_din1_mid), .Y(n1) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_3 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_neq_din1_mid), .Y(n1) );
  OR3X1_RVT U2 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U3 ( .A(din2_neq_din1_hi), .Y(n3) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_4 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_neq_din1_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_neq_din1_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_5 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U2 ( .A(din2_neq_din1_mid), .Y(n1) );
  INVX0_RVT U3 ( .A(din2_neq_din1_hi), .Y(n3) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_6 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U2 ( .A(din2_neq_din1_hi), .Y(n3) );
  INVX0_RVT U3 ( .A(din2_neq_din1_mid), .Y(n1) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3to1_7 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_neq_din1_hi), .A2(din2_neq_din1_mid), .A3(
        din2_neq_din1_lo), .Y(din2_neq_din1) );
  INVX0_RVT U2 ( .A(din2_neq_din1_hi), .Y(n3) );
  INVX0_RVT U3 ( .A(din2_neq_din1_mid), .Y(n1) );
  AO22X1_RVT U4 ( .A1(din2_neq_din1_mid), .A2(din2_gt_din1_mid), .A3(n1), .A4(
        din2_gt_din1_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_hi), .A2(din2_gt_din1_hi), .A3(n3), .A4(n2), .Y(din2_gt_din1) );
endmodule


module fpu_in2_gt_in1_3b_1 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U3 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U4 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U5 ( .A(n8), .Y(n1) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_2 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_3 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_4 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_5 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_6 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_7 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_8 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_9 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_10 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U3 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U4 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U5 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U6 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U7 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  INVX1_RVT U8 ( .A(din2[2]), .Y(n5) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_11 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U3 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U4 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U5 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U6 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U7 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  INVX1_RVT U8 ( .A(din2[2]), .Y(n5) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_12 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_13 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U3 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U4 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U5 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U6 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U7 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  INVX1_RVT U8 ( .A(din2[2]), .Y(n5) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_14 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U3 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U4 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U5 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U6 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U7 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  INVX1_RVT U8 ( .A(din2[2]), .Y(n5) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_15 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_3b_16 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX0_RVT U1 ( .A(n8), .Y(n1) );
  INVX0_RVT U2 ( .A(din2[2]), .Y(n5) );
  INVX1_RVT U3 ( .A(din1[2]), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[0]), .Y(n3) );
  NAND2X0_RVT U5 ( .A1(din2[0]), .A2(n3), .Y(n8) );
  INVX1_RVT U6 ( .A(din1[1]), .Y(n6) );
  AO222X1_RVT U7 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n6), .A5(n1), .A6(
        n6), .Y(n2) );
  AO222X1_RVT U8 ( .A1(din2[2]), .A2(n4), .A3(din2[2]), .A4(n2), .A5(n4), .A6(
        n2), .Y(din2_gt_din1) );
  OA222X1_RVT U9 ( .A1(din1[2]), .A2(n5), .A3(n4), .A4(din2[2]), .A5(din2[0]), 
        .A6(n3), .Y(n10) );
  NAND2X0_RVT U10 ( .A1(din2[1]), .A2(n6), .Y(n9) );
  OR2X1_RVT U11 ( .A1(n6), .A2(din2[1]), .Y(n7) );
  NAND4X0_RVT U12 ( .A1(n10), .A2(n9), .A3(n8), .A4(n7), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_2b_1 ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [1:0] din1;
  input [1:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   n1, n2, n3, n4, n5, n6;

  INVX0_RVT U1 ( .A(n4), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[0]), .Y(n2) );
  NAND2X0_RVT U3 ( .A1(din2[0]), .A2(n2), .Y(n4) );
  INVX1_RVT U4 ( .A(din1[1]), .Y(n3) );
  AO222X1_RVT U5 ( .A1(din2[1]), .A2(n1), .A3(din2[1]), .A4(n3), .A5(n1), .A6(
        n3), .Y(din2_gt_din1) );
  OA22X1_RVT U6 ( .A1(din2[1]), .A2(n3), .A3(din2[0]), .A4(n2), .Y(n6) );
  NAND2X0_RVT U7 ( .A1(din2[1]), .A2(n3), .Y(n5) );
  NAND3X0_RVT U8 ( .A1(n6), .A2(n5), .A3(n4), .Y(din2_neq_din1) );
endmodule


module fpu_in2_gt_in1_frac ( din1, din2, sngop, expadd11, expeq, din2_neq_din1, 
        din2_gt_din1, din2_gt1_din1 );
  input [54:0] din1;
  input [54:0] din2;
  input sngop, expadd11, expeq;
  output din2_neq_din1, din2_gt_din1, din2_gt1_din1;
  wire   din2_neq_din1_54_52, din2_gt_din1_54_52, din2_neq_din1_51_50,
         din2_gt_din1_51_50, din2_neq_din1_49_48, din2_gt_din1_49_48,
         din2_neq_din1_47_45, din2_gt_din1_47_45, din2_neq_din1_44_42,
         din2_gt_din1_44_42, din2_neq_din1_41_39, din2_gt_din1_41_39,
         din2_neq_din1_38_36, din2_gt_din1_38_36, din2_neq_din1_35_33,
         din2_gt_din1_35_33, din2_neq_din1_32_30, din2_gt_din1_32_30,
         din2_neq_din1_29_27, din2_gt_din1_29_27, din2_neq_din1_26_24,
         din2_gt_din1_26_24, din2_neq_din1_23_21, din2_gt_din1_23_21,
         din2_neq_din1_20_18, din2_gt_din1_20_18, din2_neq_din1_17_15,
         din2_gt_din1_17_15, din2_neq_din1_14_12, din2_gt_din1_14_12,
         din2_neq_din1_11_9, din2_gt_din1_11_9, din2_neq_din1_8_6,
         din2_gt_din1_8_6, din2_neq_din1_5_3, din2_gt_din1_5_3,
         din2_neq_din1_2_0, din2_gt_din1_2_0, din2_neq_din1_51_45,
         din2_gt_din1_51_45, din2_neq_din1_44_36, din2_gt_din1_44_36,
         din2_neq_din1_35_27, din2_gt_din1_35_27, din2_neq_din1_26_18,
         din2_gt_din1_26_18, din2_neq_din1_17_9, din2_gt_din1_17_9,
         din2_neq_din1_8_0, din2_gt_din1_8_0, din2_neq_din1_51_27,
         din2_gt_din1_51_27, din2_neq_din1_26_0, din2_gt_din1_26_0, n1, n2, n3,
         n4;

  fpu_in2_gt_in1_3b_0 fpu_in2_gt_in1_54_52 ( .din1(din1[54:52]), .din2(
        din2[54:52]), .din2_neq_din1(din2_neq_din1_54_52), .din2_gt_din1(
        din2_gt_din1_54_52) );
  fpu_in2_gt_in1_2b_0 fpu_in2_gt_in1_51_50 ( .din1(din1[51:50]), .din2(
        din2[51:50]), .din2_neq_din1(din2_neq_din1_51_50), .din2_gt_din1(
        din2_gt_din1_51_50) );
  fpu_in2_gt_in1_2b_1 fpu_in2_gt_in1_49_48 ( .din1(din1[49:48]), .din2(
        din2[49:48]), .din2_neq_din1(din2_neq_din1_49_48), .din2_gt_din1(
        din2_gt_din1_49_48) );
  fpu_in2_gt_in1_3b_16 fpu_in2_gt_in1_47_45 ( .din1(din1[47:45]), .din2(
        din2[47:45]), .din2_neq_din1(din2_neq_din1_47_45), .din2_gt_din1(
        din2_gt_din1_47_45) );
  fpu_in2_gt_in1_3b_15 fpu_in2_gt_in1_44_42 ( .din1(din1[44:42]), .din2(
        din2[44:42]), .din2_neq_din1(din2_neq_din1_44_42), .din2_gt_din1(
        din2_gt_din1_44_42) );
  fpu_in2_gt_in1_3b_14 fpu_in2_gt_in1_41_39 ( .din1(din1[41:39]), .din2(
        din2[41:39]), .din2_neq_din1(din2_neq_din1_41_39), .din2_gt_din1(
        din2_gt_din1_41_39) );
  fpu_in2_gt_in1_3b_13 fpu_in2_gt_in1_38_36 ( .din1(din1[38:36]), .din2(
        din2[38:36]), .din2_neq_din1(din2_neq_din1_38_36), .din2_gt_din1(
        din2_gt_din1_38_36) );
  fpu_in2_gt_in1_3b_12 fpu_in2_gt_in1_35_33 ( .din1(din1[35:33]), .din2(
        din2[35:33]), .din2_neq_din1(din2_neq_din1_35_33), .din2_gt_din1(
        din2_gt_din1_35_33) );
  fpu_in2_gt_in1_3b_11 fpu_in2_gt_in1_32_30 ( .din1(din1[32:30]), .din2(
        din2[32:30]), .din2_neq_din1(din2_neq_din1_32_30), .din2_gt_din1(
        din2_gt_din1_32_30) );
  fpu_in2_gt_in1_3b_10 fpu_in2_gt_in1_29_27 ( .din1(din1[29:27]), .din2(
        din2[29:27]), .din2_neq_din1(din2_neq_din1_29_27), .din2_gt_din1(
        din2_gt_din1_29_27) );
  fpu_in2_gt_in1_3b_9 fpu_in2_gt_in1_26_24 ( .din1(din1[26:24]), .din2(
        din2[26:24]), .din2_neq_din1(din2_neq_din1_26_24), .din2_gt_din1(
        din2_gt_din1_26_24) );
  fpu_in2_gt_in1_3b_8 fpu_in2_gt_in1_23_21 ( .din1(din1[23:21]), .din2(
        din2[23:21]), .din2_neq_din1(din2_neq_din1_23_21), .din2_gt_din1(
        din2_gt_din1_23_21) );
  fpu_in2_gt_in1_3b_7 fpu_in2_gt_in1_20_18 ( .din1(din1[20:18]), .din2(
        din2[20:18]), .din2_neq_din1(din2_neq_din1_20_18), .din2_gt_din1(
        din2_gt_din1_20_18) );
  fpu_in2_gt_in1_3b_6 fpu_in2_gt_in1_17_15 ( .din1(din1[17:15]), .din2(
        din2[17:15]), .din2_neq_din1(din2_neq_din1_17_15), .din2_gt_din1(
        din2_gt_din1_17_15) );
  fpu_in2_gt_in1_3b_5 fpu_in2_gt_in1_14_12 ( .din1(din1[14:12]), .din2(
        din2[14:12]), .din2_neq_din1(din2_neq_din1_14_12), .din2_gt_din1(
        din2_gt_din1_14_12) );
  fpu_in2_gt_in1_3b_4 fpu_in2_gt_in1_11_9 ( .din1(din1[11:9]), .din2(
        din2[11:9]), .din2_neq_din1(din2_neq_din1_11_9), .din2_gt_din1(
        din2_gt_din1_11_9) );
  fpu_in2_gt_in1_3b_3 fpu_in2_gt_in1_8_6 ( .din1(din1[8:6]), .din2(din2[8:6]), 
        .din2_neq_din1(din2_neq_din1_8_6), .din2_gt_din1(din2_gt_din1_8_6) );
  fpu_in2_gt_in1_3b_2 fpu_in2_gt_in1_5_3 ( .din1(din1[5:3]), .din2(din2[5:3]), 
        .din2_neq_din1(din2_neq_din1_5_3), .din2_gt_din1(din2_gt_din1_5_3) );
  fpu_in2_gt_in1_3b_1 fpu_in2_gt_in1_2_0 ( .din1(din1[2:0]), .din2(din2[2:0]), 
        .din2_neq_din1(din2_neq_din1_2_0), .din2_gt_din1(din2_gt_din1_2_0) );
  fpu_in2_gt_in1_3to1_0 fpu_in2_gt_in1_51_45 ( .din2_neq_din1_hi(
        din2_neq_din1_51_50), .din2_gt_din1_hi(din2_gt_din1_51_50), 
        .din2_neq_din1_mid(din2_neq_din1_49_48), .din2_gt_din1_mid(
        din2_gt_din1_49_48), .din2_neq_din1_lo(din2_neq_din1_47_45), 
        .din2_gt_din1_lo(din2_gt_din1_47_45), .din2_neq_din1(
        din2_neq_din1_51_45), .din2_gt_din1(din2_gt_din1_51_45) );
  fpu_in2_gt_in1_3to1_7 fpu_in2_gt_in1_44_36 ( .din2_neq_din1_hi(
        din2_neq_din1_44_42), .din2_gt_din1_hi(din2_gt_din1_44_42), 
        .din2_neq_din1_mid(din2_neq_din1_41_39), .din2_gt_din1_mid(
        din2_gt_din1_41_39), .din2_neq_din1_lo(din2_neq_din1_38_36), 
        .din2_gt_din1_lo(din2_gt_din1_38_36), .din2_neq_din1(
        din2_neq_din1_44_36), .din2_gt_din1(din2_gt_din1_44_36) );
  fpu_in2_gt_in1_3to1_6 fpu_in2_gt_in1_35_27 ( .din2_neq_din1_hi(
        din2_neq_din1_35_33), .din2_gt_din1_hi(din2_gt_din1_35_33), 
        .din2_neq_din1_mid(din2_neq_din1_32_30), .din2_gt_din1_mid(
        din2_gt_din1_32_30), .din2_neq_din1_lo(din2_neq_din1_29_27), 
        .din2_gt_din1_lo(din2_gt_din1_29_27), .din2_neq_din1(
        din2_neq_din1_35_27), .din2_gt_din1(din2_gt_din1_35_27) );
  fpu_in2_gt_in1_3to1_5 fpu_in2_gt_in1_26_18 ( .din2_neq_din1_hi(
        din2_neq_din1_26_24), .din2_gt_din1_hi(din2_gt_din1_26_24), 
        .din2_neq_din1_mid(din2_neq_din1_23_21), .din2_gt_din1_mid(
        din2_gt_din1_23_21), .din2_neq_din1_lo(din2_neq_din1_20_18), 
        .din2_gt_din1_lo(din2_gt_din1_20_18), .din2_neq_din1(
        din2_neq_din1_26_18), .din2_gt_din1(din2_gt_din1_26_18) );
  fpu_in2_gt_in1_3to1_4 fpu_in2_gt_in1_17_9 ( .din2_neq_din1_hi(
        din2_neq_din1_17_15), .din2_gt_din1_hi(din2_gt_din1_17_15), 
        .din2_neq_din1_mid(din2_neq_din1_14_12), .din2_gt_din1_mid(
        din2_gt_din1_14_12), .din2_neq_din1_lo(din2_neq_din1_11_9), 
        .din2_gt_din1_lo(din2_gt_din1_11_9), .din2_neq_din1(din2_neq_din1_17_9), .din2_gt_din1(din2_gt_din1_17_9) );
  fpu_in2_gt_in1_3to1_3 fpu_in2_gt_in1_8_0 ( .din2_neq_din1_hi(
        din2_neq_din1_8_6), .din2_gt_din1_hi(din2_gt_din1_8_6), 
        .din2_neq_din1_mid(din2_neq_din1_5_3), .din2_gt_din1_mid(
        din2_gt_din1_5_3), .din2_neq_din1_lo(din2_neq_din1_2_0), 
        .din2_gt_din1_lo(din2_gt_din1_2_0), .din2_neq_din1(din2_neq_din1_8_0), 
        .din2_gt_din1(din2_gt_din1_8_0) );
  fpu_in2_gt_in1_3to1_2 fpu_in2_gt_in1_51_27 ( .din2_neq_din1_hi(
        din2_neq_din1_51_45), .din2_gt_din1_hi(din2_gt_din1_51_45), 
        .din2_neq_din1_mid(din2_neq_din1_44_36), .din2_gt_din1_mid(
        din2_gt_din1_44_36), .din2_neq_din1_lo(din2_neq_din1_35_27), 
        .din2_gt_din1_lo(din2_gt_din1_35_27), .din2_neq_din1(
        din2_neq_din1_51_27), .din2_gt_din1(din2_gt_din1_51_27) );
  fpu_in2_gt_in1_3to1_1 fpu_in2_gt_in1_26_0 ( .din2_neq_din1_hi(
        din2_neq_din1_26_18), .din2_gt_din1_hi(din2_gt_din1_26_18), 
        .din2_neq_din1_mid(din2_neq_din1_17_9), .din2_gt_din1_mid(
        din2_gt_din1_17_9), .din2_neq_din1_lo(din2_neq_din1_8_0), 
        .din2_gt_din1_lo(din2_gt_din1_8_0), .din2_neq_din1(din2_neq_din1_26_0), 
        .din2_gt_din1(din2_gt_din1_26_0) );
  INVX0_RVT U1 ( .A(din2_neq_din1_51_27), .Y(n1) );
  INVX0_RVT U2 ( .A(n3), .Y(n4) );
  NAND2X0_RVT U3 ( .A1(sngop), .A2(din2_neq_din1_54_52), .Y(n3) );
  OR3X2_RVT U4 ( .A1(din2_neq_din1_51_27), .A2(n4), .A3(din2_neq_din1_26_0), 
        .Y(din2_neq_din1) );
  AO22X1_RVT U5 ( .A1(din2_neq_din1_51_27), .A2(din2_gt_din1_51_27), .A3(n1), 
        .A4(din2_gt_din1_26_0), .Y(n2) );
  AO22X1_RVT U6 ( .A1(n4), .A2(din2_gt_din1_54_52), .A3(n3), .A4(n2), .Y(
        din2_gt_din1) );
  AO21X1_RVT U7 ( .A1(din2_gt_din1), .A2(expeq), .A3(expadd11), .Y(
        din2_gt1_din1) );
endmodule


module fpu_denorm_3b_0 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3to1_0 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_1 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  INVX0_RVT U3 ( .A(din2_din1_nz_hi), .Y(n3) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_2 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  INVX0_RVT U3 ( .A(din2_din1_nz_hi), .Y(n3) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_3 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  OR3X1_RVT U1 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  INVX0_RVT U2 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U3 ( .A(din2_din1_nz_mid), .Y(n1) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_4 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_5 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_6 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3to1_7 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3;

  INVX0_RVT U1 ( .A(din2_din1_nz_hi), .Y(n3) );
  INVX0_RVT U2 ( .A(din2_din1_nz_mid), .Y(n1) );
  OR3X1_RVT U3 ( .A1(din2_din1_nz_hi), .A2(din2_din1_nz_mid), .A3(
        din2_din1_nz_lo), .Y(din2_din1_nz) );
  AO22X1_RVT U4 ( .A1(din2_din1_nz_mid), .A2(din2_din1_denorm_mid), .A3(n1), 
        .A4(din2_din1_denorm_lo), .Y(n2) );
  AO22X1_RVT U5 ( .A1(din2_din1_nz_hi), .A2(din2_din1_denorm_hi), .A3(n3), 
        .A4(n2), .Y(din2_din1_denorm) );
endmodule


module fpu_denorm_3b_1 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_2 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_3 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_4 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_5 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_6 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_7 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_8 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_9 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_10 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_11 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_12 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_13 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_14 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_15 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_16 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_3b_17 ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   n1, n2, n3, n4, n5;

  INVX0_RVT U1 ( .A(din1[1]), .Y(n1) );
  INVX1_RVT U2 ( .A(din1[2]), .Y(n3) );
  OA221X1_RVT U3 ( .A1(din2[1]), .A2(din2[0]), .A3(din2[1]), .A4(n1), .A5(n3), 
        .Y(n2) );
  OR2X1_RVT U4 ( .A1(din2[2]), .A2(n2), .Y(din2_din1_denorm) );
  NOR4X1_RVT U5 ( .A1(din2[1]), .A2(din1[1]), .A3(din2[0]), .A4(din1[0]), .Y(
        n5) );
  INVX1_RVT U6 ( .A(din2[2]), .Y(n4) );
  NAND3X0_RVT U7 ( .A1(n5), .A2(n4), .A3(n3), .Y(din2_din1_nz) );
endmodule


module fpu_denorm_frac ( din1, din2, din2_din1_denorm, din2_din1_denorm_inv, 
        din2_din1_denorma, din2_din1_denorm_inva );
  input [53:0] din1;
  input [53:0] din2;
  output din2_din1_denorm, din2_din1_denorm_inv, din2_din1_denorma,
         din2_din1_denorm_inva;
  wire   din2_din1_nz_53_51, din2_din1_denorm_53_51, din2_din1_nz_50_48,
         din2_din1_denorm_50_48, din2_din1_nz_47_45, din2_din1_denorm_47_45,
         din2_din1_nz_44_42, din2_din1_denorm_44_42, din2_din1_nz_41_39,
         din2_din1_denorm_41_39, din2_din1_nz_38_36, din2_din1_denorm_38_36,
         din2_din1_nz_35_33, din2_din1_denorm_35_33, din2_din1_nz_32_30,
         din2_din1_denorm_32_30, din2_din1_nz_29_27, din2_din1_denorm_29_27,
         din2_din1_nz_26_24, din2_din1_denorm_26_24, din2_din1_nz_23_21,
         din2_din1_denorm_23_21, din2_din1_nz_20_18, din2_din1_denorm_20_18,
         din2_din1_nz_17_15, din2_din1_denorm_17_15, din2_din1_nz_14_12,
         din2_din1_denorm_14_12, din2_din1_nz_11_9, din2_din1_denorm_11_9,
         din2_din1_nz_8_6, din2_din1_denorm_8_6, din2_din1_nz_5_3,
         din2_din1_denorm_5_3, din2_din1_nz_2_0, din2_din1_denorm_2_0,
         din2_din1_nz_53_45, din2_din1_denorm_53_45, din2_din1_nz_44_36,
         din2_din1_denorm_44_36, din2_din1_nz_35_27, din2_din1_denorm_35_27,
         din2_din1_nz_26_18, din2_din1_denorm_26_18, din2_din1_nz_17_9,
         din2_din1_denorm_17_9, din2_din1_nz_8_0, din2_din1_denorm_8_0,
         din2_din1_nz_53_27, din2_din1_denorm_53_27, din2_din1_nz_26_0,
         din2_din1_denorm_26_0, n1, n2, din2_din1_denorm;
  assign din2_din1_denorma = din2_din1_denorm;

  fpu_denorm_3b_0 i_fpu_denorm_53_51 ( .din1(din1[53:51]), .din2(din2[53:51]), 
        .din2_din1_nz(din2_din1_nz_53_51), .din2_din1_denorm(
        din2_din1_denorm_53_51) );
  fpu_denorm_3b_17 i_fpu_denorm_50_48 ( .din1(din1[50:48]), .din2(din2[50:48]), 
        .din2_din1_nz(din2_din1_nz_50_48), .din2_din1_denorm(
        din2_din1_denorm_50_48) );
  fpu_denorm_3b_16 i_fpu_denorm_47_45 ( .din1(din1[47:45]), .din2(din2[47:45]), 
        .din2_din1_nz(din2_din1_nz_47_45), .din2_din1_denorm(
        din2_din1_denorm_47_45) );
  fpu_denorm_3b_15 i_fpu_denorm_44_42 ( .din1(din1[44:42]), .din2(din2[44:42]), 
        .din2_din1_nz(din2_din1_nz_44_42), .din2_din1_denorm(
        din2_din1_denorm_44_42) );
  fpu_denorm_3b_14 i_fpu_denorm_41_39 ( .din1(din1[41:39]), .din2(din2[41:39]), 
        .din2_din1_nz(din2_din1_nz_41_39), .din2_din1_denorm(
        din2_din1_denorm_41_39) );
  fpu_denorm_3b_13 i_fpu_denorm_38_36 ( .din1(din1[38:36]), .din2(din2[38:36]), 
        .din2_din1_nz(din2_din1_nz_38_36), .din2_din1_denorm(
        din2_din1_denorm_38_36) );
  fpu_denorm_3b_12 i_fpu_denorm_35_33 ( .din1(din1[35:33]), .din2(din2[35:33]), 
        .din2_din1_nz(din2_din1_nz_35_33), .din2_din1_denorm(
        din2_din1_denorm_35_33) );
  fpu_denorm_3b_11 i_fpu_denorm_32_30 ( .din1(din1[32:30]), .din2(din2[32:30]), 
        .din2_din1_nz(din2_din1_nz_32_30), .din2_din1_denorm(
        din2_din1_denorm_32_30) );
  fpu_denorm_3b_10 i_fpu_denorm_29_27 ( .din1(din1[29:27]), .din2(din2[29:27]), 
        .din2_din1_nz(din2_din1_nz_29_27), .din2_din1_denorm(
        din2_din1_denorm_29_27) );
  fpu_denorm_3b_9 i_fpu_denorm_26_24 ( .din1(din1[26:24]), .din2(din2[26:24]), 
        .din2_din1_nz(din2_din1_nz_26_24), .din2_din1_denorm(
        din2_din1_denorm_26_24) );
  fpu_denorm_3b_8 i_fpu_denorm_23_21 ( .din1(din1[23:21]), .din2(din2[23:21]), 
        .din2_din1_nz(din2_din1_nz_23_21), .din2_din1_denorm(
        din2_din1_denorm_23_21) );
  fpu_denorm_3b_7 i_fpu_denorm_20_18 ( .din1(din1[20:18]), .din2(din2[20:18]), 
        .din2_din1_nz(din2_din1_nz_20_18), .din2_din1_denorm(
        din2_din1_denorm_20_18) );
  fpu_denorm_3b_6 i_fpu_denorm_17_15 ( .din1(din1[17:15]), .din2(din2[17:15]), 
        .din2_din1_nz(din2_din1_nz_17_15), .din2_din1_denorm(
        din2_din1_denorm_17_15) );
  fpu_denorm_3b_5 i_fpu_denorm_14_12 ( .din1(din1[14:12]), .din2(din2[14:12]), 
        .din2_din1_nz(din2_din1_nz_14_12), .din2_din1_denorm(
        din2_din1_denorm_14_12) );
  fpu_denorm_3b_4 i_fpu_denorm_11_9 ( .din1(din1[11:9]), .din2(din2[11:9]), 
        .din2_din1_nz(din2_din1_nz_11_9), .din2_din1_denorm(
        din2_din1_denorm_11_9) );
  fpu_denorm_3b_3 i_fpu_denorm_8_6 ( .din1(din1[8:6]), .din2(din2[8:6]), 
        .din2_din1_nz(din2_din1_nz_8_6), .din2_din1_denorm(
        din2_din1_denorm_8_6) );
  fpu_denorm_3b_2 i_fpu_denorm_5_3 ( .din1(din1[5:3]), .din2(din2[5:3]), 
        .din2_din1_nz(din2_din1_nz_5_3), .din2_din1_denorm(
        din2_din1_denorm_5_3) );
  fpu_denorm_3b_1 i_fpu_denorm_2_0 ( .din1(din1[2:0]), .din2(din2[2:0]), 
        .din2_din1_nz(din2_din1_nz_2_0), .din2_din1_denorm(
        din2_din1_denorm_2_0) );
  fpu_denorm_3to1_0 i_fpu_denorm_53_45 ( .din2_din1_nz_hi(din2_din1_nz_53_51), 
        .din2_din1_denorm_hi(din2_din1_denorm_53_51), .din2_din1_nz_mid(
        din2_din1_nz_50_48), .din2_din1_denorm_mid(din2_din1_denorm_50_48), 
        .din2_din1_nz_lo(din2_din1_nz_47_45), .din2_din1_denorm_lo(
        din2_din1_denorm_47_45), .din2_din1_nz(din2_din1_nz_53_45), 
        .din2_din1_denorm(din2_din1_denorm_53_45) );
  fpu_denorm_3to1_7 i_fpu_denorm_44_36 ( .din2_din1_nz_hi(din2_din1_nz_44_42), 
        .din2_din1_denorm_hi(din2_din1_denorm_44_42), .din2_din1_nz_mid(
        din2_din1_nz_41_39), .din2_din1_denorm_mid(din2_din1_denorm_41_39), 
        .din2_din1_nz_lo(din2_din1_nz_38_36), .din2_din1_denorm_lo(
        din2_din1_denorm_38_36), .din2_din1_nz(din2_din1_nz_44_36), 
        .din2_din1_denorm(din2_din1_denorm_44_36) );
  fpu_denorm_3to1_6 i_fpu_denorm_35_27 ( .din2_din1_nz_hi(din2_din1_nz_35_33), 
        .din2_din1_denorm_hi(din2_din1_denorm_35_33), .din2_din1_nz_mid(
        din2_din1_nz_32_30), .din2_din1_denorm_mid(din2_din1_denorm_32_30), 
        .din2_din1_nz_lo(din2_din1_nz_29_27), .din2_din1_denorm_lo(
        din2_din1_denorm_29_27), .din2_din1_nz(din2_din1_nz_35_27), 
        .din2_din1_denorm(din2_din1_denorm_35_27) );
  fpu_denorm_3to1_5 i_fpu_denorm_26_18 ( .din2_din1_nz_hi(din2_din1_nz_26_24), 
        .din2_din1_denorm_hi(din2_din1_denorm_26_24), .din2_din1_nz_mid(
        din2_din1_nz_23_21), .din2_din1_denorm_mid(din2_din1_denorm_23_21), 
        .din2_din1_nz_lo(din2_din1_nz_20_18), .din2_din1_denorm_lo(
        din2_din1_denorm_20_18), .din2_din1_nz(din2_din1_nz_26_18), 
        .din2_din1_denorm(din2_din1_denorm_26_18) );
  fpu_denorm_3to1_4 i_fpu_denorm_17_9 ( .din2_din1_nz_hi(din2_din1_nz_17_15), 
        .din2_din1_denorm_hi(din2_din1_denorm_17_15), .din2_din1_nz_mid(
        din2_din1_nz_14_12), .din2_din1_denorm_mid(din2_din1_denorm_14_12), 
        .din2_din1_nz_lo(din2_din1_nz_11_9), .din2_din1_denorm_lo(
        din2_din1_denorm_11_9), .din2_din1_nz(din2_din1_nz_17_9), 
        .din2_din1_denorm(din2_din1_denorm_17_9) );
  fpu_denorm_3to1_3 i_fpu_denorm_8_0 ( .din2_din1_nz_hi(din2_din1_nz_8_6), 
        .din2_din1_denorm_hi(din2_din1_denorm_8_6), .din2_din1_nz_mid(
        din2_din1_nz_5_3), .din2_din1_denorm_mid(din2_din1_denorm_5_3), 
        .din2_din1_nz_lo(din2_din1_nz_2_0), .din2_din1_denorm_lo(
        din2_din1_denorm_2_0), .din2_din1_nz(din2_din1_nz_8_0), 
        .din2_din1_denorm(din2_din1_denorm_8_0) );
  fpu_denorm_3to1_2 i_fpu_denorm_53_27 ( .din2_din1_nz_hi(din2_din1_nz_53_45), 
        .din2_din1_denorm_hi(din2_din1_denorm_53_45), .din2_din1_nz_mid(
        din2_din1_nz_44_36), .din2_din1_denorm_mid(din2_din1_denorm_44_36), 
        .din2_din1_nz_lo(din2_din1_nz_35_27), .din2_din1_denorm_lo(
        din2_din1_denorm_35_27), .din2_din1_nz(din2_din1_nz_53_27), 
        .din2_din1_denorm(din2_din1_denorm_53_27) );
  fpu_denorm_3to1_1 i_fpu_denorm_26_0 ( .din2_din1_nz_hi(din2_din1_nz_26_18), 
        .din2_din1_denorm_hi(din2_din1_denorm_26_18), .din2_din1_nz_mid(
        din2_din1_nz_17_9), .din2_din1_denorm_mid(din2_din1_denorm_17_9), 
        .din2_din1_nz_lo(din2_din1_nz_8_0), .din2_din1_denorm_lo(
        din2_din1_denorm_8_0), .din2_din1_nz(din2_din1_nz_26_0), 
        .din2_din1_denorm(din2_din1_denorm_26_0) );
  INVX1_RVT U1 ( .A(din2_din1_nz_53_27), .Y(n2) );
  INVX1_RVT U2 ( .A(din2_din1_nz_26_0), .Y(n1) );
  AO222X1_RVT U3 ( .A1(n2), .A2(din2_din1_denorm_26_0), .A3(n2), .A4(n1), .A5(
        din2_din1_denorm_53_27), .A6(din2_din1_nz_53_27), .Y(din2_din1_denorm)
         );
  INVX1_RVT U4 ( .A(din2_din1_denorm), .Y(din2_din1_denorm_inva) );
endmodule


module fpu_cnt_lead0_lvl1_0 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl2_0 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl3_0 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl4_0 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_16_eq_0), .A2(din_15_0_eq_0), .Y(din_31_0_eq_0)
         );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(din_15_8_eq_0), .A3(n1), .A4(
        din_31_24_eq_0), .Y(lead0_32b_3) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U6 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl4_7 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_16_eq_0), .A2(din_15_0_eq_0), .Y(din_31_0_eq_0)
         );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(din_15_8_eq_0), .A3(n1), .A4(
        din_31_24_eq_0), .Y(lead0_32b_3) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U6 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl3_10 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_11 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_12 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl1_40 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_41 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_42 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_43 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_44 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_45 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_46 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_47 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_48 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_49 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_50 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_51 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_52 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_53 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_54 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl2_19 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_20 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_21 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_22 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_23 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_24 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_25 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_64b ( din, lead0 );
  input [63:0] din;
  output [5:0] lead0;
  wire   din_63_60_eq_0, din_63_62_eq_0, lead0_63_60_0, din_59_56_eq_0,
         din_59_58_eq_0, lead0_59_56_0, din_55_52_eq_0, din_55_54_eq_0,
         lead0_55_52_0, din_51_48_eq_0, din_51_50_eq_0, lead0_51_48_0,
         din_47_44_eq_0, din_47_46_eq_0, lead0_47_44_0, din_43_40_eq_0,
         din_43_42_eq_0, lead0_43_40_0, din_39_36_eq_0, din_39_38_eq_0,
         lead0_39_36_0, din_35_32_eq_0, din_35_34_eq_0, lead0_35_32_0,
         din_31_28_eq_0, din_31_30_eq_0, lead0_31_28_0, din_27_24_eq_0,
         din_27_26_eq_0, lead0_27_24_0, din_23_20_eq_0, din_23_22_eq_0,
         lead0_23_20_0, din_19_16_eq_0, din_19_18_eq_0, lead0_19_16_0,
         din_15_12_eq_0, din_15_14_eq_0, lead0_15_12_0, din_11_8_eq_0,
         din_11_10_eq_0, lead0_11_8_0, din_7_4_eq_0, din_7_6_eq_0, lead0_7_4_0,
         din_3_0_eq_0, din_3_2_eq_0, lead0_3_0_0, din_63_56_eq_0,
         lead0_63_56_1, lead0_63_56_0, din_55_48_eq_0, lead0_55_48_1,
         lead0_55_48_0, din_47_40_eq_0, lead0_47_40_1, lead0_47_40_0,
         din_39_32_eq_0, lead0_39_32_1, lead0_39_32_0, din_31_24_eq_0,
         lead0_31_24_1, lead0_31_24_0, din_23_16_eq_0, lead0_23_16_1,
         lead0_23_16_0, din_15_8_eq_0, lead0_15_8_1, lead0_15_8_0,
         din_7_0_eq_0, lead0_7_0_1, lead0_7_0_0, din_63_48_eq_0, lead0_63_48_2,
         lead0_63_48_1, lead0_63_48_0, din_47_32_eq_0, lead0_47_32_2,
         lead0_47_32_1, lead0_47_32_0, din_31_16_eq_0, lead0_31_16_2,
         lead0_31_16_1, lead0_31_16_0, din_15_0_eq_0, lead0_15_0_2,
         lead0_15_0_1, lead0_15_0_0, din_63_32_eq_0, lead0_63_32_3,
         lead0_63_32_2, lead0_63_32_1, lead0_63_32_0, din_31_0_eq_0,
         lead0_31_0_3, lead0_31_0_2, lead0_31_0_1, lead0_31_0_0, n1;

  fpu_cnt_lead0_lvl1_0 i_fpu_cnt_lead0_lvl1_63_60 ( .din(din[63:60]), 
        .din_3_0_eq_0(din_63_60_eq_0), .din_3_2_eq_0(din_63_62_eq_0), 
        .lead0_4b_0(lead0_63_60_0) );
  fpu_cnt_lead0_lvl1_54 i_fpu_cnt_lead0_lvl1_59_56 ( .din(din[59:56]), 
        .din_3_0_eq_0(din_59_56_eq_0), .din_3_2_eq_0(din_59_58_eq_0), 
        .lead0_4b_0(lead0_59_56_0) );
  fpu_cnt_lead0_lvl1_53 i_fpu_cnt_lead0_lvl1_55_52 ( .din(din[55:52]), 
        .din_3_0_eq_0(din_55_52_eq_0), .din_3_2_eq_0(din_55_54_eq_0), 
        .lead0_4b_0(lead0_55_52_0) );
  fpu_cnt_lead0_lvl1_52 i_fpu_cnt_lead0_lvl1_51_48 ( .din(din[51:48]), 
        .din_3_0_eq_0(din_51_48_eq_0), .din_3_2_eq_0(din_51_50_eq_0), 
        .lead0_4b_0(lead0_51_48_0) );
  fpu_cnt_lead0_lvl1_51 i_fpu_cnt_lead0_lvl1_47_44 ( .din(din[47:44]), 
        .din_3_0_eq_0(din_47_44_eq_0), .din_3_2_eq_0(din_47_46_eq_0), 
        .lead0_4b_0(lead0_47_44_0) );
  fpu_cnt_lead0_lvl1_50 i_fpu_cnt_lead0_lvl1_43_40 ( .din(din[43:40]), 
        .din_3_0_eq_0(din_43_40_eq_0), .din_3_2_eq_0(din_43_42_eq_0), 
        .lead0_4b_0(lead0_43_40_0) );
  fpu_cnt_lead0_lvl1_49 i_fpu_cnt_lead0_lvl1_39_36 ( .din(din[39:36]), 
        .din_3_0_eq_0(din_39_36_eq_0), .din_3_2_eq_0(din_39_38_eq_0), 
        .lead0_4b_0(lead0_39_36_0) );
  fpu_cnt_lead0_lvl1_48 i_fpu_cnt_lead0_lvl1_35_32 ( .din(din[35:32]), 
        .din_3_0_eq_0(din_35_32_eq_0), .din_3_2_eq_0(din_35_34_eq_0), 
        .lead0_4b_0(lead0_35_32_0) );
  fpu_cnt_lead0_lvl1_47 i_fpu_cnt_lead0_lvl1_31_28 ( .din(din[31:28]), 
        .din_3_0_eq_0(din_31_28_eq_0), .din_3_2_eq_0(din_31_30_eq_0), 
        .lead0_4b_0(lead0_31_28_0) );
  fpu_cnt_lead0_lvl1_46 i_fpu_cnt_lead0_lvl1_27_24 ( .din(din[27:24]), 
        .din_3_0_eq_0(din_27_24_eq_0), .din_3_2_eq_0(din_27_26_eq_0), 
        .lead0_4b_0(lead0_27_24_0) );
  fpu_cnt_lead0_lvl1_45 i_fpu_cnt_lead0_lvl1_23_20 ( .din(din[23:20]), 
        .din_3_0_eq_0(din_23_20_eq_0), .din_3_2_eq_0(din_23_22_eq_0), 
        .lead0_4b_0(lead0_23_20_0) );
  fpu_cnt_lead0_lvl1_44 i_fpu_cnt_lead0_lvl1_19_16 ( .din(din[19:16]), 
        .din_3_0_eq_0(din_19_16_eq_0), .din_3_2_eq_0(din_19_18_eq_0), 
        .lead0_4b_0(lead0_19_16_0) );
  fpu_cnt_lead0_lvl1_43 i_fpu_cnt_lead0_lvl1_15_12 ( .din(din[15:12]), 
        .din_3_0_eq_0(din_15_12_eq_0), .din_3_2_eq_0(din_15_14_eq_0), 
        .lead0_4b_0(lead0_15_12_0) );
  fpu_cnt_lead0_lvl1_42 i_fpu_cnt_lead0_lvl1_11_8 ( .din(din[11:8]), 
        .din_3_0_eq_0(din_11_8_eq_0), .din_3_2_eq_0(din_11_10_eq_0), 
        .lead0_4b_0(lead0_11_8_0) );
  fpu_cnt_lead0_lvl1_41 i_fpu_cnt_lead0_lvl1_7_4 ( .din(din[7:4]), 
        .din_3_0_eq_0(din_7_4_eq_0), .din_3_2_eq_0(din_7_6_eq_0), .lead0_4b_0(
        lead0_7_4_0) );
  fpu_cnt_lead0_lvl1_40 i_fpu_cnt_lead0_lvl1_3_0 ( .din(din[3:0]), 
        .din_3_0_eq_0(din_3_0_eq_0), .din_3_2_eq_0(din_3_2_eq_0), .lead0_4b_0(
        lead0_3_0_0) );
  fpu_cnt_lead0_lvl2_0 i_fpu_cnt_lead0_lvl2_63_56 ( .din_7_4_eq_0(
        din_63_60_eq_0), .din_7_6_eq_0(din_63_62_eq_0), .lead0_4b_0_hi(
        lead0_63_60_0), .din_3_0_eq_0(din_59_56_eq_0), .din_3_2_eq_0(
        din_59_58_eq_0), .lead0_4b_0_lo(lead0_59_56_0), .din_7_0_eq_0(
        din_63_56_eq_0), .lead0_8b_1(lead0_63_56_1), .lead0_8b_0(lead0_63_56_0) );
  fpu_cnt_lead0_lvl2_25 i_fpu_cnt_lead0_lvl2_55_48 ( .din_7_4_eq_0(
        din_55_52_eq_0), .din_7_6_eq_0(din_55_54_eq_0), .lead0_4b_0_hi(
        lead0_55_52_0), .din_3_0_eq_0(din_51_48_eq_0), .din_3_2_eq_0(
        din_51_50_eq_0), .lead0_4b_0_lo(lead0_51_48_0), .din_7_0_eq_0(
        din_55_48_eq_0), .lead0_8b_1(lead0_55_48_1), .lead0_8b_0(lead0_55_48_0) );
  fpu_cnt_lead0_lvl2_24 i_fpu_cnt_lead0_lvl2_47_40 ( .din_7_4_eq_0(
        din_47_44_eq_0), .din_7_6_eq_0(din_47_46_eq_0), .lead0_4b_0_hi(
        lead0_47_44_0), .din_3_0_eq_0(din_43_40_eq_0), .din_3_2_eq_0(
        din_43_42_eq_0), .lead0_4b_0_lo(lead0_43_40_0), .din_7_0_eq_0(
        din_47_40_eq_0), .lead0_8b_1(lead0_47_40_1), .lead0_8b_0(lead0_47_40_0) );
  fpu_cnt_lead0_lvl2_23 i_fpu_cnt_lead0_lvl2_39_32 ( .din_7_4_eq_0(
        din_39_36_eq_0), .din_7_6_eq_0(din_39_38_eq_0), .lead0_4b_0_hi(
        lead0_39_36_0), .din_3_0_eq_0(din_35_32_eq_0), .din_3_2_eq_0(
        din_35_34_eq_0), .lead0_4b_0_lo(lead0_35_32_0), .din_7_0_eq_0(
        din_39_32_eq_0), .lead0_8b_1(lead0_39_32_1), .lead0_8b_0(lead0_39_32_0) );
  fpu_cnt_lead0_lvl2_22 i_fpu_cnt_lead0_lvl2_31_24 ( .din_7_4_eq_0(
        din_31_28_eq_0), .din_7_6_eq_0(din_31_30_eq_0), .lead0_4b_0_hi(
        lead0_31_28_0), .din_3_0_eq_0(din_27_24_eq_0), .din_3_2_eq_0(
        din_27_26_eq_0), .lead0_4b_0_lo(lead0_27_24_0), .din_7_0_eq_0(
        din_31_24_eq_0), .lead0_8b_1(lead0_31_24_1), .lead0_8b_0(lead0_31_24_0) );
  fpu_cnt_lead0_lvl2_21 i_fpu_cnt_lead0_lvl2_23_16 ( .din_7_4_eq_0(
        din_23_20_eq_0), .din_7_6_eq_0(din_23_22_eq_0), .lead0_4b_0_hi(
        lead0_23_20_0), .din_3_0_eq_0(din_19_16_eq_0), .din_3_2_eq_0(
        din_19_18_eq_0), .lead0_4b_0_lo(lead0_19_16_0), .din_7_0_eq_0(
        din_23_16_eq_0), .lead0_8b_1(lead0_23_16_1), .lead0_8b_0(lead0_23_16_0) );
  fpu_cnt_lead0_lvl2_20 i_fpu_cnt_lead0_lvl2_15_8 ( .din_7_4_eq_0(
        din_15_12_eq_0), .din_7_6_eq_0(din_15_14_eq_0), .lead0_4b_0_hi(
        lead0_15_12_0), .din_3_0_eq_0(din_11_8_eq_0), .din_3_2_eq_0(
        din_11_10_eq_0), .lead0_4b_0_lo(lead0_11_8_0), .din_7_0_eq_0(
        din_15_8_eq_0), .lead0_8b_1(lead0_15_8_1), .lead0_8b_0(lead0_15_8_0)
         );
  fpu_cnt_lead0_lvl2_19 i_fpu_cnt_lead0_lvl2_7_0 ( .din_7_4_eq_0(din_7_4_eq_0), 
        .din_7_6_eq_0(din_7_6_eq_0), .lead0_4b_0_hi(lead0_7_4_0), 
        .din_3_0_eq_0(din_3_0_eq_0), .din_3_2_eq_0(din_3_2_eq_0), 
        .lead0_4b_0_lo(lead0_3_0_0), .din_7_0_eq_0(din_7_0_eq_0), .lead0_8b_1(
        lead0_7_0_1), .lead0_8b_0(lead0_7_0_0) );
  fpu_cnt_lead0_lvl3_0 i_fpu_cnt_lead0_lvl3_63_48 ( .din_15_8_eq_0(
        din_63_56_eq_0), .din_15_12_eq_0(din_63_60_eq_0), .lead0_8b_1_hi(
        lead0_63_56_1), .lead0_8b_0_hi(lead0_63_56_0), .din_7_0_eq_0(
        din_55_48_eq_0), .din_7_4_eq_0(din_55_52_eq_0), .lead0_8b_1_lo(
        lead0_55_48_1), .lead0_8b_0_lo(lead0_55_48_0), .din_15_0_eq_0(
        din_63_48_eq_0), .lead0_16b_2(lead0_63_48_2), .lead0_16b_1(
        lead0_63_48_1), .lead0_16b_0(lead0_63_48_0) );
  fpu_cnt_lead0_lvl3_12 i_fpu_cnt_lead0_lvl3_47_32 ( .din_15_8_eq_0(
        din_47_40_eq_0), .din_15_12_eq_0(din_47_44_eq_0), .lead0_8b_1_hi(
        lead0_47_40_1), .lead0_8b_0_hi(lead0_47_40_0), .din_7_0_eq_0(
        din_39_32_eq_0), .din_7_4_eq_0(din_39_36_eq_0), .lead0_8b_1_lo(
        lead0_39_32_1), .lead0_8b_0_lo(lead0_39_32_0), .din_15_0_eq_0(
        din_47_32_eq_0), .lead0_16b_2(lead0_47_32_2), .lead0_16b_1(
        lead0_47_32_1), .lead0_16b_0(lead0_47_32_0) );
  fpu_cnt_lead0_lvl3_11 i_fpu_cnt_lead0_lvl3_31_16 ( .din_15_8_eq_0(
        din_31_24_eq_0), .din_15_12_eq_0(din_31_28_eq_0), .lead0_8b_1_hi(
        lead0_31_24_1), .lead0_8b_0_hi(lead0_31_24_0), .din_7_0_eq_0(
        din_23_16_eq_0), .din_7_4_eq_0(din_23_20_eq_0), .lead0_8b_1_lo(
        lead0_23_16_1), .lead0_8b_0_lo(lead0_23_16_0), .din_15_0_eq_0(
        din_31_16_eq_0), .lead0_16b_2(lead0_31_16_2), .lead0_16b_1(
        lead0_31_16_1), .lead0_16b_0(lead0_31_16_0) );
  fpu_cnt_lead0_lvl3_10 i_fpu_cnt_lead0_lvl3_15_0 ( .din_15_8_eq_0(
        din_15_8_eq_0), .din_15_12_eq_0(din_15_12_eq_0), .lead0_8b_1_hi(
        lead0_15_8_1), .lead0_8b_0_hi(lead0_15_8_0), .din_7_0_eq_0(
        din_7_0_eq_0), .din_7_4_eq_0(din_7_4_eq_0), .lead0_8b_1_lo(lead0_7_0_1), .lead0_8b_0_lo(lead0_7_0_0), .din_15_0_eq_0(din_15_0_eq_0), .lead0_16b_2(
        lead0_15_0_2), .lead0_16b_1(lead0_15_0_1), .lead0_16b_0(lead0_15_0_0)
         );
  fpu_cnt_lead0_lvl4_0 i_fpu_cnt_lead0_lvl4_63_32 ( .din_31_16_eq_0(
        din_63_48_eq_0), .din_31_24_eq_0(din_63_56_eq_0), .lead0_16b_2_hi(
        lead0_63_48_2), .lead0_16b_1_hi(lead0_63_48_1), .lead0_16b_0_hi(
        lead0_63_48_0), .din_15_0_eq_0(din_47_32_eq_0), .din_15_8_eq_0(
        din_47_40_eq_0), .lead0_16b_2_lo(lead0_47_32_2), .lead0_16b_1_lo(
        lead0_47_32_1), .lead0_16b_0_lo(lead0_47_32_0), .din_31_0_eq_0(
        din_63_32_eq_0), .lead0_32b_3(lead0_63_32_3), .lead0_32b_2(
        lead0_63_32_2), .lead0_32b_1(lead0_63_32_1), .lead0_32b_0(
        lead0_63_32_0) );
  fpu_cnt_lead0_lvl4_7 i_fpu_cnt_lead0_lvl4_31_0 ( .din_31_16_eq_0(
        din_31_16_eq_0), .din_31_24_eq_0(din_31_24_eq_0), .lead0_16b_2_hi(
        lead0_31_16_2), .lead0_16b_1_hi(lead0_31_16_1), .lead0_16b_0_hi(
        lead0_31_16_0), .din_15_0_eq_0(din_15_0_eq_0), .din_15_8_eq_0(
        din_15_8_eq_0), .lead0_16b_2_lo(lead0_15_0_2), .lead0_16b_1_lo(
        lead0_15_0_1), .lead0_16b_0_lo(lead0_15_0_0), .din_31_0_eq_0(
        din_31_0_eq_0), .lead0_32b_3(lead0_31_0_3), .lead0_32b_2(lead0_31_0_2), 
        .lead0_32b_1(lead0_31_0_1), .lead0_32b_0(lead0_31_0_0) );
  INVX1_RVT U1 ( .A(din_63_32_eq_0), .Y(n1) );
  NOR2X0_RVT U2 ( .A1(din_31_0_eq_0), .A2(n1), .Y(lead0[5]) );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(lead0[5]), .A3(din_63_48_eq_0), 
        .A4(n1), .Y(lead0[4]) );
  AO22X1_RVT U4 ( .A1(lead0_31_0_3), .A2(lead0[5]), .A3(lead0_63_32_3), .A4(n1), .Y(lead0[3]) );
  AO22X1_RVT U5 ( .A1(lead0_31_0_2), .A2(lead0[5]), .A3(lead0_63_32_2), .A4(n1), .Y(lead0[2]) );
  AO22X1_RVT U6 ( .A1(lead0_31_0_1), .A2(lead0[5]), .A3(lead0_63_32_1), .A4(n1), .Y(lead0[1]) );
  AO22X1_RVT U7 ( .A1(lead0_31_0_0), .A2(lead0[5]), .A3(lead0_63_32_0), .A4(n1), .Y(lead0[0]) );
endmodule


module clken_buf_10 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE63 ( din, en, clk, q, se, si, so );
  input [62:0] din;
  output [62:0] q;
  input [62:0] si;
  output [62:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, net24534, n3, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE63 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24534), .TE(1'b0) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24534), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24534), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24534), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24534), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24534), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24534), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24534), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24534), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24534), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24534), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24534), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24534), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24534), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24534), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24534), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24534), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24534), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24534), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24534), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24534), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24534), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24534), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24534), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24534), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24534), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24534), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24534), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24534), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24534), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24534), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24534), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24534), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24534), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24534), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24534), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24534), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24534), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24534), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24534), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24534), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24534), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24534), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24534), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24534), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24534), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24534), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24534), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24534), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24534), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24534), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24534), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24534), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24534), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24534), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24534), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24534), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24534), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24534), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24534), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24534), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24534), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24534), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24534), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n6) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n6), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n6), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n6), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n6), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n6), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n6), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n6), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n6), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n6), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n6), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n6), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n6), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n5), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n6), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n5), .Y(N66) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_0 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n3, n1, n2, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_0 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n3, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n5), .Y(N63) );
  INVX1_RVT U66 ( .A(se), .Y(n6) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n6), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n6), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n6), .Y(N66) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n6), .Y(N67) );
  OR2X1_RVT U72 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_10 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_10 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_9 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_9 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n5), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[60]), .A2(n1), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[61]), .A2(n2), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[62]), .A2(n4), .Y(N66) );
  AND2X1_RVT U69 ( .A1(din[63]), .A2(n5), .Y(N67) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_8 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6, n7;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_8 clk_gate_q_reg ( .CLK(clk), .EN(n7), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n6) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n6), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n6), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n6), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n6), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n6), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n6), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n6), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n6), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n6), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n6), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n6), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n6), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n5), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n6), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n5), .Y(N66) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n6), .Y(N67) );
  OR2X1_RVT U72 ( .A1(se), .A2(en), .Y(n7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_7 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6, n7;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_7 clk_gate_q_reg ( .CLK(clk), .EN(n7), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n6) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n6), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n6), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n6), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n6), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n6), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n6), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n6), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n6), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n6), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n6), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n6), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n6), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n2), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n4), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n5), .Y(N66) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n6), .Y(N67) );
  OR2X1_RVT U72 ( .A1(se), .A2(en), .Y(n7) );
endmodule


module dff_SIZE64_5 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n3), .Y(N57) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n4), .Y(N58) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n2), .Y(N60) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n3), .Y(N61) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n4), .Y(N62) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n2), .Y(N64) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n3), .Y(N65) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n4), .Y(N66) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_6 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, net24480, n1, n2, n4, n5, n6, n7;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_6 clk_gate_q_reg ( .CLK(clk), .EN(n7), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U29 ( .A(se), .Y(n4) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U42 ( .A(se), .Y(n5) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n5), .Y(N63) );
  INVX1_RVT U67 ( .A(se), .Y(n6) );
  AND2X1_RVT U68 ( .A1(din[60]), .A2(n6), .Y(N64) );
  AND2X1_RVT U69 ( .A1(din[61]), .A2(n6), .Y(N65) );
  AND2X1_RVT U70 ( .A1(din[62]), .A2(n6), .Y(N66) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_5 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_5 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n5), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[60]), .A2(n1), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[61]), .A2(n2), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[62]), .A2(n4), .Y(N66) );
  AND2X1_RVT U69 ( .A1(din[63]), .A2(n5), .Y(N67) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE54 ( din, en, clk, q, se, si, so );
  input [53:0] din;
  output [53:0] q;
  input [53:0] si;
  output [53:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, net24516, n3,
         n1, n2, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE54 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24516), .TE(1'b0) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24516), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24516), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24516), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24516), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24516), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24516), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24516), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24516), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24516), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24516), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24516), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24516), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24516), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24516), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24516), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24516), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24516), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24516), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24516), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24516), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24516), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24516), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24516), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24516), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24516), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24516), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24516), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24516), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24516), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24516), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24516), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24516), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24516), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24516), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24516), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24516), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24516), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24516), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24516), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24516), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24516), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24516), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24516), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24516), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24516), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24516), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24516), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24516), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24516), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24516), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24516), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24516), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24516), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24516), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n2), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n4), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n5), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n2), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n4), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n5), .Y(N57) );
  OR2X1_RVT U61 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_4 ( din, en, clk, se, si, so, \q[63] , \q[62] , \q[61] , 
        \q[60] , \q[59] , \q[58] , \q[57] , \q[56] , \q[55] , \q[54] , \q[53] , 
        \q[52] , \q[51] , \q[50] , \q[49] , \q[48] , \q[47] , \q[44] , \q[43] , 
        \q[42] , \q[41] , \q[40] , \q[39] , \q[38] , \q[37] , \q[36]_BAR , 
        \q[35] , \q[32] , \q[31] , \q[29] , \q[28] , \q[27] , \q[26] , \q[25] , 
        \q[24] , \q[23] , \q[22] , \q[21] , \q[20] , \q[19] , \q[18] , \q[17] , 
        \q[16] , \q[15] , \q[14] , \q[13] , \q[12] , \q[11] , \q[10] , \q[9] , 
        \q[8] , \q[7] , \q[6] , \q[5] , \q[4] , \q[3] , \q[2] , \q[1] , \q[0] , 
        \q[46]_BAR , \q[45]_BAR , \q[34]_BAR , \q[33]_BAR , \q[30]_BAR  );
  input [63:0] din;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  output \q[63] , \q[62] , \q[61] , \q[60] , \q[59] , \q[58] , \q[57] ,
         \q[56] , \q[55] , \q[54] , \q[53] , \q[52] , \q[51] , \q[50] ,
         \q[49] , \q[48] , \q[47] , \q[44] , \q[43] , \q[42] , \q[41] ,
         \q[40] , \q[39] , \q[38] , \q[37] , \q[36]_BAR , \q[35] , \q[32] ,
         \q[31] , \q[29] , \q[28] , \q[27] , \q[26] , \q[25] , \q[24] ,
         \q[23] , \q[22] , \q[21] , \q[20] , \q[19] , \q[18] , \q[17] ,
         \q[16] , \q[15] , \q[14] , \q[13] , \q[12] , \q[11] , \q[10] , \q[9] ,
         \q[8] , \q[7] , \q[6] , \q[5] , \q[4] , \q[3] , \q[2] , \q[1] ,
         \q[0] , \q[46]_BAR , \q[45]_BAR , \q[34]_BAR , \q[33]_BAR ,
         \q[30]_BAR ;
  wire   N4, N6, N8, N9, N10, N11, N12, N16, N17, N18, N19, N20, N21, N22, N25,
         N28, N31, N34, N36, N38, N40, N44, N45, N46, N64, net24480, n1, n2,
         n10;
  wire   [63:0] q;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_4 clk_gate_q_reg ( .CLK(clk), .EN(n10), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N64), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N64), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N46), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N46), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N46), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[52]  ( .D(N45), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N45), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N45), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N45), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N45), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N44), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N44), .CLK(net24480), .QN(\q[46]_BAR ) );
  DFFX1_RVT \q_reg[45]  ( .D(N44), .CLK(net24480), .QN(\q[45]_BAR ) );
  DFFX1_RVT \q_reg[44]  ( .D(N44), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N44), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N38), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N36), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N34), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .QN(\q[36]_BAR ) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .QN(\q[34]_BAR ) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(net24480), .QN(\q[33]_BAR ) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .QN(\q[30]_BAR ) );
  DFFX1_RVT \q_reg[29]  ( .D(N31), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(din[42]), .Y(N64) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U7 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U8 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U9 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U10 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U11 ( .A1(din[12]), .A2(n1), .Y(N16) );
  AND2X1_RVT U12 ( .A1(din[13]), .A2(n1), .Y(N17) );
  AND2X1_RVT U13 ( .A1(din[14]), .A2(n1), .Y(N18) );
  AND2X1_RVT U14 ( .A1(din[15]), .A2(n1), .Y(N19) );
  AND2X1_RVT U15 ( .A1(din[16]), .A2(n1), .Y(N20) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U18 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U19 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U20 ( .A1(din[24]), .A2(n2), .Y(N28) );
  AND2X1_RVT U21 ( .A1(din[27]), .A2(n2), .Y(N31) );
  AND2X1_RVT U22 ( .A1(din[30]), .A2(n2), .Y(N34) );
  AND2X1_RVT U23 ( .A1(din[32]), .A2(n2), .Y(N36) );
  AND2X1_RVT U24 ( .A1(din[34]), .A2(n2), .Y(N38) );
  AND2X1_RVT U25 ( .A1(din[36]), .A2(n2), .Y(N40) );
  AND2X1_RVT U26 ( .A1(din[40]), .A2(n2), .Y(N44) );
  AND2X1_RVT U27 ( .A1(din[41]), .A2(n2), .Y(N45) );
  AND2X1_RVT U28 ( .A1(din[42]), .A2(n2), .Y(N46) );
  OR2X1_RVT U30 ( .A1(se), .A2(en), .Y(n10) );
endmodule


module dff_SIZE64_4 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61,
         N62, N63, N64, N65, N66, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[13]), .A2(n1), .Y(N16) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[23]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[24]), .A2(n2), .Y(N27) );
  AND2X1_RVT U28 ( .A1(din[25]), .A2(n2), .Y(N28) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n3), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n3), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n3), .Y(N40) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[48]), .A2(n4), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[49]), .A2(n4), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[54]), .A2(n3), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[55]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[57]), .A2(n2), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[58]), .A2(n3), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[59]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[61]), .A2(n2), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[63]), .A2(n2), .Y(N66) );
endmodule


module dff_SIZE64_3 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N15) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n2), .Y(N27) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n3), .Y(N38) );
  AND2X1_RVT U41 ( .A1(din[36]), .A2(n3), .Y(N39) );
  AND2X1_RVT U42 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[38]), .A2(n2), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[39]), .A2(n3), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[41]), .A2(n2), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[42]), .A2(n3), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[44]), .A2(n2), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[45]), .A2(n3), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[47]), .A2(n2), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[48]), .A2(n3), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n4) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n4), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n4), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n4), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n4), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n4), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n4), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n4), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[60]), .A2(n4), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[61]), .A2(n4), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[62]), .A2(n4), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[63]), .A2(n4), .Y(N66) );
endmodule


module dff_SIZE64_2 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n3), .Y(N57) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n4), .Y(N58) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n2), .Y(N60) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n3), .Y(N61) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n4), .Y(N62) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n2), .Y(N64) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n3), .Y(N65) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n4), .Y(N66) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_3 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_3 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n5), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[60]), .A2(n1), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[61]), .A2(n2), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[62]), .A2(n4), .Y(N66) );
  AND2X1_RVT U69 ( .A1(din[63]), .A2(n5), .Y(N67) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE58 ( din, en, clk, q, se, si, so );
  input [57:0] din;
  output [57:0] q;
  input [57:0] si;
  output [57:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, net24498, n3, n1, n2, n4, n5;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE58 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24498), .TE(1'b0) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24498), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24498), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24498), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24498), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24498), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24498), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24498), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24498), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24498), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24498), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24498), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24498), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24498), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24498), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24498), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24498), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24498), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24498), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24498), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24498), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24498), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24498), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24498), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24498), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24498), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24498), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24498), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24498), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24498), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24498), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24498), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24498), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24498), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24498), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24498), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24498), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24498), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24498), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24498), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24498), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24498), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24498), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24498), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24498), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24498), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24498), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24498), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24498), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24498), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24498), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24498), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24498), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24498), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24498), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24498), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24498), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24498), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24498), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  OR2X1_RVT U65 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_2 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_2 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[55]), .A2(n5), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[56]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[57]), .A2(n2), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[58]), .A2(n4), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[59]), .A2(n5), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[60]), .A2(n1), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[61]), .A2(n2), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[62]), .A2(n4), .Y(N66) );
  AND2X1_RVT U69 ( .A1(din[63]), .A2(n5), .Y(N67) );
  OR2X1_RVT U71 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE64_1 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, net24480, n1, n2, n4, n5, n6, n7;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE64_1 clk_gate_q_reg ( .CLK(clk), .EN(n7), 
        .ENCLK(net24480), .TE(1'b0) );
  DFFX1_RVT \q_reg[63]  ( .D(N67), .CLK(net24480), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N66), .CLK(net24480), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N65), .CLK(net24480), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N64), .CLK(net24480), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N63), .CLK(net24480), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N62), .CLK(net24480), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N61), .CLK(net24480), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N60), .CLK(net24480), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N59), .CLK(net24480), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24480), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24480), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24480), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24480), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24480), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24480), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24480), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24480), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24480), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24480), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24480), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24480), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24480), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24480), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24480), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24480), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24480), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24480), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24480), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24480), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24480), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24480), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24480), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24480), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24480), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24480), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24480), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24480), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24480), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24480), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24480), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24480), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24480), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24480), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24480), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24480), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24480), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24480), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24480), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24480), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24480), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24480), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24480), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24480), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24480), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24480), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24480), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24480), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24480), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24480), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24480), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24480), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24480), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24480), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24480), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  INVX1_RVT U54 ( .A(se), .Y(n6) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n6), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n6), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n6), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n6), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n6), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n6), .Y(N57) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n6), .Y(N58) );
  AND2X1_RVT U62 ( .A1(din[55]), .A2(n6), .Y(N59) );
  AND2X1_RVT U63 ( .A1(din[56]), .A2(n6), .Y(N60) );
  AND2X1_RVT U64 ( .A1(din[57]), .A2(n6), .Y(N61) );
  AND2X1_RVT U65 ( .A1(din[58]), .A2(n6), .Y(N62) );
  AND2X1_RVT U66 ( .A1(din[59]), .A2(n6), .Y(N63) );
  AND2X1_RVT U67 ( .A1(din[60]), .A2(n2), .Y(N64) );
  AND2X1_RVT U68 ( .A1(din[61]), .A2(n4), .Y(N65) );
  AND2X1_RVT U69 ( .A1(din[62]), .A2(n5), .Y(N66) );
  AND2X1_RVT U70 ( .A1(din[63]), .A2(n6), .Y(N67) );
  OR2X1_RVT U72 ( .A1(se), .A2(en), .Y(n7) );
endmodule


module fpu_add_frac_dp ( inq_in1, inq_in2, a1stg_step, a1stg_sngop, 
        a1stg_expadd3_11, a1stg_norm_dbl_in1, a1stg_denorm_dbl_in1, 
        a1stg_norm_sng_in1, a1stg_denorm_sng_in1, a1stg_norm_dbl_in2, 
        a1stg_denorm_dbl_in2, a1stg_norm_sng_in2, a1stg_denorm_sng_in2, 
        a1stg_intlngop, a2stg_frac1_in_frac1, a2stg_frac1_in_frac2, 
        a1stg_2nan_in_inv, a1stg_faddsubop_inv, a2stg_frac1_in_qnan, 
        a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, a6stg_step, 
        a2stg_frac2_in_frac1, a2stg_frac2_in_qnan, a2stg_shr_cnt_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int, 
        a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max, 
        a2stg_expadd_11, a2stg_sub_step, a2stg_fracadd_frac2_inv_in, 
        a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2, 
        a2stg_fracadd_cin_in, a2stg_exp, a2stg_expdec_neq_0, a3stg_faddsubopa, 
        a3stg_sub_in, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, a3stg_exp_0, 
        a4stg_rnd_frac_add_inv, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, 
        a4stg_rnd_sng, a4stg_rnd_dbl, a4stg_shl_cnt_in, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0, 
        fadd_clken_l, rclk, a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, 
        a1stg_in2_eq_in1_exp, a2stg_frac2_63, a2stg_frac2hi_neq_0, 
        a2stg_frac2lo_neq_0, a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a3stg_denorm, 
        a3stg_denorm_inv, a3stg_lead0, a4stg_shl_cnt, a4stg_denorm_inv, 
        a3stg_inc_exp_inv, a3stg_same_exp_inv, a3stg_dec_exp_inv, 
        a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac_11, 
        a4stg_rnd_frac_10, a4stg_rndadd_cout, a4stg_frac_9_0_nx, 
        a4stg_frac_dbl_nx, a4stg_frac_38_0_nx, a4stg_frac_sng_nx, 
        a4stg_frac_neq_0, a4stg_shl_data_neq_0, add_of_out_cout, add_frac_out, 
        se, si, so, a4stg_round_BAR );
  input [62:0] inq_in1;
  input [63:0] inq_in2;
  input [5:0] a2stg_shr_cnt_in;
  input [5:0] a2stg_exp;
  input [1:0] a3stg_faddsubopa;
  input [9:0] a4stg_shl_cnt_in;
  output [5:0] a3stg_lead0;
  output [5:0] a4stg_shl_cnt;
  output [63:0] add_frac_out;
  input a1stg_step, a1stg_sngop, a1stg_expadd3_11, a1stg_norm_dbl_in1,
         a1stg_denorm_dbl_in1, a1stg_norm_sng_in1, a1stg_denorm_sng_in1,
         a1stg_norm_dbl_in2, a1stg_denorm_dbl_in2, a1stg_norm_sng_in2,
         a1stg_denorm_sng_in2, a1stg_intlngop, a2stg_frac1_in_frac1,
         a2stg_frac1_in_frac2, a1stg_2nan_in_inv, a1stg_faddsubop_inv,
         a2stg_frac1_in_qnan, a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl,
         a6stg_step, a2stg_frac2_in_frac1, a2stg_frac2_in_qnan,
         a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_expadd_11, a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a2stg_expdec_neq_0, a3stg_sub_in,
         a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, a3stg_exp_0,
         a4stg_rnd_frac_add_inv, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0,
         fadd_clken_l, rclk, se, si;
  output a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, a1stg_in2_eq_in1_exp,
         a2stg_frac2_63, a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0,
         a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a3stg_denorm, a3stg_denorm_inv,
         a4stg_denorm_inv, a3stg_inc_exp_inv, a3stg_same_exp_inv,
         a3stg_dec_exp_inv, a4stg_rnd_frac_40, a4stg_rnd_frac_39,
         a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_rndadd_cout,
         a4stg_frac_9_0_nx, a4stg_frac_dbl_nx, a4stg_frac_38_0_nx,
         a4stg_frac_sng_nx, a4stg_frac_neq_0, a4stg_shl_data_neq_0,
         add_of_out_cout, so, a4stg_round_BAR;
  wire   a4stg_round, clk, a1stg_in2_gt_in1, a2stg_fsdtoi_nx, a2stg_fsdtoix_nx,
         a2stg_fracadd_frac2_inv, a2stg_fracadd_frac2_inv_shr1,
         a2stg_fracadd_cin, a3stg_ld0_dnrm_10, a3stg_denorm_inva, a3stg_suba,
         \a4stg_shl_cnt_dec54_2[0] , \a4stg_shl_cnt_dec54_3[0] ,
         a4stg_round_in, a4stg_rnd_frac_63, a4stg_rnd_frac_62,
         a4stg_rnd_frac_61, a4stg_rnd_frac_60, a4stg_rnd_frac_59,
         a4stg_rnd_frac_58, a4stg_rnd_frac_57, a4stg_rnd_frac_56,
         a4stg_rnd_frac_55, a4stg_rnd_frac_54, a4stg_rnd_frac_53,
         a4stg_rnd_frac_52, a4stg_rnd_frac_51, a4stg_rnd_frac_50,
         a4stg_rnd_frac_49, a4stg_rnd_frac_48, a4stg_rnd_frac_47,
         a4stg_rnd_frac_46, a4stg_rnd_frac_45, a4stg_rnd_frac_44,
         a4stg_rnd_frac_43, a4stg_rnd_frac_42, a4stg_rnd_frac_41,
         a4stg_rnd_frac_9, a4stg_rnd_frac_8, a4stg_rnd_frac_7,
         a4stg_rnd_frac_6, a4stg_rnd_frac_5, a4stg_rnd_frac_4,
         a4stg_rnd_frac_3, a4stg_rnd_frac_2, a4stg_rnd_frac_1,
         a5stg_frac_out_rndadd, a5stg_frac_out_rnd_frac, a5stg_in_of,
         a5stg_frac_out_shl, a5stg_to_0, N1198, N1206, N1214, N1222, N1230,
         N1238, N1246, N1254, N1262, N1270, N1278, N1601, N1607, N1613, N1619,
         N1625, N1631, N1637, N1643, N1649, N1655, N1661, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, \DP_OP_16J2_123_4718/n1 , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2542, n2543;
  wire   [62:0] a1stg_in1;
  wire   [54:0] a1stg_in1a;
  wire   [63:0] a1stg_in2;
  wire   [54:0] a1stg_in2a;
  wire   [63:0] a2stg_frac1_in;
  wire   [63:0] a2stg_frac1;
  wire   [63:0] a2stg_frac2_in;
  wire   [62:0] a2stg_frac2;
  wire   [63:0] a2stg_frac2a;
  wire   [3:0] a2stg_shr_cnt_5;
  wire   [3:0] a2stg_shr_cnt_5_inv;
  wire   [4:0] a2stg_shr_cnt_4;
  wire   [4:0] a2stg_shr_cnt_3;
  wire   [1:0] a2stg_shr_cnt_2;
  wire   [1:0] a2stg_shr_cnt_1;
  wire   [1:0] a2stg_shr_cnt_0;
  wire   [5:0] a2stg_shr_cnt;
  wire   [63:0] a3stg_frac2;
  wire   [63:0] a3stg_frac1;
  wire   [63:0] a2stg_fracadd;
  wire   [63:0] a3stg_ld0_frac;
  wire   [53:0] a2stg_expdec;
  wire   [53:0] a3stg_expdec;
  wire   [2:0] a4stg_shl_cnt_dec54_0;
  wire   [2:0] a4stg_shl_cnt_dec54_1;
  wire   [63:2] a4stg_rnd_frac_pre1_in;
  wire   [63:0] a4stg_rnd_frac_pre1;
  wire   [63:1] a4stg_rnd_frac_pre3_in;
  wire   [63:0] a4stg_rnd_frac_pre3;
  wire   [63:0] a4stg_shl;
  wire   [38:12] a4stg_rnd_frac;
  wire   [63:0] a4stg_rnd_frac_pre2_in;
  wire   [63:0] a4stg_rnd_frac_pre2;
  wire   [63:0] a4stg_shl_data_in;
  wire   [63:0] a4stg_shl_data;
  wire   [51:0] a4stg_rndadd_tmp;
  wire   [51:0] a5stg_rndadd;
  wire   [63:0] a5stg_rnd_frac;
  wire   [63:0] a5stg_shl;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign a4stg_round_BAR = a4stg_round;
  assign so = 1'b0;

  clken_buf_10 ckbuf_add_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fadd_clken_l), .tmb_l(n2543) );
  dffe_SIZE63 i_a1stg_in1 ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_0 i_a1stg_in1a ( .din(inq_in1[54:0]), .en(a1stg_step), .clk(clk), 
        .q(a1stg_in1a), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_0 i_a1stg_in2 ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_10 i_a1stg_in2a ( .din(inq_in2[54:0]), .en(a1stg_step), .clk(clk), .q(a1stg_in2a), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  fpu_in2_gt_in1_frac i_a1stg_in2_gt_in1_frac ( .din1(a1stg_in1a), .din2(
        a1stg_in2a), .sngop(a1stg_sngop), .expadd11(a1stg_expadd3_11), .expeq(
        a1stg_in2_eq_in1_exp), .din2_neq_din1(a1stg_in2_neq_in1_frac), 
        .din2_gt_din1(a1stg_in2_gt_in1_frac), .din2_gt1_din1(a1stg_in2_gt_in1)
         );
  dffe_SIZE64_9 i_a2stg_frac1 ( .din({a2stg_frac1_in[63:11], N1198, N1206, 
        N1214, N1222, N1230, N1238, N1246, N1254, N1262, N1270, N1278}), .en(
        a6stg_step), .clk(clk), .q(a2stg_frac1), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dffe_SIZE64_8 i_a2stg_frac2 ( .din({a2stg_frac2_in[63:11], N1601, N1607, 
        N1613, N1619, N1625, N1631, N1637, N1643, N1649, N1655, N1661}), .en(
        a6stg_step), .clk(clk), .q({a2stg_frac2_63, a2stg_frac2}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_7 i_a2stg_frac2a ( .din({a2stg_frac2_in[63:11], N1601, N1607, 
        N1613, N1619, N1625, N1631, N1637, N1643, N1649, N1655, N1661}), .en(
        a6stg_step), .clk(clk), .q(a2stg_frac2a), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dff_SIZE64_5 i_a3stg_frac2 ( .din({n1731, n1730, n1729, n1728, n1727, n1726, 
        n1725, n1724, n1723, n1722, n1721, n1720, n1719, n1718, n1717, n1716, 
        n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, n1707, n1706, 
        n1705, n1704, n1703, n1702, n1701, n1700, n1699, n1698, n1697, n1696, 
        n1695, n1694, n1693, n1692, n1691, n1690, n1689, n1688, n1687, n1686, 
        n1685, n1684, n1683, n1682, n1681, n1680, n1679, n1678, n1677, n1676, 
        n1668, n1675, n1674, n1673, n1672, n1671, n1670, n1669}), .clk(clk), 
        .q({\DP_OP_16J2_123_4718/n1 , a3stg_frac2[62:0]}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_6 i_a3stg_frac1 ( .din({1'b0, a2stg_frac1[63:1]}), .en(
        a6stg_step), .clk(clk), .q({SYNOPSYS_UNCONNECTED__0, a3stg_frac1[62:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_5 i_a3stg_ld0_frac ( .din(a2stg_fracadd), .en(a6stg_step), .clk(
        clk), .q(a3stg_ld0_frac), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE54 i_a3stg_expdec ( .din(a2stg_expdec), .en(a6stg_step), .clk(clk), 
        .q(a3stg_expdec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  fpu_denorm_frac i_a3stg_denorm ( .din1({a3stg_ld0_frac[63:11], 
        a3stg_ld0_dnrm_10}), .din2(a3stg_expdec), .din2_din1_denorm(
        a3stg_denorm), .din2_din1_denorma(n5), .din2_din1_denorm_inva(
        a3stg_denorm_inva) );
  fpu_cnt_lead0_64b i_a3stg_lead0 ( .din(a3stg_ld0_frac), .lead0(a3stg_lead0)
         );
  dffe_SIZE64_4 i_astg_xtra_regs ( .din({a2stg_shr_cnt_5_inv_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_cnt_5_inv_in, a2stg_shr_cnt_5_inv_in, 
        a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], 1'b0, 
        1'b0, 1'b0, 1'b0, a2stg_shr_cnt_in[4], a2stg_shr_cnt_in[4], 
        a2stg_shr_cnt_in[4], a2stg_shr_cnt_in[4], a2stg_shr_cnt_in[4:3], 
        a2stg_shr_cnt_in[3], a2stg_shr_cnt_in[3], a2stg_shr_cnt_in[3], 
        a2stg_shr_cnt_in[3], a2stg_shr_cnt_in[5:3], 1'b0, 1'b0, 1'b0, 
        a4stg_round_in, 1'b0, a2stg_shr_cnt_in[2], 1'b0, a2stg_shr_cnt_in[1], 
        1'b0, a2stg_shr_cnt_in[0], 1'b0, 1'b0, a4stg_shl_cnt_in[6], 1'b0, 
        a4stg_shl_cnt_in[7], a4stg_shl_cnt_in[7], 1'b0, 1'b0, 
        a4stg_shl_cnt_in[8], 1'b0, 1'b0, a4stg_shl_cnt_in[9], 
        a4stg_shl_cnt_in[5:0], 1'b0, 1'b0, 1'b0, a2stg_fracadd_frac2_inv_in, 
        a2stg_fracadd_frac2_inv_shr1_in, a3stg_denorm_inva, a2stg_fsdtoix_nx, 
        a2stg_fsdtoi_nx, 1'b0, a2stg_fracadd_cin_in, 1'b0, a3stg_sub_in}), 
        .en(a6stg_step), .clk(clk), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .\q[63] (a2stg_shr_cnt_5_inv[3]), .\q[62] (a2stg_shr_cnt_5_inv[2]), 
        .\q[61] (a2stg_shr_cnt_5_inv[1]), .\q[60] (a2stg_shr_cnt_5_inv[0]), 
        .\q[59] (a2stg_shr_cnt_5[3]), .\q[58] (a2stg_shr_cnt_5[2]), .\q[57] (
        a2stg_shr_cnt_5[1]), .\q[52] (a2stg_shr_cnt_4[4]), .\q[51] (
        a2stg_shr_cnt_4[3]), .\q[50] (a2stg_shr_cnt_4[2]), .\q[49] (
        a2stg_shr_cnt_4[1]), .\q[48] (a2stg_shr_cnt_4[0]), .\q[47] (
        a2stg_shr_cnt_3[4]), .\q[44] (a2stg_shr_cnt_3[1]), .\q[43] (
        a2stg_shr_cnt_3[0]), .\q[42] (a2stg_shr_cnt[5]), .\q[41] (
        a2stg_shr_cnt[4]), .\q[40] (a2stg_shr_cnt[3]), .\q[39] (
        a2stg_shr_cnt[2]), .\q[38] (a2stg_shr_cnt[1]), .\q[37] (
        a2stg_shr_cnt[0]), .\q[36]_BAR (a4stg_round), .\q[35] (
        a2stg_shr_cnt_2[1]), .\q[32] (a2stg_shr_cnt_1[0]), .\q[31] (
        a2stg_shr_cnt_0[1]), .\q[29] (a4stg_shl_cnt_dec54_0[2]), .\q[28] (
        a4stg_shl_cnt_dec54_0[1]), .\q[27] (a4stg_shl_cnt_dec54_0[0]), 
        .\q[25] (a4stg_shl_cnt_dec54_1[1]), .\q[24] (a4stg_shl_cnt_dec54_1[0]), 
        .\q[21] (\a4stg_shl_cnt_dec54_2[0] ), .\q[18] (
        \a4stg_shl_cnt_dec54_3[0] ), .\q[17] (a4stg_shl_cnt[5]), .\q[16] (
        a4stg_shl_cnt[4]), .\q[15] (a4stg_shl_cnt[3]), .\q[14] (
        a4stg_shl_cnt[2]), .\q[13] (a4stg_shl_cnt[1]), .\q[12] (
        a4stg_shl_cnt[0]), .\q[8] (a2stg_fracadd_frac2_inv), .\q[7] (
        a2stg_fracadd_frac2_inv_shr1), .\q[6] (a4stg_denorm_inv), .\q[5] (
        a3stg_fsdtoix_nx), .\q[4] (a3stg_fsdtoi_nx), .\q[2] (a2stg_fracadd_cin), .\q[0] (a3stg_suba), .\q[46]_BAR (a2stg_shr_cnt_3[3]), .\q[45]_BAR (
        a2stg_shr_cnt_3[2]), .\q[34]_BAR (a2stg_shr_cnt_2[0]), .\q[33]_BAR (
        a2stg_shr_cnt_1[1]), .\q[30]_BAR (a2stg_shr_cnt_0[0]) );
  dff_SIZE64_4 i_a4stg_rnd_frac_pre1 ( .din({n2542, 
        a4stg_rnd_frac_pre1_in[62:2], 1'b0, 1'b0}), .clk(clk), .q({
        a4stg_rnd_frac_pre1[63:2], SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE64_3 i_a4stg_rnd_frac_pre3 ( .din({a4stg_rnd_frac_pre3_in, 1'b0}), 
        .clk(clk), .q({a4stg_rnd_frac_pre3[63:1], SYNOPSYS_UNCONNECTED__3}), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE64_2 i_a4stg_rnd_frac_pre2 ( .din(a4stg_rnd_frac_pre2_in), .clk(clk), 
        .q(a4stg_rnd_frac_pre2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_3 i_a4stg_shl_data ( .din(a4stg_shl_data_in), .en(a6stg_step), 
        .clk(clk), .q(a4stg_shl_data), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE58 i_a5stg_rndadd ( .din({a4stg_rndadd_cout, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0, 
        a4stg_rndadd_tmp}), .en(a6stg_step), .clk(clk), .q({add_of_out_cout, 
        a5stg_frac_out_rndadd, a5stg_frac_out_rnd_frac, a5stg_in_of, 
        a5stg_frac_out_shl, a5stg_to_0, a5stg_rndadd}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_2 i_a5stg_rnd_frac ( .din({a4stg_rnd_frac_63, a4stg_rnd_frac_62, 
        a4stg_rnd_frac_61, a4stg_rnd_frac_60, a4stg_rnd_frac_59, 
        a4stg_rnd_frac_58, a4stg_rnd_frac_57, a4stg_rnd_frac_56, 
        a4stg_rnd_frac_55, a4stg_rnd_frac_54, a4stg_rnd_frac_53, 
        a4stg_rnd_frac_52, a4stg_rnd_frac_51, a4stg_rnd_frac_50, 
        a4stg_rnd_frac_49, a4stg_rnd_frac_48, a4stg_rnd_frac_47, 
        a4stg_rnd_frac_46, a4stg_rnd_frac_45, a4stg_rnd_frac_44, 
        a4stg_rnd_frac_43, a4stg_rnd_frac_42, a4stg_rnd_frac_41, 
        a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac, 
        a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_rnd_frac_9, 
        a4stg_rnd_frac_8, a4stg_rnd_frac_7, a4stg_rnd_frac_6, a4stg_rnd_frac_5, 
        a4stg_rnd_frac_4, a4stg_rnd_frac_3, a4stg_rnd_frac_2, a4stg_rnd_frac_1, 
        a4stg_rnd_frac_pre2[0]}), .en(a6stg_step), .clk(clk), .q(
        a5stg_rnd_frac), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE64_1 i_a5stg_shl ( .din(a4stg_shl), .en(a6stg_step), .clk(clk), .q(
        a5stg_shl), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  INVX0_RVT U3 ( .A(n618), .Y(n617) );
  INVX0_RVT U4 ( .A(a1stg_in2_gt_in1), .Y(n1032) );
  INVX0_RVT U5 ( .A(n1927), .Y(n1923) );
  INVX0_RVT U6 ( .A(n2500), .Y(n2509) );
  INVX0_RVT U7 ( .A(n245), .Y(n246) );
  INVX0_RVT U8 ( .A(n244), .Y(n247) );
  INVX0_RVT U9 ( .A(n281), .Y(n282) );
  INVX0_RVT U10 ( .A(n2256), .Y(n2203) );
  INVX0_RVT U11 ( .A(a4stg_frac_sng_nx), .Y(n1885) );
  INVX0_RVT U12 ( .A(n277), .Y(n283) );
  INVX0_RVT U13 ( .A(n308), .Y(n309) );
  INVX0_RVT U14 ( .A(n2278), .Y(n2259) );
  INVX0_RVT U15 ( .A(n2518), .Y(n800) );
  INVX0_RVT U16 ( .A(n2515), .Y(n789) );
  INVX0_RVT U17 ( .A(n2346), .Y(n2327) );
  INVX0_RVT U18 ( .A(n2475), .Y(n2477) );
  INVX0_RVT U19 ( .A(n307), .Y(n310) );
  INVX0_RVT U20 ( .A(n1251), .Y(n1291) );
  INVX0_RVT U21 ( .A(n346), .Y(n348) );
  INVX0_RVT U22 ( .A(n2220), .Y(n695) );
  INVX0_RVT U23 ( .A(n326), .Y(n328) );
  INVX0_RVT U24 ( .A(n339), .Y(n341) );
  INVX0_RVT U25 ( .A(n2296), .Y(n704) );
  INVX0_RVT U26 ( .A(n334), .Y(n336) );
  INVX0_RVT U27 ( .A(n290), .Y(n284) );
  INVX0_RVT U28 ( .A(n351), .Y(n345) );
  INVX0_RVT U29 ( .A(n321), .Y(n323) );
  INVX0_RVT U30 ( .A(n285), .Y(n287) );
  INVX0_RVT U31 ( .A(n1965), .Y(n1968) );
  INVX0_RVT U32 ( .A(n361), .Y(n363) );
  INVX0_RVT U33 ( .A(n260), .Y(n262) );
  INVX0_RVT U34 ( .A(n255), .Y(n257) );
  INVX0_RVT U35 ( .A(n248), .Y(n250) );
  INVX0_RVT U36 ( .A(n241), .Y(n147) );
  INVX0_RVT U37 ( .A(n356), .Y(n358) );
  INVX0_RVT U38 ( .A(n1294), .Y(n1346) );
  INVX0_RVT U39 ( .A(n272), .Y(n266) );
  INVX0_RVT U40 ( .A(n267), .Y(n269) );
  INVX0_RVT U41 ( .A(n312), .Y(n314) );
  INVX0_RVT U42 ( .A(n302), .Y(n295) );
  INVX0_RVT U43 ( .A(n297), .Y(n299) );
  INVX0_RVT U44 ( .A(n317), .Y(n311) );
  INVX0_RVT U45 ( .A(n2508), .Y(n2488) );
  INVX0_RVT U46 ( .A(n2516), .Y(n817) );
  OR3X1_RVT U47 ( .A1(a4stg_frac_dbl_nx), .A2(n409), .A3(n408), .Y(
        a4stg_frac_38_0_nx) );
  INVX0_RVT U48 ( .A(n1257), .Y(n1260) );
  INVX0_RVT U49 ( .A(n784), .Y(n787) );
  INVX0_RVT U50 ( .A(n1258), .Y(n1259) );
  INVX0_RVT U51 ( .A(n1347), .Y(n1370) );
  INVX0_RVT U52 ( .A(n2490), .Y(n2496) );
  INVX0_RVT U53 ( .A(n1324), .Y(n1325) );
  INVX0_RVT U54 ( .A(n1323), .Y(n1326) );
  INVX0_RVT U55 ( .A(n1297), .Y(n1298) );
  INVX0_RVT U56 ( .A(n1293), .Y(n1299) );
  INVX0_RVT U57 ( .A(n826), .Y(n758) );
  INVX0_RVT U58 ( .A(n366), .Y(n368) );
  INVX0_RVT U59 ( .A(n821), .Y(n822) );
  INVX0_RVT U60 ( .A(n2467), .Y(n2326) );
  OR3X1_RVT U61 ( .A1(n897), .A2(a1stg_norm_sng_in1), .A3(a1stg_norm_dbl_in1), 
        .Y(n1034) );
  INVX0_RVT U62 ( .A(n2456), .Y(n2476) );
  INVX0_RVT U63 ( .A(n1254), .Y(n392) );
  INVX0_RVT U64 ( .A(n1265), .Y(n389) );
  INVX0_RVT U65 ( .A(n1262), .Y(n388) );
  INVX0_RVT U66 ( .A(n676), .Y(n675) );
  INVX0_RVT U67 ( .A(n1382), .Y(n1384) );
  INVX0_RVT U68 ( .A(n1271), .Y(n1273) );
  INVX0_RVT U69 ( .A(n1276), .Y(n1278) );
  INVX0_RVT U70 ( .A(n1377), .Y(n1379) );
  INVX0_RVT U71 ( .A(n1292), .Y(n1307) );
  INVX0_RVT U72 ( .A(n1318), .Y(n1311) );
  INVX0_RVT U73 ( .A(n1313), .Y(n1315) );
  INVX0_RVT U74 ( .A(n1310), .Y(n1319) );
  INVX0_RVT U75 ( .A(n1288), .Y(n1282) );
  INVX0_RVT U76 ( .A(n1283), .Y(n1285) );
  INVX0_RVT U77 ( .A(n1281), .Y(n1289) );
  INVX0_RVT U78 ( .A(n1306), .Y(n1300) );
  INVX0_RVT U79 ( .A(n1301), .Y(n1303) );
  INVX0_RVT U80 ( .A(n1337), .Y(n1339) );
  INVX0_RVT U81 ( .A(n1342), .Y(n1344) );
  INVX0_RVT U82 ( .A(n1350), .Y(n1352) );
  INVX0_RVT U83 ( .A(n1355), .Y(n1357) );
  INVX0_RVT U84 ( .A(n1367), .Y(n1361) );
  INVX0_RVT U85 ( .A(n1362), .Y(n1364) );
  INVX0_RVT U86 ( .A(n1360), .Y(n1368) );
  INVX0_RVT U87 ( .A(n1372), .Y(n1374) );
  INVX0_RVT U88 ( .A(n1333), .Y(n1327) );
  INVX0_RVT U89 ( .A(n1328), .Y(n1330) );
  INVX0_RVT U90 ( .A(n1322), .Y(n1334) );
  INVX0_RVT U91 ( .A(a1stg_in2[52]), .Y(n872) );
  INVX0_RVT U92 ( .A(a1stg_in2[54]), .Y(n870) );
  INVX0_RVT U93 ( .A(a1stg_in1[52]), .Y(n873) );
  INVX0_RVT U94 ( .A(a1stg_in1[54]), .Y(n869) );
  INVX0_RVT U95 ( .A(a2stg_frac2[0]), .Y(n103) );
  INVX0_RVT U96 ( .A(a2stg_shr_cnt_0[0]), .Y(n1957) );
  INVX0_RVT U97 ( .A(a2stg_shr_cnt_0[1]), .Y(n1958) );
  INVX0_RVT U98 ( .A(a4stg_rnd_frac_5), .Y(n400) );
  INVX0_RVT U99 ( .A(a3stg_ld0_frac[5]), .Y(n1206) );
  INVX0_RVT U100 ( .A(a3stg_ld0_frac[4]), .Y(n1207) );
  INVX0_RVT U101 ( .A(a4stg_rnd_frac_4), .Y(n399) );
  INVX0_RVT U102 ( .A(a2stg_shr_cnt_4[3]), .Y(n710) );
  INVX0_RVT U103 ( .A(a2stg_shr_cnt[3]), .Y(n2486) );
  INVX0_RVT U104 ( .A(a2stg_shr_cnt_3[2]), .Y(n2254) );
  INVX0_RVT U105 ( .A(a2stg_frac2a[11]), .Y(n792) );
  INVX0_RVT U106 ( .A(a2stg_frac2a[6]), .Y(n737) );
  INVX0_RVT U107 ( .A(a2stg_frac2a[10]), .Y(n776) );
  INVX0_RVT U108 ( .A(a2stg_frac2a[2]), .Y(n754) );
  INVX0_RVT U109 ( .A(n866), .Y(n411) );
  INVX0_RVT U110 ( .A(a2stg_frac1_in_frac1), .Y(n414) );
  INVX0_RVT U111 ( .A(a2stg_shr_frac2_shr_int), .Y(n1986) );
  INVX0_RVT U112 ( .A(a2stg_sub_step), .Y(n2483) );
  OR3X1_RVT U113 ( .A1(a4stg_rnd_frac_pre1[2]), .A2(a4stg_rnd_frac_pre2[2]), 
        .A3(a4stg_rnd_frac_pre3[2]), .Y(a4stg_rnd_frac_2) );
  OR3X1_RVT U114 ( .A1(a4stg_rnd_frac_pre1[3]), .A2(a4stg_rnd_frac_pre2[3]), 
        .A3(a4stg_rnd_frac_pre3[3]), .Y(a4stg_rnd_frac_3) );
  OR3X1_RVT U115 ( .A1(a4stg_rnd_frac_pre1[9]), .A2(a4stg_rnd_frac_pre2[9]), 
        .A3(a4stg_rnd_frac_pre3[9]), .Y(a4stg_rnd_frac_9) );
  OR3X1_RVT U116 ( .A1(a4stg_rnd_frac_pre1[8]), .A2(a4stg_rnd_frac_pre2[8]), 
        .A3(a4stg_rnd_frac_pre3[8]), .Y(a4stg_rnd_frac_8) );
  OR3X1_RVT U117 ( .A1(a4stg_rnd_frac_pre1[7]), .A2(a4stg_rnd_frac_pre2[7]), 
        .A3(a4stg_rnd_frac_pre3[7]), .Y(a4stg_rnd_frac_7) );
  INVX0_RVT U118 ( .A(a1stg_norm_dbl_in2), .Y(n894) );
  INVX0_RVT U119 ( .A(a1stg_norm_sng_in2), .Y(n895) );
  INVX0_RVT U120 ( .A(a3stg_faddsubopa[0]), .Y(n1211) );
  OA222X1_RVT U121 ( .A1(a4stg_rnd_frac_pre3_in[63]), .A2(n1386), .A3(
        a4stg_rnd_frac_pre3_in[63]), .A4(a3stg_exp10_1_eq0), .A5(
        a4stg_rnd_frac_pre3_in[63]), .A6(a3stg_exp_0), .Y(n1) );
  OR2X1_RVT U122 ( .A1(a2stg_frac1[20]), .A2(n146), .Y(n2) );
  OR2X1_RVT U123 ( .A1(a3stg_frac1[21]), .A2(a3stg_frac2[21]), .Y(n3) );
  OR2X1_RVT U124 ( .A1(a3stg_frac1[20]), .A2(a3stg_frac2[20]), .Y(n4) );
  INVX1_RVT U125 ( .A(a6stg_step), .Y(n2526) );
  AOI22X1_RVT U126 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[46]), .A3(
        a1stg_in2[54]), .A4(a1stg_intlngop), .Y(n6) );
  AOI22X1_RVT U127 ( .A1(n2176), .A2(n1987), .A3(a3stg_frac2[55]), .A4(n2526), 
        .Y(n7) );
  AOI22X1_RVT U128 ( .A1(n2176), .A2(n2148), .A3(a3stg_frac2[37]), .A4(n2526), 
        .Y(n8) );
  AOI22X1_RVT U129 ( .A1(n2176), .A2(n2155), .A3(a3stg_frac2[36]), .A4(n2526), 
        .Y(n9) );
  AOI22X1_RVT U130 ( .A1(n2176), .A2(n2164), .A3(a3stg_frac2[35]), .A4(n2526), 
        .Y(n10) );
  AOI22X1_RVT U131 ( .A1(n2176), .A2(n2172), .A3(a3stg_frac2[34]), .A4(n2526), 
        .Y(n11) );
  AOI22X1_RVT U132 ( .A1(n2176), .A2(n2177), .A3(a3stg_frac2[33]), .A4(n2526), 
        .Y(n12) );
  AOI22X1_RVT U133 ( .A1(n2176), .A2(n2180), .A3(a3stg_frac2[32]), .A4(n2526), 
        .Y(n13) );
  AOI22X1_RVT U134 ( .A1(n2525), .A2(n2421), .A3(a3stg_frac2[6]), .A4(n2526), 
        .Y(n14) );
  AOI22X1_RVT U135 ( .A1(n2525), .A2(n2429), .A3(a3stg_frac2[5]), .A4(n2526), 
        .Y(n15) );
  AOI22X1_RVT U136 ( .A1(n2525), .A2(n2437), .A3(a3stg_frac2[4]), .A4(n2526), 
        .Y(n16) );
  AOI22X1_RVT U137 ( .A1(n2525), .A2(n2445), .A3(a3stg_frac2[3]), .A4(n2526), 
        .Y(n17) );
  AOI22X1_RVT U138 ( .A1(n2525), .A2(n2460), .A3(a3stg_frac2[2]), .A4(n2526), 
        .Y(n18) );
  AOI22X1_RVT U139 ( .A1(n2525), .A2(n2463), .A3(a3stg_frac2[1]), .A4(n2526), 
        .Y(n19) );
  AOI22X1_RVT U140 ( .A1(n2176), .A2(n2049), .A3(a3stg_frac2[48]), .A4(n2526), 
        .Y(n20) );
  AOI22X1_RVT U141 ( .A1(n2176), .A2(n2098), .A3(a3stg_frac2[43]), .A4(n2526), 
        .Y(n21) );
  AOI22X1_RVT U142 ( .A1(n2176), .A2(n2118), .A3(a3stg_frac2[41]), .A4(n2526), 
        .Y(n22) );
  AOI22X1_RVT U143 ( .A1(n2176), .A2(n2127), .A3(a3stg_frac2[40]), .A4(n2526), 
        .Y(n23) );
  AOI22X1_RVT U144 ( .A1(n2176), .A2(n2134), .A3(a3stg_frac2[39]), .A4(n2526), 
        .Y(n24) );
  AOI22X1_RVT U145 ( .A1(n2176), .A2(n2141), .A3(a3stg_frac2[38]), .A4(n2526), 
        .Y(n25) );
  AOI22X1_RVT U146 ( .A1(a1stg_intlngop), .A2(a1stg_in2[61]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[49]), .Y(n26) );
  AOI22X1_RVT U147 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[47]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[46]), .Y(n27) );
  AOI22X1_RVT U148 ( .A1(a1stg_intlngop), .A2(a1stg_in2[60]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[48]), .Y(n28) );
  AOI22X1_RVT U149 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[48]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[47]), .Y(n29) );
  AOI22X1_RVT U150 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[46]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[45]), .Y(n30) );
  AOI22X1_RVT U151 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[44]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[43]), .Y(n31) );
  AOI22X1_RVT U152 ( .A1(a1stg_intlngop), .A2(a1stg_in2[52]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[40]), .Y(n32) );
  INVX1_RVT U153 ( .A(a2stg_frac2_63), .Y(n150) );
  INVX1_RVT U154 ( .A(a2stg_frac2[62]), .Y(n34) );
  AO22X1_RVT U155 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n150), .A3(
        a2stg_fracadd_frac2_inv), .A4(n34), .Y(n33) );
  AO21X1_RVT U156 ( .A1(a2stg_frac2[62]), .A2(a2stg_fracadd_frac2), .A3(n33), 
        .Y(n155) );
  INVX1_RVT U157 ( .A(a2stg_frac2[61]), .Y(n1137) );
  AO22X1_RVT U158 ( .A1(a2stg_fracadd_frac2_inv), .A2(n1137), .A3(
        a2stg_fracadd_frac2_inv_shr1), .A4(n34), .Y(n35) );
  AO21X1_RVT U159 ( .A1(a2stg_frac2[61]), .A2(a2stg_fracadd_frac2), .A3(n35), 
        .Y(n157) );
  INVX1_RVT U160 ( .A(a2stg_frac2[60]), .Y(n1138) );
  AO22X1_RVT U161 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1137), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1138), .Y(n36) );
  AO21X1_RVT U162 ( .A1(a2stg_frac2[60]), .A2(a2stg_fracadd_frac2), .A3(n36), 
        .Y(n159) );
  INVX1_RVT U163 ( .A(a2stg_frac2[59]), .Y(n1139) );
  AO22X1_RVT U164 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1138), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1139), .Y(n37) );
  AO21X1_RVT U165 ( .A1(a2stg_frac2[59]), .A2(a2stg_fracadd_frac2), .A3(n37), 
        .Y(n161) );
  INVX1_RVT U166 ( .A(a2stg_frac2[58]), .Y(n1140) );
  AO22X1_RVT U167 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1139), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1140), .Y(n38) );
  AO21X1_RVT U168 ( .A1(a2stg_frac2[58]), .A2(a2stg_fracadd_frac2), .A3(n38), 
        .Y(n163) );
  INVX1_RVT U169 ( .A(a2stg_frac2[57]), .Y(n1141) );
  AO22X1_RVT U170 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1140), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1141), .Y(n39) );
  AO21X1_RVT U171 ( .A1(a2stg_frac2[57]), .A2(a2stg_fracadd_frac2), .A3(n39), 
        .Y(n165) );
  INVX1_RVT U172 ( .A(a2stg_frac2[56]), .Y(n1142) );
  AO22X1_RVT U173 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1141), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1142), .Y(n40) );
  AO21X1_RVT U174 ( .A1(a2stg_frac2[56]), .A2(a2stg_fracadd_frac2), .A3(n40), 
        .Y(n167) );
  INVX1_RVT U175 ( .A(a2stg_frac2[55]), .Y(n1143) );
  AO22X1_RVT U176 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1142), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1143), .Y(n41) );
  AO21X1_RVT U177 ( .A1(a2stg_frac2[55]), .A2(a2stg_fracadd_frac2), .A3(n41), 
        .Y(n169) );
  INVX1_RVT U178 ( .A(a2stg_frac2[54]), .Y(n1144) );
  AO22X1_RVT U179 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1143), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1144), .Y(n42) );
  AO21X1_RVT U180 ( .A1(a2stg_frac2[54]), .A2(a2stg_fracadd_frac2), .A3(n42), 
        .Y(n171) );
  INVX1_RVT U181 ( .A(a2stg_frac2[53]), .Y(n1129) );
  AO22X1_RVT U182 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1144), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1129), .Y(n43) );
  AO21X1_RVT U183 ( .A1(a2stg_frac2[53]), .A2(a2stg_fracadd_frac2), .A3(n43), 
        .Y(n173) );
  INVX1_RVT U184 ( .A(a2stg_frac2[52]), .Y(n1130) );
  AO22X1_RVT U185 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1129), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1130), .Y(n44) );
  AO21X1_RVT U186 ( .A1(a2stg_frac2[52]), .A2(a2stg_fracadd_frac2), .A3(n44), 
        .Y(n175) );
  INVX1_RVT U187 ( .A(a2stg_frac2[51]), .Y(n1131) );
  AO22X1_RVT U188 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1130), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1131), .Y(n45) );
  AO21X1_RVT U189 ( .A1(a2stg_frac2[51]), .A2(a2stg_fracadd_frac2), .A3(n45), 
        .Y(n177) );
  INVX1_RVT U190 ( .A(a2stg_frac2[50]), .Y(n1132) );
  AO22X1_RVT U191 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1131), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1132), .Y(n46) );
  AO21X1_RVT U192 ( .A1(a2stg_frac2[50]), .A2(a2stg_fracadd_frac2), .A3(n46), 
        .Y(n179) );
  INVX1_RVT U193 ( .A(a2stg_frac2[49]), .Y(n1133) );
  AO22X1_RVT U194 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1132), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1133), .Y(n47) );
  AO21X1_RVT U195 ( .A1(a2stg_frac2[49]), .A2(a2stg_fracadd_frac2), .A3(n47), 
        .Y(n181) );
  INVX1_RVT U196 ( .A(a2stg_frac2[48]), .Y(n1134) );
  AO22X1_RVT U197 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1133), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1134), .Y(n48) );
  AO21X1_RVT U198 ( .A1(a2stg_frac2[48]), .A2(a2stg_fracadd_frac2), .A3(n48), 
        .Y(n183) );
  INVX1_RVT U199 ( .A(a2stg_frac2[47]), .Y(n1135) );
  AO22X1_RVT U200 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1134), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1135), .Y(n49) );
  AO21X1_RVT U201 ( .A1(a2stg_frac2[47]), .A2(a2stg_fracadd_frac2), .A3(n49), 
        .Y(n185) );
  INVX1_RVT U202 ( .A(a2stg_frac2[46]), .Y(n1136) );
  AO22X1_RVT U203 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1135), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1136), .Y(n50) );
  AO21X1_RVT U204 ( .A1(a2stg_frac2[46]), .A2(a2stg_fracadd_frac2), .A3(n50), 
        .Y(n187) );
  INVX1_RVT U205 ( .A(a2stg_frac2[45]), .Y(n1121) );
  AO22X1_RVT U206 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1136), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1121), .Y(n51) );
  AO21X1_RVT U207 ( .A1(a2stg_frac2[45]), .A2(a2stg_fracadd_frac2), .A3(n51), 
        .Y(n189) );
  INVX1_RVT U208 ( .A(a2stg_frac2[44]), .Y(n1122) );
  AO22X1_RVT U209 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1121), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1122), .Y(n52) );
  AO21X1_RVT U210 ( .A1(a2stg_frac2[44]), .A2(a2stg_fracadd_frac2), .A3(n52), 
        .Y(n191) );
  INVX1_RVT U211 ( .A(a2stg_frac2[43]), .Y(n1123) );
  AO22X1_RVT U212 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1122), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1123), .Y(n53) );
  AO21X1_RVT U213 ( .A1(a2stg_frac2[43]), .A2(a2stg_fracadd_frac2), .A3(n53), 
        .Y(n193) );
  INVX1_RVT U214 ( .A(a2stg_frac2[42]), .Y(n1124) );
  AO22X1_RVT U215 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1123), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1124), .Y(n54) );
  AO21X1_RVT U216 ( .A1(a2stg_frac2[42]), .A2(a2stg_fracadd_frac2), .A3(n54), 
        .Y(n195) );
  INVX1_RVT U217 ( .A(a2stg_frac2[41]), .Y(n1125) );
  AO22X1_RVT U218 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1124), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1125), .Y(n55) );
  AO21X1_RVT U219 ( .A1(a2stg_frac2[41]), .A2(a2stg_fracadd_frac2), .A3(n55), 
        .Y(n197) );
  INVX1_RVT U220 ( .A(a2stg_frac2[40]), .Y(n1126) );
  AO22X1_RVT U221 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1125), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1126), .Y(n56) );
  AO21X1_RVT U222 ( .A1(a2stg_frac2[40]), .A2(a2stg_fracadd_frac2), .A3(n56), 
        .Y(n199) );
  INVX1_RVT U223 ( .A(a2stg_frac2[39]), .Y(n1127) );
  AO22X1_RVT U224 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1126), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1127), .Y(n57) );
  AO21X1_RVT U225 ( .A1(a2stg_frac2[39]), .A2(a2stg_fracadd_frac2), .A3(n57), 
        .Y(n201) );
  INVX1_RVT U226 ( .A(a2stg_frac2[38]), .Y(n1128) );
  AO22X1_RVT U227 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1127), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1128), .Y(n58) );
  AO21X1_RVT U228 ( .A1(a2stg_frac2[38]), .A2(a2stg_fracadd_frac2), .A3(n58), 
        .Y(n203) );
  INVX1_RVT U229 ( .A(a2stg_frac2[37]), .Y(n1116) );
  AO22X1_RVT U230 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1128), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1116), .Y(n59) );
  AO21X1_RVT U231 ( .A1(a2stg_frac2[37]), .A2(a2stg_fracadd_frac2), .A3(n59), 
        .Y(n205) );
  INVX1_RVT U232 ( .A(a2stg_frac2[36]), .Y(n1117) );
  AO22X1_RVT U233 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1116), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1117), .Y(n60) );
  AO21X1_RVT U234 ( .A1(a2stg_frac2[36]), .A2(a2stg_fracadd_frac2), .A3(n60), 
        .Y(n207) );
  INVX1_RVT U235 ( .A(a2stg_frac2[35]), .Y(n1118) );
  AO22X1_RVT U236 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1117), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1118), .Y(n61) );
  AO21X1_RVT U237 ( .A1(a2stg_frac2[35]), .A2(a2stg_fracadd_frac2), .A3(n61), 
        .Y(n209) );
  INVX1_RVT U238 ( .A(a2stg_frac2[34]), .Y(n1119) );
  AO22X1_RVT U239 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1118), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1119), .Y(n62) );
  AO21X1_RVT U240 ( .A1(a2stg_frac2[34]), .A2(a2stg_fracadd_frac2), .A3(n62), 
        .Y(n211) );
  INVX1_RVT U241 ( .A(a2stg_frac2[33]), .Y(n64) );
  AO22X1_RVT U242 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1119), .A3(
        a2stg_fracadd_frac2_inv), .A4(n64), .Y(n63) );
  AO21X1_RVT U243 ( .A1(a2stg_frac2[33]), .A2(a2stg_fracadd_frac2), .A3(n63), 
        .Y(n213) );
  INVX1_RVT U244 ( .A(a2stg_frac2[32]), .Y(n66) );
  AO22X1_RVT U245 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n64), .A3(
        a2stg_fracadd_frac2_inv), .A4(n66), .Y(n65) );
  AO21X1_RVT U246 ( .A1(a2stg_frac2[32]), .A2(a2stg_fracadd_frac2), .A3(n65), 
        .Y(n215) );
  INVX1_RVT U247 ( .A(a2stg_frac2[31]), .Y(n1163) );
  AO22X1_RVT U248 ( .A1(a2stg_fracadd_frac2_inv), .A2(n1163), .A3(
        a2stg_fracadd_frac2_inv_shr1), .A4(n66), .Y(n67) );
  AO21X1_RVT U249 ( .A1(a2stg_frac2[31]), .A2(a2stg_fracadd_frac2), .A3(n67), 
        .Y(n217) );
  INVX1_RVT U250 ( .A(a2stg_frac2[30]), .Y(n1164) );
  AO22X1_RVT U251 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1163), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1164), .Y(n68) );
  AO21X1_RVT U252 ( .A1(a2stg_frac2[30]), .A2(a2stg_fracadd_frac2), .A3(n68), 
        .Y(n219) );
  INVX1_RVT U253 ( .A(a2stg_frac2[29]), .Y(n1173) );
  AO22X1_RVT U254 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1164), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1173), .Y(n69) );
  AO21X1_RVT U255 ( .A1(a2stg_frac2[29]), .A2(a2stg_fracadd_frac2), .A3(n69), 
        .Y(n221) );
  INVX1_RVT U256 ( .A(a2stg_frac2[28]), .Y(n1157) );
  AO22X1_RVT U257 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1173), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1157), .Y(n70) );
  AO21X1_RVT U258 ( .A1(a2stg_frac2[28]), .A2(a2stg_fracadd_frac2), .A3(n70), 
        .Y(n223) );
  INVX1_RVT U259 ( .A(a2stg_frac2[27]), .Y(n1158) );
  AO22X1_RVT U260 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1157), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1158), .Y(n71) );
  AO21X1_RVT U261 ( .A1(a2stg_frac2[27]), .A2(a2stg_fracadd_frac2), .A3(n71), 
        .Y(n225) );
  INVX1_RVT U262 ( .A(a2stg_frac2[26]), .Y(n1159) );
  AO22X1_RVT U263 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1158), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1159), .Y(n72) );
  AO21X1_RVT U264 ( .A1(a2stg_frac2[26]), .A2(a2stg_fracadd_frac2), .A3(n72), 
        .Y(n227) );
  INVX1_RVT U265 ( .A(a2stg_frac2[25]), .Y(n1160) );
  AO22X1_RVT U266 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1159), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1160), .Y(n73) );
  AO21X1_RVT U267 ( .A1(a2stg_frac2[25]), .A2(a2stg_fracadd_frac2), .A3(n73), 
        .Y(n229) );
  INVX1_RVT U268 ( .A(a2stg_frac2[24]), .Y(n1153) );
  AO22X1_RVT U269 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1160), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1153), .Y(n74) );
  AO21X1_RVT U270 ( .A1(a2stg_frac2[24]), .A2(a2stg_fracadd_frac2), .A3(n74), 
        .Y(n231) );
  INVX1_RVT U271 ( .A(a2stg_frac2[23]), .Y(n1154) );
  AO22X1_RVT U272 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1153), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1154), .Y(n75) );
  AO21X1_RVT U273 ( .A1(a2stg_frac2[23]), .A2(a2stg_fracadd_frac2), .A3(n75), 
        .Y(n233) );
  INVX1_RVT U274 ( .A(a2stg_frac2[22]), .Y(n1155) );
  AO22X1_RVT U275 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1154), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1155), .Y(n76) );
  AO21X1_RVT U276 ( .A1(a2stg_frac2[22]), .A2(a2stg_fracadd_frac2), .A3(n76), 
        .Y(n235) );
  INVX1_RVT U277 ( .A(a2stg_frac2[21]), .Y(n1156) );
  AO22X1_RVT U278 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1155), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1156), .Y(n77) );
  AO21X1_RVT U279 ( .A1(a2stg_frac2[21]), .A2(a2stg_fracadd_frac2), .A3(n77), 
        .Y(n237) );
  INVX1_RVT U280 ( .A(a2stg_frac2[20]), .Y(n1165) );
  AO22X1_RVT U281 ( .A1(a2stg_fracadd_frac2_inv), .A2(n1165), .A3(
        a2stg_fracadd_frac2_inv_shr1), .A4(n1156), .Y(n78) );
  AO21X1_RVT U282 ( .A1(a2stg_frac2[20]), .A2(a2stg_fracadd_frac2), .A3(n78), 
        .Y(n146) );
  INVX1_RVT U283 ( .A(a2stg_frac2[19]), .Y(n1166) );
  AO22X1_RVT U284 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1165), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1166), .Y(n79) );
  AO21X1_RVT U285 ( .A1(a2stg_frac2[19]), .A2(a2stg_fracadd_frac2), .A3(n79), 
        .Y(n145) );
  NOR2X0_RVT U286 ( .A1(a2stg_frac1[19]), .A2(n145), .Y(n248) );
  INVX1_RVT U287 ( .A(a2stg_frac2[18]), .Y(n1167) );
  AO22X1_RVT U288 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1166), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1167), .Y(n80) );
  AO21X1_RVT U289 ( .A1(a2stg_frac2[18]), .A2(a2stg_fracadd_frac2), .A3(n80), 
        .Y(n142) );
  NOR2X0_RVT U290 ( .A1(a2stg_frac1[18]), .A2(n142), .Y(n255) );
  INVX1_RVT U291 ( .A(a2stg_frac2[17]), .Y(n1168) );
  AO22X1_RVT U292 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1167), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1168), .Y(n81) );
  AO21X1_RVT U293 ( .A1(a2stg_frac2[17]), .A2(a2stg_fracadd_frac2), .A3(n81), 
        .Y(n141) );
  NOR2X0_RVT U294 ( .A1(a2stg_frac1[17]), .A2(n141), .Y(n260) );
  NOR2X0_RVT U295 ( .A1(n255), .A2(n260), .Y(n144) );
  INVX1_RVT U296 ( .A(a2stg_frac2[16]), .Y(n1169) );
  AO22X1_RVT U297 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1168), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1169), .Y(n82) );
  AO21X1_RVT U298 ( .A1(a2stg_frac2[16]), .A2(a2stg_fracadd_frac2), .A3(n82), 
        .Y(n140) );
  NOR2X0_RVT U299 ( .A1(a2stg_frac1[16]), .A2(n140), .Y(n267) );
  INVX1_RVT U300 ( .A(a2stg_frac2[15]), .Y(n1170) );
  AO22X1_RVT U301 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1169), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1170), .Y(n83) );
  AO21X1_RVT U302 ( .A1(a2stg_frac2[15]), .A2(a2stg_fracadd_frac2), .A3(n83), 
        .Y(n139) );
  NOR2X0_RVT U303 ( .A1(a2stg_frac1[15]), .A2(n139), .Y(n265) );
  NOR2X0_RVT U304 ( .A1(n267), .A2(n265), .Y(n254) );
  NAND2X0_RVT U305 ( .A1(n144), .A2(n254), .Y(n244) );
  NOR2X0_RVT U306 ( .A1(n248), .A2(n244), .Y(n240) );
  NAND2X0_RVT U307 ( .A1(n2), .A2(n240), .Y(n149) );
  INVX1_RVT U308 ( .A(a2stg_frac2[14]), .Y(n1171) );
  INVX1_RVT U309 ( .A(a2stg_frac2[13]), .Y(n1172) );
  AO22X1_RVT U310 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1171), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1172), .Y(n84) );
  AO21X1_RVT U311 ( .A1(a2stg_frac2[13]), .A2(a2stg_fracadd_frac2), .A3(n84), 
        .Y(n131) );
  NOR2X0_RVT U312 ( .A1(a2stg_frac1[13]), .A2(n131), .Y(n276) );
  AO22X1_RVT U313 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1170), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1171), .Y(n85) );
  AO21X1_RVT U314 ( .A1(a2stg_frac2[14]), .A2(a2stg_fracadd_frac2), .A3(n85), 
        .Y(n132) );
  NOR2X0_RVT U315 ( .A1(a2stg_frac1[14]), .A2(n132), .Y(n285) );
  NOR2X0_RVT U316 ( .A1(n276), .A2(n285), .Y(n134) );
  INVX1_RVT U317 ( .A(a2stg_frac2[12]), .Y(n1161) );
  AO22X1_RVT U318 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1172), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1161), .Y(n86) );
  AO21X1_RVT U319 ( .A1(a2stg_frac2[12]), .A2(a2stg_fracadd_frac2), .A3(n86), 
        .Y(n130) );
  NOR2X0_RVT U320 ( .A1(a2stg_frac1[12]), .A2(n130), .Y(n297) );
  INVX1_RVT U321 ( .A(a2stg_frac2[11]), .Y(n1162) );
  AO22X1_RVT U322 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n1161), .A3(
        a2stg_fracadd_frac2_inv), .A4(n1162), .Y(n87) );
  AO21X1_RVT U323 ( .A1(a2stg_frac2[11]), .A2(a2stg_fracadd_frac2), .A3(n87), 
        .Y(n129) );
  NOR2X0_RVT U324 ( .A1(a2stg_frac1[11]), .A2(n129), .Y(n294) );
  NOR2X0_RVT U325 ( .A1(n297), .A2(n294), .Y(n277) );
  NAND2X0_RVT U326 ( .A1(n134), .A2(n277), .Y(n136) );
  INVX1_RVT U327 ( .A(a2stg_frac2[8]), .Y(n89) );
  INVX1_RVT U328 ( .A(a2stg_frac2[7]), .Y(n95) );
  AO22X1_RVT U329 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n89), .A3(
        a2stg_fracadd_frac2_inv), .A4(n95), .Y(n88) );
  AO21X1_RVT U330 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[7]), .A3(n88), 
        .Y(n123) );
  NOR2X0_RVT U331 ( .A1(a2stg_frac1[7]), .A2(n123), .Y(n326) );
  INVX1_RVT U332 ( .A(a2stg_frac2[9]), .Y(n91) );
  AO22X1_RVT U333 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n91), .A3(
        a2stg_fracadd_frac2_inv), .A4(n89), .Y(n90) );
  AO21X1_RVT U334 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[8]), .A3(n90), 
        .Y(n124) );
  NOR2X0_RVT U335 ( .A1(a2stg_frac1[8]), .A2(n124), .Y(n321) );
  NOR2X0_RVT U336 ( .A1(n326), .A2(n321), .Y(n307) );
  INVX1_RVT U337 ( .A(a2stg_frac2[10]), .Y(n93) );
  AO22X1_RVT U338 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n93), .A3(
        a2stg_fracadd_frac2_inv), .A4(n91), .Y(n92) );
  AO21X1_RVT U339 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[9]), .A3(n92), 
        .Y(n125) );
  NOR2X0_RVT U340 ( .A1(a2stg_frac1[9]), .A2(n125), .Y(n306) );
  AO22X1_RVT U341 ( .A1(a2stg_fracadd_frac2_inv), .A2(n93), .A3(
        a2stg_fracadd_frac2_inv_shr1), .A4(n1162), .Y(n94) );
  AO21X1_RVT U342 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[10]), .A3(n94), 
        .Y(n126) );
  NOR2X0_RVT U343 ( .A1(a2stg_frac1[10]), .A2(n126), .Y(n312) );
  NOR2X0_RVT U344 ( .A1(n306), .A2(n312), .Y(n128) );
  NAND2X0_RVT U345 ( .A1(n307), .A2(n128), .Y(n280) );
  NOR2X0_RVT U346 ( .A1(n136), .A2(n280), .Y(n138) );
  INVX1_RVT U347 ( .A(a2stg_frac2[6]), .Y(n97) );
  AO22X1_RVT U348 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n95), .A3(
        a2stg_fracadd_frac2_inv), .A4(n97), .Y(n96) );
  AO21X1_RVT U349 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[6]), .A3(n96), 
        .Y(n118) );
  NOR2X0_RVT U350 ( .A1(a2stg_frac1[6]), .A2(n118), .Y(n334) );
  INVX1_RVT U351 ( .A(a2stg_frac2[5]), .Y(n99) );
  AO22X1_RVT U352 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n97), .A3(
        a2stg_fracadd_frac2_inv), .A4(n99), .Y(n98) );
  AO21X1_RVT U353 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[5]), .A3(n98), 
        .Y(n117) );
  NOR2X0_RVT U354 ( .A1(a2stg_frac1[5]), .A2(n117), .Y(n339) );
  NOR2X0_RVT U355 ( .A1(n334), .A2(n339), .Y(n120) );
  INVX1_RVT U356 ( .A(a2stg_frac2[4]), .Y(n101) );
  AO22X1_RVT U357 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n99), .A3(
        a2stg_fracadd_frac2_inv), .A4(n101), .Y(n100) );
  AO21X1_RVT U358 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[4]), .A3(n100), 
        .Y(n116) );
  NOR2X0_RVT U359 ( .A1(a2stg_frac1[4]), .A2(n116), .Y(n346) );
  INVX1_RVT U360 ( .A(a2stg_frac2[3]), .Y(n106) );
  AO22X1_RVT U361 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n101), .A3(
        a2stg_fracadd_frac2_inv), .A4(n106), .Y(n102) );
  AO21X1_RVT U362 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[3]), .A3(n102), 
        .Y(n115) );
  NOR2X0_RVT U363 ( .A1(a2stg_frac1[3]), .A2(n115), .Y(n344) );
  NOR2X0_RVT U364 ( .A1(n346), .A2(n344), .Y(n333) );
  NAND2X0_RVT U365 ( .A1(n120), .A2(n333), .Y(n122) );
  NOR2X0_RVT U366 ( .A1(a2stg_fracadd_cin), .A2(a2stg_frac1[0]), .Y(n366) );
  INVX1_RVT U367 ( .A(a2stg_frac2[1]), .Y(n108) );
  AO22X1_RVT U368 ( .A1(n108), .A2(a2stg_fracadd_frac2_inv_shr1), .A3(n103), 
        .A4(a2stg_fracadd_frac2_inv), .Y(n104) );
  AO21X1_RVT U369 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[0]), .A3(n104), 
        .Y(n370) );
  INVX1_RVT U370 ( .A(n370), .Y(n105) );
  NAND2X0_RVT U371 ( .A1(a2stg_fracadd_cin), .A2(a2stg_frac1[0]), .Y(n367) );
  OAI21X1_RVT U372 ( .A1(n366), .A2(n105), .A3(n367), .Y(n355) );
  INVX1_RVT U373 ( .A(a2stg_frac2[2]), .Y(n109) );
  AO22X1_RVT U374 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n106), .A3(
        a2stg_fracadd_frac2_inv), .A4(n109), .Y(n107) );
  AO21X1_RVT U375 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[2]), .A3(n107), 
        .Y(n112) );
  NOR2X0_RVT U376 ( .A1(a2stg_frac1[2]), .A2(n112), .Y(n356) );
  AO22X1_RVT U377 ( .A1(a2stg_fracadd_frac2_inv_shr1), .A2(n109), .A3(
        a2stg_fracadd_frac2_inv), .A4(n108), .Y(n110) );
  AO21X1_RVT U378 ( .A1(a2stg_fracadd_frac2), .A2(a2stg_frac2[1]), .A3(n110), 
        .Y(n111) );
  NOR2X0_RVT U379 ( .A1(a2stg_frac1[1]), .A2(n111), .Y(n361) );
  NOR2X0_RVT U380 ( .A1(n356), .A2(n361), .Y(n114) );
  NAND2X0_RVT U381 ( .A1(a2stg_frac1[1]), .A2(n111), .Y(n362) );
  NAND2X0_RVT U382 ( .A1(a2stg_frac1[2]), .A2(n112), .Y(n357) );
  OAI21X1_RVT U383 ( .A1(n362), .A2(n356), .A3(n357), .Y(n113) );
  AOI21X1_RVT U384 ( .A1(n355), .A2(n114), .A3(n113), .Y(n331) );
  NAND2X0_RVT U385 ( .A1(a2stg_frac1[3]), .A2(n115), .Y(n351) );
  NAND2X0_RVT U386 ( .A1(a2stg_frac1[4]), .A2(n116), .Y(n347) );
  OAI21X1_RVT U387 ( .A1(n351), .A2(n346), .A3(n347), .Y(n332) );
  NAND2X0_RVT U388 ( .A1(a2stg_frac1[5]), .A2(n117), .Y(n340) );
  NAND2X0_RVT U389 ( .A1(a2stg_frac1[6]), .A2(n118), .Y(n335) );
  OAI21X1_RVT U390 ( .A1(n340), .A2(n334), .A3(n335), .Y(n119) );
  AOI21X1_RVT U391 ( .A1(n120), .A2(n332), .A3(n119), .Y(n121) );
  OAI21X1_RVT U392 ( .A1(n122), .A2(n331), .A3(n121), .Y(n278) );
  NAND2X0_RVT U393 ( .A1(a2stg_frac1[7]), .A2(n123), .Y(n327) );
  NAND2X0_RVT U394 ( .A1(a2stg_frac1[8]), .A2(n124), .Y(n322) );
  OAI21X1_RVT U395 ( .A1(n327), .A2(n321), .A3(n322), .Y(n308) );
  NAND2X0_RVT U396 ( .A1(a2stg_frac1[9]), .A2(n125), .Y(n317) );
  NAND2X0_RVT U397 ( .A1(a2stg_frac1[10]), .A2(n126), .Y(n313) );
  OAI21X1_RVT U398 ( .A1(n317), .A2(n312), .A3(n313), .Y(n127) );
  AOI21X1_RVT U399 ( .A1(n308), .A2(n128), .A3(n127), .Y(n279) );
  NAND2X0_RVT U400 ( .A1(a2stg_frac1[11]), .A2(n129), .Y(n302) );
  NAND2X0_RVT U401 ( .A1(a2stg_frac1[12]), .A2(n130), .Y(n298) );
  OAI21X1_RVT U402 ( .A1(n302), .A2(n297), .A3(n298), .Y(n281) );
  NAND2X0_RVT U403 ( .A1(a2stg_frac1[13]), .A2(n131), .Y(n290) );
  NAND2X0_RVT U404 ( .A1(a2stg_frac1[14]), .A2(n132), .Y(n286) );
  OAI21X1_RVT U405 ( .A1(n290), .A2(n285), .A3(n286), .Y(n133) );
  AOI21X1_RVT U406 ( .A1(n134), .A2(n281), .A3(n133), .Y(n135) );
  OAI21X1_RVT U407 ( .A1(n136), .A2(n279), .A3(n135), .Y(n137) );
  AOI21X1_RVT U408 ( .A1(n138), .A2(n278), .A3(n137), .Y(n238) );
  NAND2X0_RVT U409 ( .A1(a2stg_frac1[15]), .A2(n139), .Y(n272) );
  NAND2X0_RVT U410 ( .A1(a2stg_frac1[16]), .A2(n140), .Y(n268) );
  OAI21X1_RVT U411 ( .A1(n272), .A2(n267), .A3(n268), .Y(n253) );
  NAND2X0_RVT U412 ( .A1(a2stg_frac1[17]), .A2(n141), .Y(n261) );
  NAND2X0_RVT U413 ( .A1(a2stg_frac1[18]), .A2(n142), .Y(n256) );
  OAI21X1_RVT U414 ( .A1(n261), .A2(n255), .A3(n256), .Y(n143) );
  AOI21X1_RVT U415 ( .A1(n144), .A2(n253), .A3(n143), .Y(n245) );
  NAND2X0_RVT U416 ( .A1(a2stg_frac1[19]), .A2(n145), .Y(n249) );
  OAI21X1_RVT U417 ( .A1(n248), .A2(n245), .A3(n249), .Y(n239) );
  NAND2X0_RVT U418 ( .A1(a2stg_frac1[20]), .A2(n146), .Y(n241) );
  AOI21X1_RVT U419 ( .A1(n2), .A2(n239), .A3(n147), .Y(n148) );
  OAI21X1_RVT U420 ( .A1(n149), .A2(n238), .A3(n148), .Y(n236) );
  AO221X1_RVT U421 ( .A1(a2stg_frac2_63), .A2(a2stg_fracadd_frac2), .A3(n150), 
        .A4(a2stg_fracadd_frac2_inv), .A5(a2stg_fracadd_frac2_inv_shr1), .Y(
        n151) );
  XOR2X1_RVT U422 ( .A1(n151), .A2(a2stg_frac1[63]), .Y(n152) );
  XOR2X1_RVT U423 ( .A1(n153), .A2(n152), .Y(a2stg_fracadd[63]) );
  FADDX1_RVT U424 ( .A(a2stg_frac1[62]), .B(n155), .CI(n154), .CO(n153), .S(
        a2stg_fracadd[62]) );
  FADDX1_RVT U425 ( .A(a2stg_frac1[61]), .B(n157), .CI(n156), .CO(n154), .S(
        a2stg_fracadd[61]) );
  FADDX1_RVT U426 ( .A(a2stg_frac1[60]), .B(n159), .CI(n158), .CO(n156), .S(
        a2stg_fracadd[60]) );
  FADDX1_RVT U427 ( .A(a2stg_frac1[59]), .B(n161), .CI(n160), .CO(n158), .S(
        a2stg_fracadd[59]) );
  FADDX1_RVT U428 ( .A(a2stg_frac1[58]), .B(n163), .CI(n162), .CO(n160), .S(
        a2stg_fracadd[58]) );
  FADDX1_RVT U429 ( .A(a2stg_frac1[57]), .B(n165), .CI(n164), .CO(n162), .S(
        a2stg_fracadd[57]) );
  FADDX1_RVT U430 ( .A(a2stg_frac1[56]), .B(n167), .CI(n166), .CO(n164), .S(
        a2stg_fracadd[56]) );
  FADDX1_RVT U431 ( .A(a2stg_frac1[55]), .B(n169), .CI(n168), .CO(n166), .S(
        a2stg_fracadd[55]) );
  FADDX1_RVT U432 ( .A(a2stg_frac1[54]), .B(n171), .CI(n170), .CO(n168), .S(
        a2stg_fracadd[54]) );
  FADDX1_RVT U433 ( .A(a2stg_frac1[53]), .B(n173), .CI(n172), .CO(n170), .S(
        a2stg_fracadd[53]) );
  FADDX1_RVT U434 ( .A(a2stg_frac1[52]), .B(n175), .CI(n174), .CO(n172), .S(
        a2stg_fracadd[52]) );
  FADDX1_RVT U435 ( .A(a2stg_frac1[51]), .B(n177), .CI(n176), .CO(n174), .S(
        a2stg_fracadd[51]) );
  FADDX1_RVT U436 ( .A(a2stg_frac1[50]), .B(n179), .CI(n178), .CO(n176), .S(
        a2stg_fracadd[50]) );
  FADDX1_RVT U437 ( .A(a2stg_frac1[49]), .B(n181), .CI(n180), .CO(n178), .S(
        a2stg_fracadd[49]) );
  FADDX1_RVT U438 ( .A(a2stg_frac1[48]), .B(n183), .CI(n182), .CO(n180), .S(
        a2stg_fracadd[48]) );
  FADDX1_RVT U439 ( .A(a2stg_frac1[47]), .B(n185), .CI(n184), .CO(n182), .S(
        a2stg_fracadd[47]) );
  FADDX1_RVT U440 ( .A(a2stg_frac1[46]), .B(n187), .CI(n186), .CO(n184), .S(
        a2stg_fracadd[46]) );
  FADDX1_RVT U441 ( .A(a2stg_frac1[45]), .B(n189), .CI(n188), .CO(n186), .S(
        a2stg_fracadd[45]) );
  FADDX1_RVT U442 ( .A(a2stg_frac1[44]), .B(n191), .CI(n190), .CO(n188), .S(
        a2stg_fracadd[44]) );
  FADDX1_RVT U443 ( .A(a2stg_frac1[43]), .B(n193), .CI(n192), .CO(n190), .S(
        a2stg_fracadd[43]) );
  FADDX1_RVT U444 ( .A(a2stg_frac1[42]), .B(n195), .CI(n194), .CO(n192), .S(
        a2stg_fracadd[42]) );
  FADDX1_RVT U445 ( .A(a2stg_frac1[41]), .B(n197), .CI(n196), .CO(n194), .S(
        a2stg_fracadd[41]) );
  FADDX1_RVT U446 ( .A(a2stg_frac1[40]), .B(n199), .CI(n198), .CO(n196), .S(
        a2stg_fracadd[40]) );
  FADDX1_RVT U447 ( .A(a2stg_frac1[39]), .B(n201), .CI(n200), .CO(n198), .S(
        a2stg_fracadd[39]) );
  FADDX1_RVT U448 ( .A(a2stg_frac1[38]), .B(n203), .CI(n202), .CO(n200), .S(
        a2stg_fracadd[38]) );
  FADDX1_RVT U449 ( .A(a2stg_frac1[37]), .B(n205), .CI(n204), .CO(n202), .S(
        a2stg_fracadd[37]) );
  FADDX1_RVT U450 ( .A(a2stg_frac1[36]), .B(n207), .CI(n206), .CO(n204), .S(
        a2stg_fracadd[36]) );
  FADDX1_RVT U451 ( .A(a2stg_frac1[35]), .B(n209), .CI(n208), .CO(n206), .S(
        a2stg_fracadd[35]) );
  FADDX1_RVT U452 ( .A(a2stg_frac1[34]), .B(n211), .CI(n210), .CO(n208), .S(
        a2stg_fracadd[34]) );
  FADDX1_RVT U453 ( .A(a2stg_frac1[33]), .B(n213), .CI(n212), .CO(n210), .S(
        a2stg_fracadd[33]) );
  FADDX1_RVT U454 ( .A(a2stg_frac1[32]), .B(n215), .CI(n214), .CO(n212), .S(
        a2stg_fracadd[32]) );
  FADDX1_RVT U455 ( .A(a2stg_frac1[31]), .B(n217), .CI(n216), .CO(n214), .S(
        a2stg_fracadd[31]) );
  FADDX1_RVT U456 ( .A(a2stg_frac1[30]), .B(n219), .CI(n218), .CO(n216), .S(
        a2stg_fracadd[30]) );
  FADDX1_RVT U457 ( .A(a2stg_frac1[29]), .B(n221), .CI(n220), .CO(n218), .S(
        a2stg_fracadd[29]) );
  FADDX1_RVT U458 ( .A(a2stg_frac1[28]), .B(n223), .CI(n222), .CO(n220), .S(
        a2stg_fracadd[28]) );
  FADDX1_RVT U459 ( .A(a2stg_frac1[27]), .B(n225), .CI(n224), .CO(n222), .S(
        a2stg_fracadd[27]) );
  FADDX1_RVT U460 ( .A(a2stg_frac1[26]), .B(n227), .CI(n226), .CO(n224), .S(
        a2stg_fracadd[26]) );
  FADDX1_RVT U461 ( .A(a2stg_frac1[25]), .B(n229), .CI(n228), .CO(n226), .S(
        a2stg_fracadd[25]) );
  FADDX1_RVT U462 ( .A(a2stg_frac1[24]), .B(n231), .CI(n230), .CO(n228), .S(
        a2stg_fracadd[24]) );
  FADDX1_RVT U463 ( .A(a2stg_frac1[23]), .B(n233), .CI(n232), .CO(n230), .S(
        a2stg_fracadd[23]) );
  FADDX1_RVT U464 ( .A(a2stg_frac1[22]), .B(n235), .CI(n234), .CO(n232), .S(
        a2stg_fracadd[22]) );
  FADDX1_RVT U465 ( .A(a2stg_frac1[21]), .B(n237), .CI(n236), .CO(n234), .S(
        a2stg_fracadd[21]) );
  INVX1_RVT U466 ( .A(n238), .Y(n275) );
  AOI21X1_RVT U467 ( .A1(n240), .A2(n275), .A3(n239), .Y(n243) );
  NAND2X0_RVT U468 ( .A1(n2), .A2(n241), .Y(n242) );
  XOR2X1_RVT U469 ( .A1(n243), .A2(n242), .Y(a2stg_fracadd[20]) );
  AOI21X1_RVT U470 ( .A1(n247), .A2(n275), .A3(n246), .Y(n252) );
  NAND2X0_RVT U471 ( .A1(n250), .A2(n249), .Y(n251) );
  XOR2X1_RVT U472 ( .A1(n252), .A2(n251), .Y(a2stg_fracadd[19]) );
  AOI21X1_RVT U473 ( .A1(n254), .A2(n275), .A3(n253), .Y(n264) );
  OAI21X1_RVT U474 ( .A1(n260), .A2(n264), .A3(n261), .Y(n259) );
  NAND2X0_RVT U475 ( .A1(n257), .A2(n256), .Y(n258) );
  XNOR2X1_RVT U476 ( .A1(n259), .A2(n258), .Y(a2stg_fracadd[18]) );
  NAND2X0_RVT U477 ( .A1(n262), .A2(n261), .Y(n263) );
  XOR2X1_RVT U478 ( .A1(n264), .A2(n263), .Y(a2stg_fracadd[17]) );
  INVX1_RVT U479 ( .A(n265), .Y(n273) );
  AOI21X1_RVT U480 ( .A1(n273), .A2(n275), .A3(n266), .Y(n271) );
  NAND2X0_RVT U481 ( .A1(n269), .A2(n268), .Y(n270) );
  XOR2X1_RVT U482 ( .A1(n271), .A2(n270), .Y(a2stg_fracadd[16]) );
  NAND2X0_RVT U483 ( .A1(n273), .A2(n272), .Y(n274) );
  XNOR2X1_RVT U484 ( .A1(n275), .A2(n274), .Y(a2stg_fracadd[15]) );
  INVX1_RVT U485 ( .A(n276), .Y(n291) );
  INVX1_RVT U486 ( .A(n278), .Y(n330) );
  OAI21X1_RVT U487 ( .A1(n280), .A2(n330), .A3(n279), .Y(n296) );
  INVX1_RVT U488 ( .A(n296), .Y(n305) );
  OAI21X1_RVT U489 ( .A1(n283), .A2(n305), .A3(n282), .Y(n293) );
  AOI21X1_RVT U490 ( .A1(n291), .A2(n293), .A3(n284), .Y(n289) );
  NAND2X0_RVT U491 ( .A1(n287), .A2(n286), .Y(n288) );
  XOR2X1_RVT U492 ( .A1(n289), .A2(n288), .Y(a2stg_fracadd[14]) );
  NAND2X0_RVT U493 ( .A1(n291), .A2(n290), .Y(n292) );
  XNOR2X1_RVT U494 ( .A1(n293), .A2(n292), .Y(a2stg_fracadd[13]) );
  INVX1_RVT U495 ( .A(n294), .Y(n303) );
  AOI21X1_RVT U496 ( .A1(n303), .A2(n296), .A3(n295), .Y(n301) );
  NAND2X0_RVT U497 ( .A1(n299), .A2(n298), .Y(n300) );
  XOR2X1_RVT U498 ( .A1(n301), .A2(n300), .Y(a2stg_fracadd[12]) );
  NAND2X0_RVT U499 ( .A1(n303), .A2(n302), .Y(n304) );
  XOR2X1_RVT U500 ( .A1(n305), .A2(n304), .Y(a2stg_fracadd[11]) );
  INVX1_RVT U501 ( .A(n306), .Y(n318) );
  OAI21X1_RVT U502 ( .A1(n310), .A2(n330), .A3(n309), .Y(n320) );
  AOI21X1_RVT U503 ( .A1(n318), .A2(n320), .A3(n311), .Y(n316) );
  NAND2X0_RVT U504 ( .A1(n314), .A2(n313), .Y(n315) );
  XOR2X1_RVT U505 ( .A1(n316), .A2(n315), .Y(a2stg_fracadd[10]) );
  NAND2X0_RVT U506 ( .A1(n318), .A2(n317), .Y(n319) );
  XNOR2X1_RVT U507 ( .A1(n320), .A2(n319), .Y(a2stg_fracadd[9]) );
  OAI21X1_RVT U508 ( .A1(n326), .A2(n330), .A3(n327), .Y(n325) );
  NAND2X0_RVT U509 ( .A1(n323), .A2(n322), .Y(n324) );
  XNOR2X1_RVT U510 ( .A1(n325), .A2(n324), .Y(a2stg_fracadd[8]) );
  NAND2X0_RVT U511 ( .A1(n328), .A2(n327), .Y(n329) );
  XOR2X1_RVT U512 ( .A1(n330), .A2(n329), .Y(a2stg_fracadd[7]) );
  INVX1_RVT U513 ( .A(n331), .Y(n354) );
  AOI21X1_RVT U514 ( .A1(n333), .A2(n354), .A3(n332), .Y(n343) );
  OAI21X1_RVT U515 ( .A1(n339), .A2(n343), .A3(n340), .Y(n338) );
  NAND2X0_RVT U516 ( .A1(n336), .A2(n335), .Y(n337) );
  XNOR2X1_RVT U517 ( .A1(n338), .A2(n337), .Y(a2stg_fracadd[6]) );
  NAND2X0_RVT U518 ( .A1(n341), .A2(n340), .Y(n342) );
  XOR2X1_RVT U519 ( .A1(n343), .A2(n342), .Y(a2stg_fracadd[5]) );
  INVX1_RVT U520 ( .A(n344), .Y(n352) );
  AOI21X1_RVT U521 ( .A1(n352), .A2(n354), .A3(n345), .Y(n350) );
  NAND2X0_RVT U522 ( .A1(n348), .A2(n347), .Y(n349) );
  XOR2X1_RVT U523 ( .A1(n350), .A2(n349), .Y(a2stg_fracadd[4]) );
  NAND2X0_RVT U524 ( .A1(n352), .A2(n351), .Y(n353) );
  XNOR2X1_RVT U525 ( .A1(n354), .A2(n353), .Y(a2stg_fracadd[3]) );
  INVX1_RVT U526 ( .A(n355), .Y(n364) );
  OAI21X1_RVT U527 ( .A1(n361), .A2(n364), .A3(n362), .Y(n360) );
  NAND2X0_RVT U528 ( .A1(n358), .A2(n357), .Y(n359) );
  XNOR2X1_RVT U529 ( .A1(n360), .A2(n359), .Y(a2stg_fracadd[2]) );
  NAND2X0_RVT U530 ( .A1(n363), .A2(n362), .Y(n365) );
  XOR2X1_RVT U531 ( .A1(n365), .A2(n364), .Y(a2stg_fracadd[1]) );
  NAND2X0_RVT U532 ( .A1(n368), .A2(n367), .Y(n369) );
  XNOR2X1_RVT U533 ( .A1(n370), .A2(n369), .Y(a2stg_fracadd[0]) );
  INVX1_RVT U534 ( .A(a4stg_shl_cnt[1]), .Y(n1813) );
  INVX1_RVT U535 ( .A(se), .Y(n2543) );
  AND2X1_RVT U536 ( .A1(n1546), .A2(n1826), .Y(n1874) );
  AND2X1_RVT U537 ( .A1(a4stg_shl_data[0]), .A2(a4stg_shl_cnt_dec54_0[2]), .Y(
        n1819) );
  INVX1_RVT U538 ( .A(a4stg_shl_cnt[0]), .Y(n1800) );
  OA221X1_RVT U539 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[2]), .A3(n1800), 
        .A4(a4stg_shl_data[1]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1794) );
  OA222X1_RVT U540 ( .A1(n1813), .A2(n1819), .A3(n1813), .A4(n1800), .A5(
        a4stg_shl_cnt[1]), .A6(n1794), .Y(n1832) );
  AND2X1_RVT U541 ( .A1(n1874), .A2(n1832), .Y(a4stg_shl[2]) );
  NOR2X0_RVT U542 ( .A1(a3stg_frac1[19]), .A2(a3stg_frac2[19]), .Y(n1261) );
  INVX1_RVT U543 ( .A(n1261), .Y(n1266) );
  NAND2X0_RVT U544 ( .A1(n4), .A2(n1266), .Y(n391) );
  NOR2X0_RVT U545 ( .A1(a3stg_frac1[18]), .A2(a3stg_frac2[18]), .Y(n1271) );
  NOR2X0_RVT U546 ( .A1(a3stg_frac1[17]), .A2(a3stg_frac2[17]), .Y(n1276) );
  NOR2X0_RVT U547 ( .A1(n1271), .A2(n1276), .Y(n387) );
  NOR2X0_RVT U548 ( .A1(a3stg_frac1[16]), .A2(a3stg_frac2[16]), .Y(n1283) );
  NOR2X0_RVT U549 ( .A1(a3stg_frac1[15]), .A2(a3stg_frac2[15]), .Y(n1281) );
  NOR2X0_RVT U550 ( .A1(n1283), .A2(n1281), .Y(n1270) );
  NAND2X0_RVT U551 ( .A1(n387), .A2(n1270), .Y(n1257) );
  NOR2X0_RVT U552 ( .A1(n391), .A2(n1257), .Y(n1253) );
  NAND2X0_RVT U553 ( .A1(n3), .A2(n1253), .Y(n394) );
  NOR2X0_RVT U554 ( .A1(a3stg_frac1[14]), .A2(a3stg_frac2[14]), .Y(n1301) );
  NOR2X0_RVT U555 ( .A1(a3stg_frac1[13]), .A2(a3stg_frac2[13]), .Y(n1292) );
  NOR2X0_RVT U556 ( .A1(n1301), .A2(n1292), .Y(n381) );
  NOR2X0_RVT U557 ( .A1(a3stg_frac1[12]), .A2(a3stg_frac2[12]), .Y(n1313) );
  NOR2X0_RVT U558 ( .A1(a3stg_frac1[11]), .A2(a3stg_frac2[11]), .Y(n1310) );
  NOR2X0_RVT U559 ( .A1(n1313), .A2(n1310), .Y(n1293) );
  NAND2X0_RVT U560 ( .A1(n381), .A2(n1293), .Y(n383) );
  NOR2X0_RVT U561 ( .A1(a3stg_frac1[10]), .A2(a3stg_frac2[10]), .Y(n1328) );
  NOR2X0_RVT U562 ( .A1(a3stg_frac1[9]), .A2(a3stg_frac2[9]), .Y(n1322) );
  NOR2X0_RVT U563 ( .A1(n1328), .A2(n1322), .Y(n379) );
  NOR2X0_RVT U564 ( .A1(a3stg_frac1[8]), .A2(a3stg_frac2[8]), .Y(n1337) );
  NOR2X0_RVT U565 ( .A1(a3stg_frac1[7]), .A2(a3stg_frac2[7]), .Y(n1342) );
  NOR2X0_RVT U566 ( .A1(n1337), .A2(n1342), .Y(n1323) );
  NAND2X0_RVT U567 ( .A1(n379), .A2(n1323), .Y(n1296) );
  NOR2X0_RVT U568 ( .A1(n383), .A2(n1296), .Y(n385) );
  NOR2X0_RVT U569 ( .A1(a3stg_frac1[6]), .A2(a3stg_frac2[6]), .Y(n1350) );
  NOR2X0_RVT U570 ( .A1(a3stg_frac1[5]), .A2(a3stg_frac2[5]), .Y(n1355) );
  NOR2X0_RVT U571 ( .A1(n1350), .A2(n1355), .Y(n375) );
  NOR2X0_RVT U572 ( .A1(a3stg_frac1[4]), .A2(a3stg_frac2[4]), .Y(n1362) );
  NOR2X0_RVT U573 ( .A1(a3stg_frac1[3]), .A2(a3stg_frac2[3]), .Y(n1360) );
  NOR2X0_RVT U574 ( .A1(n1362), .A2(n1360), .Y(n1349) );
  NAND2X0_RVT U575 ( .A1(n375), .A2(n1349), .Y(n377) );
  NOR2X0_RVT U576 ( .A1(a3stg_frac1[2]), .A2(a3stg_frac2[2]), .Y(n1372) );
  NOR2X0_RVT U577 ( .A1(a3stg_frac1[1]), .A2(a3stg_frac2[1]), .Y(n1377) );
  NOR2X0_RVT U578 ( .A1(n1372), .A2(n1377), .Y(n373) );
  INVX1_RVT U579 ( .A(a3stg_frac2[0]), .Y(n371) );
  NOR2X0_RVT U580 ( .A1(a3stg_suba), .A2(a3stg_frac1[0]), .Y(n1382) );
  NAND2X0_RVT U581 ( .A1(a3stg_suba), .A2(a3stg_frac1[0]), .Y(n1383) );
  OAI21X1_RVT U582 ( .A1(n371), .A2(n1382), .A3(n1383), .Y(n1371) );
  NAND2X0_RVT U583 ( .A1(a3stg_frac1[1]), .A2(a3stg_frac2[1]), .Y(n1378) );
  NAND2X0_RVT U584 ( .A1(a3stg_frac1[2]), .A2(a3stg_frac2[2]), .Y(n1373) );
  OAI21X1_RVT U585 ( .A1(n1378), .A2(n1372), .A3(n1373), .Y(n372) );
  AOI21X1_RVT U586 ( .A1(n373), .A2(n1371), .A3(n372), .Y(n1347) );
  NAND2X0_RVT U587 ( .A1(a3stg_frac1[3]), .A2(a3stg_frac2[3]), .Y(n1367) );
  NAND2X0_RVT U588 ( .A1(a3stg_frac1[4]), .A2(a3stg_frac2[4]), .Y(n1363) );
  OAI21X1_RVT U589 ( .A1(n1367), .A2(n1362), .A3(n1363), .Y(n1348) );
  NAND2X0_RVT U590 ( .A1(a3stg_frac1[5]), .A2(a3stg_frac2[5]), .Y(n1356) );
  NAND2X0_RVT U591 ( .A1(a3stg_frac1[6]), .A2(a3stg_frac2[6]), .Y(n1351) );
  OAI21X1_RVT U592 ( .A1(n1356), .A2(n1350), .A3(n1351), .Y(n374) );
  AOI21X1_RVT U593 ( .A1(n375), .A2(n1348), .A3(n374), .Y(n376) );
  OAI21X1_RVT U594 ( .A1(n377), .A2(n1347), .A3(n376), .Y(n1294) );
  NAND2X0_RVT U595 ( .A1(a3stg_frac1[7]), .A2(a3stg_frac2[7]), .Y(n1343) );
  NAND2X0_RVT U596 ( .A1(a3stg_frac1[8]), .A2(a3stg_frac2[8]), .Y(n1338) );
  OAI21X1_RVT U597 ( .A1(n1343), .A2(n1337), .A3(n1338), .Y(n1324) );
  NAND2X0_RVT U598 ( .A1(a3stg_frac1[9]), .A2(a3stg_frac2[9]), .Y(n1333) );
  NAND2X0_RVT U599 ( .A1(a3stg_frac1[10]), .A2(a3stg_frac2[10]), .Y(n1329) );
  OAI21X1_RVT U600 ( .A1(n1333), .A2(n1328), .A3(n1329), .Y(n378) );
  AOI21X1_RVT U601 ( .A1(n379), .A2(n1324), .A3(n378), .Y(n1295) );
  NAND2X0_RVT U602 ( .A1(a3stg_frac1[11]), .A2(a3stg_frac2[11]), .Y(n1318) );
  NAND2X0_RVT U603 ( .A1(a3stg_frac1[12]), .A2(a3stg_frac2[12]), .Y(n1314) );
  OAI21X1_RVT U604 ( .A1(n1318), .A2(n1313), .A3(n1314), .Y(n1297) );
  NAND2X0_RVT U605 ( .A1(a3stg_frac1[13]), .A2(a3stg_frac2[13]), .Y(n1306) );
  NAND2X0_RVT U606 ( .A1(a3stg_frac1[14]), .A2(a3stg_frac2[14]), .Y(n1302) );
  OAI21X1_RVT U607 ( .A1(n1306), .A2(n1301), .A3(n1302), .Y(n380) );
  AOI21X1_RVT U608 ( .A1(n381), .A2(n1297), .A3(n380), .Y(n382) );
  OAI21X1_RVT U609 ( .A1(n383), .A2(n1295), .A3(n382), .Y(n384) );
  AOI21X1_RVT U610 ( .A1(n385), .A2(n1294), .A3(n384), .Y(n1251) );
  NAND2X0_RVT U611 ( .A1(a3stg_frac1[15]), .A2(a3stg_frac2[15]), .Y(n1288) );
  NAND2X0_RVT U612 ( .A1(a3stg_frac1[16]), .A2(a3stg_frac2[16]), .Y(n1284) );
  OAI21X1_RVT U613 ( .A1(n1288), .A2(n1283), .A3(n1284), .Y(n1269) );
  NAND2X0_RVT U614 ( .A1(a3stg_frac1[17]), .A2(a3stg_frac2[17]), .Y(n1277) );
  NAND2X0_RVT U615 ( .A1(a3stg_frac1[18]), .A2(a3stg_frac2[18]), .Y(n1272) );
  OAI21X1_RVT U616 ( .A1(n1277), .A2(n1271), .A3(n1272), .Y(n386) );
  AOI21X1_RVT U617 ( .A1(n387), .A2(n1269), .A3(n386), .Y(n1258) );
  NAND2X0_RVT U618 ( .A1(a3stg_frac1[19]), .A2(a3stg_frac2[19]), .Y(n1265) );
  NAND2X0_RVT U619 ( .A1(a3stg_frac1[20]), .A2(a3stg_frac2[20]), .Y(n1262) );
  AOI21X1_RVT U620 ( .A1(n389), .A2(n4), .A3(n388), .Y(n390) );
  OAI21X1_RVT U621 ( .A1(n391), .A2(n1258), .A3(n390), .Y(n1252) );
  NAND2X0_RVT U622 ( .A1(a3stg_frac1[21]), .A2(a3stg_frac2[21]), .Y(n1254) );
  AOI21X1_RVT U623 ( .A1(n3), .A2(n1252), .A3(n392), .Y(n393) );
  OAI21X1_RVT U624 ( .A1(n394), .A2(n1251), .A3(n393), .Y(n1250) );
  XOR2X1_RVT U625 ( .A1(n395), .A2(\DP_OP_16J2_123_4718/n1 ), .Y(n1920) );
  INVX1_RVT U626 ( .A(n1920), .Y(a3stg_inc_exp_inv) );
  INVX1_RVT U627 ( .A(a3stg_exp10_0_eq0), .Y(n1921) );
  FADDX1_RVT U628 ( .A(a3stg_frac1[62]), .B(a3stg_frac2[62]), .CI(n396), .CO(
        n395), .S(n1404) );
  NAND2X0_RVT U629 ( .A1(a6stg_step), .A2(a3stg_faddsubopa[1]), .Y(n866) );
  AND4X1_RVT U630 ( .A1(a3stg_inc_exp_inv), .A2(n1921), .A3(n1404), .A4(n411), 
        .Y(a4stg_rnd_frac_pre3_in[63]) );
  OR3X2_RVT U631 ( .A1(a4stg_rnd_frac_pre1[39]), .A2(a4stg_rnd_frac_pre2[39]), 
        .A3(a4stg_rnd_frac_pre3[39]), .Y(a4stg_rnd_frac_39) );
  OR3X2_RVT U632 ( .A1(a4stg_rnd_frac_pre1[10]), .A2(a4stg_rnd_frac_pre2[10]), 
        .A3(a4stg_rnd_frac_pre3[10]), .Y(a4stg_rnd_frac_10) );
  OR3X2_RVT U633 ( .A1(a4stg_rnd_frac_pre1[5]), .A2(a4stg_rnd_frac_pre2[5]), 
        .A3(a4stg_rnd_frac_pre3[5]), .Y(a4stg_rnd_frac_5) );
  OR3X2_RVT U634 ( .A1(a4stg_rnd_frac_pre1[4]), .A2(a4stg_rnd_frac_pre2[4]), 
        .A3(a4stg_rnd_frac_pre3[4]), .Y(a4stg_rnd_frac_4) );
  OR2X1_RVT U635 ( .A1(a4stg_rnd_frac_pre2[1]), .A2(a4stg_rnd_frac_pre3[1]), 
        .Y(a4stg_rnd_frac_1) );
  NOR4X1_RVT U636 ( .A1(a4stg_rnd_frac_pre2[0]), .A2(a4stg_rnd_frac_2), .A3(
        a4stg_rnd_frac_3), .A4(a4stg_rnd_frac_1), .Y(n398) );
  OR3X2_RVT U637 ( .A1(a4stg_rnd_frac_pre1[6]), .A2(a4stg_rnd_frac_pre2[6]), 
        .A3(a4stg_rnd_frac_pre3[6]), .Y(a4stg_rnd_frac_6) );
  NOR4X1_RVT U638 ( .A1(a4stg_rnd_frac_9), .A2(a4stg_rnd_frac_8), .A3(
        a4stg_rnd_frac_7), .A4(a4stg_rnd_frac_6), .Y(n397) );
  NAND4X0_RVT U639 ( .A1(n400), .A2(n399), .A3(n398), .A4(n397), .Y(
        a4stg_frac_9_0_nx) );
  OR2X1_RVT U640 ( .A1(a4stg_rnd_frac_10), .A2(a4stg_frac_9_0_nx), .Y(
        a4stg_frac_dbl_nx) );
  OR3X2_RVT U641 ( .A1(a4stg_rnd_frac_pre1[14]), .A2(a4stg_rnd_frac_pre2[14]), 
        .A3(a4stg_rnd_frac_pre3[14]), .Y(a4stg_rnd_frac[14]) );
  OR3X2_RVT U642 ( .A1(a4stg_rnd_frac_pre1[13]), .A2(a4stg_rnd_frac_pre2[13]), 
        .A3(a4stg_rnd_frac_pre3[13]), .Y(a4stg_rnd_frac[13]) );
  OR3X2_RVT U643 ( .A1(a4stg_rnd_frac_pre1[12]), .A2(a4stg_rnd_frac_pre2[12]), 
        .A3(a4stg_rnd_frac_pre3[12]), .Y(a4stg_rnd_frac[12]) );
  OR3X2_RVT U644 ( .A1(a4stg_rnd_frac_pre1[11]), .A2(a4stg_rnd_frac_pre2[11]), 
        .A3(a4stg_rnd_frac_pre3[11]), .Y(a4stg_rnd_frac_11) );
  NOR4X1_RVT U645 ( .A1(a4stg_rnd_frac[14]), .A2(a4stg_rnd_frac[13]), .A3(
        a4stg_rnd_frac[12]), .A4(a4stg_rnd_frac_11), .Y(n403) );
  OR3X2_RVT U646 ( .A1(a4stg_rnd_frac_pre1[19]), .A2(a4stg_rnd_frac_pre2[19]), 
        .A3(a4stg_rnd_frac_pre3[19]), .Y(a4stg_rnd_frac[19]) );
  OR3X2_RVT U647 ( .A1(a4stg_rnd_frac_pre1[17]), .A2(a4stg_rnd_frac_pre2[17]), 
        .A3(a4stg_rnd_frac_pre3[17]), .Y(a4stg_rnd_frac[17]) );
  OR3X2_RVT U648 ( .A1(a4stg_rnd_frac_pre1[16]), .A2(a4stg_rnd_frac_pre2[16]), 
        .A3(a4stg_rnd_frac_pre3[16]), .Y(a4stg_rnd_frac[16]) );
  OR3X2_RVT U649 ( .A1(a4stg_rnd_frac_pre1[15]), .A2(a4stg_rnd_frac_pre2[15]), 
        .A3(a4stg_rnd_frac_pre3[15]), .Y(a4stg_rnd_frac[15]) );
  NOR4X1_RVT U650 ( .A1(a4stg_rnd_frac[19]), .A2(a4stg_rnd_frac[17]), .A3(
        a4stg_rnd_frac[16]), .A4(a4stg_rnd_frac[15]), .Y(n402) );
  OR3X2_RVT U651 ( .A1(a4stg_rnd_frac_pre1[38]), .A2(a4stg_rnd_frac_pre2[38]), 
        .A3(a4stg_rnd_frac_pre3[38]), .Y(a4stg_rnd_frac[38]) );
  OR3X2_RVT U652 ( .A1(a4stg_rnd_frac_pre1[37]), .A2(a4stg_rnd_frac_pre2[37]), 
        .A3(a4stg_rnd_frac_pre3[37]), .Y(a4stg_rnd_frac[37]) );
  OR3X2_RVT U653 ( .A1(a4stg_rnd_frac_pre1[36]), .A2(a4stg_rnd_frac_pre2[36]), 
        .A3(a4stg_rnd_frac_pre3[36]), .Y(a4stg_rnd_frac[36]) );
  OR3X2_RVT U654 ( .A1(a4stg_rnd_frac_pre1[34]), .A2(a4stg_rnd_frac_pre2[34]), 
        .A3(a4stg_rnd_frac_pre3[34]), .Y(a4stg_rnd_frac[34]) );
  NOR4X1_RVT U655 ( .A1(a4stg_rnd_frac[38]), .A2(a4stg_rnd_frac[37]), .A3(
        a4stg_rnd_frac[36]), .A4(a4stg_rnd_frac[34]), .Y(n401) );
  NAND3X0_RVT U656 ( .A1(n403), .A2(n402), .A3(n401), .Y(n409) );
  OR3X2_RVT U657 ( .A1(a4stg_rnd_frac_pre1[26]), .A2(a4stg_rnd_frac_pre2[26]), 
        .A3(a4stg_rnd_frac_pre3[26]), .Y(a4stg_rnd_frac[26]) );
  OR3X2_RVT U658 ( .A1(a4stg_rnd_frac_pre1[25]), .A2(a4stg_rnd_frac_pre2[25]), 
        .A3(a4stg_rnd_frac_pre3[25]), .Y(a4stg_rnd_frac[25]) );
  OR3X2_RVT U659 ( .A1(a4stg_rnd_frac_pre1[24]), .A2(a4stg_rnd_frac_pre2[24]), 
        .A3(a4stg_rnd_frac_pre3[24]), .Y(a4stg_rnd_frac[24]) );
  OR3X2_RVT U660 ( .A1(a4stg_rnd_frac_pre1[23]), .A2(a4stg_rnd_frac_pre2[23]), 
        .A3(a4stg_rnd_frac_pre3[23]), .Y(a4stg_rnd_frac[23]) );
  NOR4X1_RVT U661 ( .A1(a4stg_rnd_frac[26]), .A2(a4stg_rnd_frac[25]), .A3(
        a4stg_rnd_frac[24]), .A4(a4stg_rnd_frac[23]), .Y(n407) );
  OR3X2_RVT U662 ( .A1(a4stg_rnd_frac_pre1[22]), .A2(a4stg_rnd_frac_pre2[22]), 
        .A3(a4stg_rnd_frac_pre3[22]), .Y(a4stg_rnd_frac[22]) );
  OR3X2_RVT U663 ( .A1(a4stg_rnd_frac_pre1[21]), .A2(a4stg_rnd_frac_pre2[21]), 
        .A3(a4stg_rnd_frac_pre3[21]), .Y(a4stg_rnd_frac[21]) );
  OR3X2_RVT U664 ( .A1(a4stg_rnd_frac_pre1[20]), .A2(a4stg_rnd_frac_pre2[20]), 
        .A3(a4stg_rnd_frac_pre3[20]), .Y(a4stg_rnd_frac[20]) );
  OR3X2_RVT U665 ( .A1(a4stg_rnd_frac_pre1[18]), .A2(a4stg_rnd_frac_pre2[18]), 
        .A3(a4stg_rnd_frac_pre3[18]), .Y(a4stg_rnd_frac[18]) );
  NOR4X1_RVT U666 ( .A1(a4stg_rnd_frac[22]), .A2(a4stg_rnd_frac[21]), .A3(
        a4stg_rnd_frac[20]), .A4(a4stg_rnd_frac[18]), .Y(n406) );
  OR3X2_RVT U667 ( .A1(a4stg_rnd_frac_pre1[35]), .A2(a4stg_rnd_frac_pre2[35]), 
        .A3(a4stg_rnd_frac_pre3[35]), .Y(a4stg_rnd_frac[35]) );
  OR3X2_RVT U668 ( .A1(a4stg_rnd_frac_pre1[33]), .A2(a4stg_rnd_frac_pre2[33]), 
        .A3(a4stg_rnd_frac_pre3[33]), .Y(a4stg_rnd_frac[33]) );
  OR3X2_RVT U669 ( .A1(a4stg_rnd_frac_pre1[32]), .A2(a4stg_rnd_frac_pre2[32]), 
        .A3(a4stg_rnd_frac_pre3[32]), .Y(a4stg_rnd_frac[32]) );
  OR3X2_RVT U670 ( .A1(a4stg_rnd_frac_pre1[30]), .A2(a4stg_rnd_frac_pre2[30]), 
        .A3(a4stg_rnd_frac_pre3[30]), .Y(a4stg_rnd_frac[30]) );
  NOR4X1_RVT U671 ( .A1(a4stg_rnd_frac[35]), .A2(a4stg_rnd_frac[33]), .A3(
        a4stg_rnd_frac[32]), .A4(a4stg_rnd_frac[30]), .Y(n405) );
  OR3X2_RVT U672 ( .A1(a4stg_rnd_frac_pre1[31]), .A2(a4stg_rnd_frac_pre2[31]), 
        .A3(a4stg_rnd_frac_pre3[31]), .Y(a4stg_rnd_frac[31]) );
  OR3X2_RVT U673 ( .A1(a4stg_rnd_frac_pre1[29]), .A2(a4stg_rnd_frac_pre2[29]), 
        .A3(a4stg_rnd_frac_pre3[29]), .Y(a4stg_rnd_frac[29]) );
  OR3X2_RVT U674 ( .A1(a4stg_rnd_frac_pre1[28]), .A2(a4stg_rnd_frac_pre2[28]), 
        .A3(a4stg_rnd_frac_pre3[28]), .Y(a4stg_rnd_frac[28]) );
  OR3X2_RVT U675 ( .A1(a4stg_rnd_frac_pre1[27]), .A2(a4stg_rnd_frac_pre2[27]), 
        .A3(a4stg_rnd_frac_pre3[27]), .Y(a4stg_rnd_frac[27]) );
  NOR4X1_RVT U676 ( .A1(a4stg_rnd_frac[31]), .A2(a4stg_rnd_frac[29]), .A3(
        a4stg_rnd_frac[28]), .A4(a4stg_rnd_frac[27]), .Y(n404) );
  NAND4X0_RVT U677 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .Y(n408) );
  OR2X1_RVT U678 ( .A1(a4stg_rnd_frac_39), .A2(a4stg_frac_38_0_nx), .Y(
        a4stg_frac_sng_nx) );
  OR3X2_RVT U679 ( .A1(a4stg_rnd_frac_pre1[40]), .A2(a4stg_rnd_frac_pre2[40]), 
        .A3(a4stg_rnd_frac_pre3[40]), .Y(a4stg_rnd_frac_40) );
  NAND4X0_RVT U680 ( .A1(a4stg_rnd_dbl), .A2(a4stg_rnd_frac[13]), .A3(
        a4stg_rnd_frac[12]), .A4(a4stg_rnd_frac_11), .Y(n674) );
  INVX1_RVT U681 ( .A(n674), .Y(n673) );
  NAND2X0_RVT U682 ( .A1(n673), .A2(a4stg_rnd_frac[14]), .Y(n672) );
  INVX1_RVT U683 ( .A(n672), .Y(n671) );
  NAND2X0_RVT U684 ( .A1(n671), .A2(a4stg_rnd_frac[15]), .Y(n670) );
  INVX1_RVT U685 ( .A(n670), .Y(n669) );
  NAND2X0_RVT U686 ( .A1(n669), .A2(a4stg_rnd_frac[16]), .Y(n668) );
  INVX1_RVT U687 ( .A(n668), .Y(n667) );
  NAND2X0_RVT U688 ( .A1(n667), .A2(a4stg_rnd_frac[17]), .Y(n666) );
  INVX1_RVT U689 ( .A(n666), .Y(n665) );
  NAND2X0_RVT U690 ( .A1(n665), .A2(a4stg_rnd_frac[18]), .Y(n664) );
  INVX1_RVT U691 ( .A(n664), .Y(n663) );
  NAND2X0_RVT U692 ( .A1(n663), .A2(a4stg_rnd_frac[19]), .Y(n662) );
  INVX1_RVT U693 ( .A(n662), .Y(n661) );
  NAND2X0_RVT U694 ( .A1(n661), .A2(a4stg_rnd_frac[20]), .Y(n660) );
  INVX1_RVT U695 ( .A(n660), .Y(n659) );
  NAND2X0_RVT U696 ( .A1(n659), .A2(a4stg_rnd_frac[21]), .Y(n658) );
  INVX1_RVT U697 ( .A(n658), .Y(n657) );
  NAND2X0_RVT U698 ( .A1(n657), .A2(a4stg_rnd_frac[22]), .Y(n656) );
  INVX1_RVT U699 ( .A(n656), .Y(n655) );
  NAND2X0_RVT U700 ( .A1(n655), .A2(a4stg_rnd_frac[23]), .Y(n654) );
  INVX1_RVT U701 ( .A(n654), .Y(n653) );
  NAND2X0_RVT U702 ( .A1(n653), .A2(a4stg_rnd_frac[24]), .Y(n652) );
  INVX1_RVT U703 ( .A(n652), .Y(n651) );
  NAND2X0_RVT U704 ( .A1(n651), .A2(a4stg_rnd_frac[25]), .Y(n650) );
  INVX1_RVT U705 ( .A(n650), .Y(n649) );
  NAND2X0_RVT U706 ( .A1(n649), .A2(a4stg_rnd_frac[26]), .Y(n648) );
  INVX1_RVT U707 ( .A(n648), .Y(n647) );
  NAND2X0_RVT U708 ( .A1(n647), .A2(a4stg_rnd_frac[27]), .Y(n646) );
  INVX1_RVT U709 ( .A(n646), .Y(n645) );
  NAND2X0_RVT U710 ( .A1(n645), .A2(a4stg_rnd_frac[28]), .Y(n644) );
  INVX1_RVT U711 ( .A(n644), .Y(n643) );
  NAND2X0_RVT U712 ( .A1(n643), .A2(a4stg_rnd_frac[29]), .Y(n642) );
  INVX1_RVT U713 ( .A(n642), .Y(n641) );
  NAND2X0_RVT U714 ( .A1(n641), .A2(a4stg_rnd_frac[30]), .Y(n640) );
  INVX1_RVT U715 ( .A(n640), .Y(n639) );
  NAND2X0_RVT U716 ( .A1(n639), .A2(a4stg_rnd_frac[31]), .Y(n638) );
  INVX1_RVT U717 ( .A(n638), .Y(n637) );
  NAND2X0_RVT U718 ( .A1(n637), .A2(a4stg_rnd_frac[32]), .Y(n636) );
  INVX1_RVT U719 ( .A(n636), .Y(n635) );
  NAND2X0_RVT U720 ( .A1(n635), .A2(a4stg_rnd_frac[33]), .Y(n634) );
  INVX1_RVT U721 ( .A(n634), .Y(n633) );
  NAND2X0_RVT U722 ( .A1(n633), .A2(a4stg_rnd_frac[34]), .Y(n632) );
  INVX1_RVT U723 ( .A(n632), .Y(n631) );
  NAND2X0_RVT U724 ( .A1(n631), .A2(a4stg_rnd_frac[35]), .Y(n630) );
  INVX1_RVT U725 ( .A(n630), .Y(n629) );
  NAND2X0_RVT U726 ( .A1(n629), .A2(a4stg_rnd_frac[36]), .Y(n628) );
  INVX1_RVT U727 ( .A(n628), .Y(n627) );
  NAND2X0_RVT U728 ( .A1(n627), .A2(a4stg_rnd_frac[37]), .Y(n626) );
  INVX1_RVT U729 ( .A(n626), .Y(n625) );
  NAND2X0_RVT U730 ( .A1(n625), .A2(a4stg_rnd_frac[38]), .Y(n624) );
  INVX1_RVT U731 ( .A(n624), .Y(n623) );
  NAND2X0_RVT U732 ( .A1(n623), .A2(a4stg_rnd_frac_39), .Y(n622) );
  INVX1_RVT U733 ( .A(n622), .Y(n621) );
  OR3X2_RVT U734 ( .A1(a4stg_rnd_frac_pre1[43]), .A2(a4stg_rnd_frac_pre2[43]), 
        .A3(a4stg_rnd_frac_pre3[43]), .Y(a4stg_rnd_frac_43) );
  OR3X2_RVT U735 ( .A1(a4stg_rnd_frac_pre1[42]), .A2(a4stg_rnd_frac_pre2[42]), 
        .A3(a4stg_rnd_frac_pre3[42]), .Y(a4stg_rnd_frac_42) );
  OR3X2_RVT U736 ( .A1(a4stg_rnd_frac_pre1[41]), .A2(a4stg_rnd_frac_pre2[41]), 
        .A3(a4stg_rnd_frac_pre3[41]), .Y(a4stg_rnd_frac_41) );
  NAND4X0_RVT U737 ( .A1(n620), .A2(a4stg_rnd_frac_43), .A3(a4stg_rnd_frac_42), 
        .A4(a4stg_rnd_frac_41), .Y(n616) );
  INVX1_RVT U738 ( .A(n616), .Y(n615) );
  OR3X2_RVT U739 ( .A1(a4stg_rnd_frac_pre1[44]), .A2(a4stg_rnd_frac_pre2[44]), 
        .A3(a4stg_rnd_frac_pre3[44]), .Y(a4stg_rnd_frac_44) );
  NAND2X0_RVT U740 ( .A1(n615), .A2(a4stg_rnd_frac_44), .Y(n614) );
  INVX1_RVT U741 ( .A(n614), .Y(n613) );
  OR3X2_RVT U742 ( .A1(a4stg_rnd_frac_pre1[45]), .A2(a4stg_rnd_frac_pre2[45]), 
        .A3(a4stg_rnd_frac_pre3[45]), .Y(a4stg_rnd_frac_45) );
  NAND2X0_RVT U743 ( .A1(n613), .A2(a4stg_rnd_frac_45), .Y(n612) );
  INVX1_RVT U744 ( .A(n612), .Y(n611) );
  OR3X2_RVT U745 ( .A1(a4stg_rnd_frac_pre1[46]), .A2(a4stg_rnd_frac_pre2[46]), 
        .A3(a4stg_rnd_frac_pre3[46]), .Y(a4stg_rnd_frac_46) );
  NAND2X0_RVT U746 ( .A1(n611), .A2(a4stg_rnd_frac_46), .Y(n610) );
  INVX1_RVT U747 ( .A(n610), .Y(n609) );
  OR3X2_RVT U748 ( .A1(a4stg_rnd_frac_pre1[47]), .A2(a4stg_rnd_frac_pre2[47]), 
        .A3(a4stg_rnd_frac_pre3[47]), .Y(a4stg_rnd_frac_47) );
  NAND2X0_RVT U749 ( .A1(n609), .A2(a4stg_rnd_frac_47), .Y(n608) );
  INVX1_RVT U750 ( .A(n608), .Y(n607) );
  OR3X2_RVT U751 ( .A1(a4stg_rnd_frac_pre1[48]), .A2(a4stg_rnd_frac_pre2[48]), 
        .A3(a4stg_rnd_frac_pre3[48]), .Y(a4stg_rnd_frac_48) );
  NAND2X0_RVT U752 ( .A1(n607), .A2(a4stg_rnd_frac_48), .Y(n606) );
  INVX1_RVT U753 ( .A(n606), .Y(n605) );
  OR3X2_RVT U754 ( .A1(a4stg_rnd_frac_pre1[49]), .A2(a4stg_rnd_frac_pre2[49]), 
        .A3(a4stg_rnd_frac_pre3[49]), .Y(a4stg_rnd_frac_49) );
  NAND2X0_RVT U755 ( .A1(n605), .A2(a4stg_rnd_frac_49), .Y(n604) );
  INVX1_RVT U756 ( .A(n604), .Y(n603) );
  OR3X2_RVT U757 ( .A1(a4stg_rnd_frac_pre1[50]), .A2(a4stg_rnd_frac_pre2[50]), 
        .A3(a4stg_rnd_frac_pre3[50]), .Y(a4stg_rnd_frac_50) );
  NAND2X0_RVT U758 ( .A1(n603), .A2(a4stg_rnd_frac_50), .Y(n602) );
  INVX1_RVT U759 ( .A(n602), .Y(n601) );
  OR3X2_RVT U760 ( .A1(a4stg_rnd_frac_pre1[51]), .A2(a4stg_rnd_frac_pre2[51]), 
        .A3(a4stg_rnd_frac_pre3[51]), .Y(a4stg_rnd_frac_51) );
  NAND2X0_RVT U761 ( .A1(n601), .A2(a4stg_rnd_frac_51), .Y(n600) );
  INVX1_RVT U762 ( .A(n600), .Y(n599) );
  OR3X2_RVT U763 ( .A1(a4stg_rnd_frac_pre1[52]), .A2(a4stg_rnd_frac_pre2[52]), 
        .A3(a4stg_rnd_frac_pre3[52]), .Y(a4stg_rnd_frac_52) );
  NAND2X0_RVT U764 ( .A1(n599), .A2(a4stg_rnd_frac_52), .Y(n598) );
  INVX1_RVT U765 ( .A(n598), .Y(n597) );
  OR3X2_RVT U766 ( .A1(a4stg_rnd_frac_pre1[53]), .A2(a4stg_rnd_frac_pre2[53]), 
        .A3(a4stg_rnd_frac_pre3[53]), .Y(a4stg_rnd_frac_53) );
  NAND2X0_RVT U767 ( .A1(n597), .A2(a4stg_rnd_frac_53), .Y(n596) );
  INVX1_RVT U768 ( .A(n596), .Y(n595) );
  OR3X2_RVT U769 ( .A1(a4stg_rnd_frac_pre1[54]), .A2(a4stg_rnd_frac_pre2[54]), 
        .A3(a4stg_rnd_frac_pre3[54]), .Y(a4stg_rnd_frac_54) );
  NAND2X0_RVT U770 ( .A1(n595), .A2(a4stg_rnd_frac_54), .Y(n594) );
  INVX1_RVT U771 ( .A(n594), .Y(n593) );
  OR3X2_RVT U772 ( .A1(a4stg_rnd_frac_pre1[55]), .A2(a4stg_rnd_frac_pre2[55]), 
        .A3(a4stg_rnd_frac_pre3[55]), .Y(a4stg_rnd_frac_55) );
  NAND2X0_RVT U773 ( .A1(n593), .A2(a4stg_rnd_frac_55), .Y(n592) );
  INVX1_RVT U774 ( .A(n592), .Y(n591) );
  OR3X2_RVT U775 ( .A1(a4stg_rnd_frac_pre1[56]), .A2(a4stg_rnd_frac_pre2[56]), 
        .A3(a4stg_rnd_frac_pre3[56]), .Y(a4stg_rnd_frac_56) );
  NAND2X0_RVT U776 ( .A1(n591), .A2(a4stg_rnd_frac_56), .Y(n590) );
  INVX1_RVT U777 ( .A(n590), .Y(n589) );
  OR3X2_RVT U778 ( .A1(a4stg_rnd_frac_pre1[57]), .A2(a4stg_rnd_frac_pre2[57]), 
        .A3(a4stg_rnd_frac_pre3[57]), .Y(a4stg_rnd_frac_57) );
  NAND2X0_RVT U779 ( .A1(n589), .A2(a4stg_rnd_frac_57), .Y(n588) );
  INVX1_RVT U780 ( .A(n588), .Y(n587) );
  OR3X2_RVT U781 ( .A1(a4stg_rnd_frac_pre1[58]), .A2(a4stg_rnd_frac_pre2[58]), 
        .A3(a4stg_rnd_frac_pre3[58]), .Y(a4stg_rnd_frac_58) );
  NAND2X0_RVT U782 ( .A1(n587), .A2(a4stg_rnd_frac_58), .Y(n586) );
  INVX1_RVT U783 ( .A(n586), .Y(n585) );
  OR3X2_RVT U784 ( .A1(a4stg_rnd_frac_pre1[59]), .A2(a4stg_rnd_frac_pre2[59]), 
        .A3(a4stg_rnd_frac_pre3[59]), .Y(a4stg_rnd_frac_59) );
  NAND2X0_RVT U785 ( .A1(n585), .A2(a4stg_rnd_frac_59), .Y(n584) );
  INVX1_RVT U786 ( .A(n584), .Y(n583) );
  OR3X2_RVT U787 ( .A1(a4stg_rnd_frac_pre1[60]), .A2(a4stg_rnd_frac_pre2[60]), 
        .A3(a4stg_rnd_frac_pre3[60]), .Y(a4stg_rnd_frac_60) );
  NAND2X0_RVT U788 ( .A1(n583), .A2(a4stg_rnd_frac_60), .Y(n582) );
  INVX1_RVT U789 ( .A(n582), .Y(n581) );
  OR3X2_RVT U790 ( .A1(a4stg_rnd_frac_pre1[61]), .A2(a4stg_rnd_frac_pre2[61]), 
        .A3(a4stg_rnd_frac_pre3[61]), .Y(a4stg_rnd_frac_61) );
  NAND2X0_RVT U791 ( .A1(n581), .A2(a4stg_rnd_frac_61), .Y(n580) );
  INVX1_RVT U792 ( .A(n580), .Y(n579) );
  OR3X2_RVT U793 ( .A1(a4stg_rnd_frac_pre1[62]), .A2(a4stg_rnd_frac_pre2[62]), 
        .A3(a4stg_rnd_frac_pre3[62]), .Y(a4stg_rnd_frac_62) );
  NAND2X0_RVT U794 ( .A1(n579), .A2(a4stg_rnd_frac_62), .Y(n578) );
  INVX1_RVT U795 ( .A(n578), .Y(a4stg_rndadd_cout) );
  FADDX1_RVT U796 ( .A(a3stg_frac1[61]), .B(a3stg_frac2[61]), .CI(n410), .CO(
        n396), .S(n1919) );
  OR3X2_RVT U797 ( .A1(n1404), .A2(n1920), .A3(n1919), .Y(a4stg_round_in) );
  OR3X2_RVT U798 ( .A1(a4stg_rnd_frac_pre1[63]), .A2(a4stg_rnd_frac_pre2[63]), 
        .A3(a4stg_rnd_frac_pre3[63]), .Y(a4stg_rnd_frac_63) );
  INVX1_RVT U799 ( .A(n1404), .Y(n1922) );
  AND4X1_RVT U800 ( .A1(n411), .A2(n1919), .A3(n1922), .A4(a3stg_inc_exp_inv), 
        .Y(n1386) );
  INVX1_RVT U801 ( .A(a3stg_exp10_1_eq0), .Y(n412) );
  AND2X1_RVT U802 ( .A1(n1386), .A2(n412), .Y(n2542) );
  NAND2X0_RVT U811 ( .A1(a1stg_in2_gt_in1), .A2(a1stg_2nan_in_inv), .Y(n413)
         );
  AO21X1_RVT U812 ( .A1(n414), .A2(n413), .A3(a1stg_faddsubop_inv), .Y(n1024)
         );
  AND2X1_RVT U813 ( .A1(a1stg_norm_dbl_in1), .A2(n1024), .Y(n1027) );
  AND2X1_RVT U814 ( .A1(a1stg_denorm_dbl_in1), .A2(n1024), .Y(n470) );
  AOI22X1_RVT U815 ( .A1(n1027), .A2(a1stg_in1[1]), .A3(n470), .A4(
        a1stg_in1[0]), .Y(n417) );
  OR2X1_RVT U816 ( .A1(a2stg_frac1_in_frac2), .A2(n1024), .Y(n907) );
  AND2X1_RVT U817 ( .A1(a2stg_frac1_in_nv_dbl), .A2(n907), .Y(n1029) );
  INVX1_RVT U818 ( .A(n1029), .Y(n416) );
  OA21X1_RVT U819 ( .A1(a1stg_in2_gt_in1), .A2(a2stg_frac1_in_frac1), .A3(
        a2stg_frac1_in_frac2), .Y(n1030) );
  AO222X1_RVT U820 ( .A1(a1stg_intlngop), .A2(a1stg_in2[12]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[0]), .A5(a1stg_in2[1]), .A6(
        a1stg_norm_dbl_in2), .Y(n1111) );
  NAND2X0_RVT U821 ( .A1(n1030), .A2(n1111), .Y(n415) );
  NAND3X0_RVT U822 ( .A1(n417), .A2(n416), .A3(n415), .Y(a2stg_frac1_in[12])
         );
  AOI22X1_RVT U823 ( .A1(n1027), .A2(a1stg_in1[2]), .A3(n470), .A4(
        a1stg_in1[1]), .Y(n419) );
  AO222X1_RVT U824 ( .A1(a1stg_intlngop), .A2(a1stg_in2[13]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[1]), .A5(a1stg_in2[2]), .A6(
        a1stg_norm_dbl_in2), .Y(n1109) );
  NAND2X0_RVT U825 ( .A1(n1030), .A2(n1109), .Y(n418) );
  NAND3X0_RVT U826 ( .A1(n419), .A2(n416), .A3(n418), .Y(a2stg_frac1_in[13])
         );
  AOI22X1_RVT U827 ( .A1(n1027), .A2(a1stg_in1[3]), .A3(n470), .A4(
        a1stg_in1[2]), .Y(n421) );
  AO222X1_RVT U828 ( .A1(a1stg_intlngop), .A2(a1stg_in2[14]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[2]), .A5(a1stg_in2[3]), .A6(
        a1stg_norm_dbl_in2), .Y(n1108) );
  NAND2X0_RVT U829 ( .A1(n1030), .A2(n1108), .Y(n420) );
  NAND3X0_RVT U830 ( .A1(n421), .A2(n416), .A3(n420), .Y(a2stg_frac1_in[14])
         );
  AOI22X1_RVT U831 ( .A1(n1027), .A2(a1stg_in1[4]), .A3(n470), .A4(
        a1stg_in1[3]), .Y(n423) );
  AO222X1_RVT U832 ( .A1(a1stg_intlngop), .A2(a1stg_in2[15]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[3]), .A5(a1stg_in2[4]), .A6(
        a1stg_norm_dbl_in2), .Y(n1107) );
  NAND2X0_RVT U833 ( .A1(n1030), .A2(n1107), .Y(n422) );
  NAND3X0_RVT U834 ( .A1(n423), .A2(n416), .A3(n422), .Y(a2stg_frac1_in[15])
         );
  AOI22X1_RVT U835 ( .A1(n1027), .A2(a1stg_in1[5]), .A3(n470), .A4(
        a1stg_in1[4]), .Y(n425) );
  AO222X1_RVT U836 ( .A1(a1stg_intlngop), .A2(a1stg_in2[16]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[4]), .A5(a1stg_in2[5]), .A6(
        a1stg_norm_dbl_in2), .Y(n1106) );
  NAND2X0_RVT U837 ( .A1(n1030), .A2(n1106), .Y(n424) );
  NAND3X0_RVT U838 ( .A1(n425), .A2(n416), .A3(n424), .Y(a2stg_frac1_in[16])
         );
  AOI22X1_RVT U839 ( .A1(n1027), .A2(a1stg_in1[6]), .A3(n470), .A4(
        a1stg_in1[5]), .Y(n427) );
  AO222X1_RVT U840 ( .A1(a1stg_intlngop), .A2(a1stg_in2[17]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[5]), .A5(a1stg_in2[6]), .A6(
        a1stg_norm_dbl_in2), .Y(n1105) );
  NAND2X0_RVT U841 ( .A1(n1030), .A2(n1105), .Y(n426) );
  NAND3X0_RVT U842 ( .A1(n427), .A2(n416), .A3(n426), .Y(a2stg_frac1_in[17])
         );
  AOI22X1_RVT U843 ( .A1(n1027), .A2(a1stg_in1[7]), .A3(n470), .A4(
        a1stg_in1[6]), .Y(n429) );
  AO222X1_RVT U844 ( .A1(a1stg_intlngop), .A2(a1stg_in2[18]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[6]), .A5(a1stg_in2[7]), .A6(
        a1stg_norm_dbl_in2), .Y(n1104) );
  NAND2X0_RVT U845 ( .A1(n1030), .A2(n1104), .Y(n428) );
  NAND3X0_RVT U846 ( .A1(n429), .A2(n416), .A3(n428), .Y(a2stg_frac1_in[18])
         );
  AOI22X1_RVT U847 ( .A1(n1027), .A2(a1stg_in1[8]), .A3(n470), .A4(
        a1stg_in1[7]), .Y(n431) );
  AO222X1_RVT U848 ( .A1(a1stg_intlngop), .A2(a1stg_in2[19]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[7]), .A5(a1stg_in2[8]), .A6(
        a1stg_norm_dbl_in2), .Y(n1103) );
  NAND2X0_RVT U849 ( .A1(n1030), .A2(n1103), .Y(n430) );
  NAND3X0_RVT U850 ( .A1(n431), .A2(n416), .A3(n430), .Y(a2stg_frac1_in[19])
         );
  AOI22X1_RVT U851 ( .A1(n1027), .A2(a1stg_in1[9]), .A3(n470), .A4(
        a1stg_in1[8]), .Y(n433) );
  AO222X1_RVT U852 ( .A1(a1stg_intlngop), .A2(a1stg_in2[20]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[8]), .A5(a1stg_in2[9]), .A6(
        a1stg_norm_dbl_in2), .Y(n1102) );
  NAND2X0_RVT U853 ( .A1(n1030), .A2(n1102), .Y(n432) );
  NAND3X0_RVT U854 ( .A1(n433), .A2(n416), .A3(n432), .Y(a2stg_frac1_in[20])
         );
  AOI22X1_RVT U855 ( .A1(n1027), .A2(a1stg_in1[10]), .A3(n470), .A4(
        a1stg_in1[9]), .Y(n435) );
  AO222X1_RVT U856 ( .A1(a1stg_intlngop), .A2(a1stg_in2[21]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[9]), .A5(a1stg_in2[10]), .A6(
        a1stg_norm_dbl_in2), .Y(n1101) );
  NAND2X0_RVT U857 ( .A1(n1030), .A2(n1101), .Y(n434) );
  NAND3X0_RVT U858 ( .A1(n435), .A2(n416), .A3(n434), .Y(a2stg_frac1_in[21])
         );
  AOI22X1_RVT U859 ( .A1(n1027), .A2(a1stg_in1[11]), .A3(n470), .A4(
        a1stg_in1[10]), .Y(n437) );
  AO222X1_RVT U860 ( .A1(a1stg_intlngop), .A2(a1stg_in2[22]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[10]), .A5(a1stg_in2[11]), .A6(
        a1stg_norm_dbl_in2), .Y(n1100) );
  NAND2X0_RVT U861 ( .A1(n1030), .A2(n1100), .Y(n436) );
  NAND3X0_RVT U862 ( .A1(n437), .A2(n416), .A3(n436), .Y(a2stg_frac1_in[22])
         );
  AOI22X1_RVT U863 ( .A1(n1027), .A2(a1stg_in1[12]), .A3(n470), .A4(
        a1stg_in1[11]), .Y(n439) );
  AO222X1_RVT U864 ( .A1(a1stg_intlngop), .A2(a1stg_in2[23]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[11]), .A5(a1stg_in2[12]), .A6(
        a1stg_norm_dbl_in2), .Y(n1099) );
  NAND2X0_RVT U865 ( .A1(n1030), .A2(n1099), .Y(n438) );
  NAND3X0_RVT U866 ( .A1(n439), .A2(n416), .A3(n438), .Y(a2stg_frac1_in[23])
         );
  AOI22X1_RVT U867 ( .A1(n1027), .A2(a1stg_in1[13]), .A3(n470), .A4(
        a1stg_in1[12]), .Y(n441) );
  AO222X1_RVT U868 ( .A1(a1stg_intlngop), .A2(a1stg_in2[24]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[12]), .A5(a1stg_in2[13]), .A6(
        a1stg_norm_dbl_in2), .Y(n1098) );
  NAND2X0_RVT U869 ( .A1(n1030), .A2(n1098), .Y(n440) );
  NAND3X0_RVT U870 ( .A1(n441), .A2(n416), .A3(n440), .Y(a2stg_frac1_in[24])
         );
  AOI22X1_RVT U871 ( .A1(n1027), .A2(a1stg_in1[14]), .A3(n470), .A4(
        a1stg_in1[13]), .Y(n443) );
  AO222X1_RVT U872 ( .A1(a1stg_intlngop), .A2(a1stg_in2[25]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[13]), .A5(a1stg_in2[14]), .A6(
        a1stg_norm_dbl_in2), .Y(n1097) );
  NAND2X0_RVT U873 ( .A1(n1030), .A2(n1097), .Y(n442) );
  NAND3X0_RVT U874 ( .A1(n443), .A2(n416), .A3(n442), .Y(a2stg_frac1_in[25])
         );
  AOI22X1_RVT U875 ( .A1(n1027), .A2(a1stg_in1[15]), .A3(n470), .A4(
        a1stg_in1[14]), .Y(n445) );
  AO222X1_RVT U876 ( .A1(a1stg_intlngop), .A2(a1stg_in2[26]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[14]), .A5(a1stg_in2[15]), .A6(
        a1stg_norm_dbl_in2), .Y(n1096) );
  NAND2X0_RVT U877 ( .A1(n1030), .A2(n1096), .Y(n444) );
  NAND3X0_RVT U878 ( .A1(n445), .A2(n416), .A3(n444), .Y(a2stg_frac1_in[26])
         );
  AOI22X1_RVT U879 ( .A1(n1027), .A2(a1stg_in1[16]), .A3(n470), .A4(
        a1stg_in1[15]), .Y(n447) );
  AO222X1_RVT U880 ( .A1(a1stg_intlngop), .A2(a1stg_in2[27]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[15]), .A5(a1stg_in2[16]), .A6(
        a1stg_norm_dbl_in2), .Y(n1095) );
  NAND2X0_RVT U881 ( .A1(n1030), .A2(n1095), .Y(n446) );
  NAND3X0_RVT U882 ( .A1(n447), .A2(n416), .A3(n446), .Y(a2stg_frac1_in[27])
         );
  AOI22X1_RVT U883 ( .A1(n1027), .A2(a1stg_in1[17]), .A3(n470), .A4(
        a1stg_in1[16]), .Y(n449) );
  AO222X1_RVT U884 ( .A1(a1stg_intlngop), .A2(a1stg_in2[28]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[16]), .A5(a1stg_in2[17]), .A6(
        a1stg_norm_dbl_in2), .Y(n1094) );
  NAND2X0_RVT U885 ( .A1(n1030), .A2(n1094), .Y(n448) );
  NAND3X0_RVT U886 ( .A1(n449), .A2(n416), .A3(n448), .Y(a2stg_frac1_in[28])
         );
  AOI22X1_RVT U887 ( .A1(n1027), .A2(a1stg_in1[18]), .A3(n470), .A4(
        a1stg_in1[17]), .Y(n451) );
  AO222X1_RVT U888 ( .A1(a1stg_intlngop), .A2(a1stg_in2[29]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[17]), .A5(a1stg_in2[18]), .A6(
        a1stg_norm_dbl_in2), .Y(n1093) );
  NAND2X0_RVT U889 ( .A1(n1030), .A2(n1093), .Y(n450) );
  NAND3X0_RVT U890 ( .A1(n451), .A2(n416), .A3(n450), .Y(a2stg_frac1_in[29])
         );
  AOI22X1_RVT U891 ( .A1(n1027), .A2(a1stg_in1[19]), .A3(n470), .A4(
        a1stg_in1[18]), .Y(n453) );
  AO222X1_RVT U892 ( .A1(a1stg_intlngop), .A2(a1stg_in2[30]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[18]), .A5(a1stg_in2[19]), .A6(
        a1stg_norm_dbl_in2), .Y(n1092) );
  NAND2X0_RVT U893 ( .A1(n1030), .A2(n1092), .Y(n452) );
  NAND3X0_RVT U894 ( .A1(n453), .A2(n416), .A3(n452), .Y(a2stg_frac1_in[30])
         );
  AOI22X1_RVT U895 ( .A1(n1027), .A2(a1stg_in1[20]), .A3(n470), .A4(
        a1stg_in1[19]), .Y(n455) );
  AO222X1_RVT U896 ( .A1(a1stg_intlngop), .A2(a1stg_in2[31]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[19]), .A5(a1stg_in2[20]), .A6(
        a1stg_norm_dbl_in2), .Y(n1091) );
  NAND2X0_RVT U897 ( .A1(n1030), .A2(n1091), .Y(n454) );
  NAND3X0_RVT U898 ( .A1(n455), .A2(n416), .A3(n454), .Y(a2stg_frac1_in[31])
         );
  AOI22X1_RVT U899 ( .A1(n1027), .A2(a1stg_in1[21]), .A3(n470), .A4(
        a1stg_in1[20]), .Y(n457) );
  AO222X1_RVT U900 ( .A1(a1stg_intlngop), .A2(a1stg_in2[32]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[20]), .A5(a1stg_in2[21]), .A6(
        a1stg_norm_dbl_in2), .Y(n1090) );
  NAND2X0_RVT U901 ( .A1(n1030), .A2(n1090), .Y(n456) );
  NAND3X0_RVT U902 ( .A1(n457), .A2(n416), .A3(n456), .Y(a2stg_frac1_in[32])
         );
  AOI22X1_RVT U903 ( .A1(n1027), .A2(a1stg_in1[22]), .A3(n470), .A4(
        a1stg_in1[21]), .Y(n459) );
  AO222X1_RVT U904 ( .A1(a1stg_intlngop), .A2(a1stg_in2[33]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[21]), .A5(a1stg_in2[22]), .A6(
        a1stg_norm_dbl_in2), .Y(n1089) );
  NAND2X0_RVT U905 ( .A1(n1030), .A2(n1089), .Y(n458) );
  NAND3X0_RVT U906 ( .A1(n459), .A2(n416), .A3(n458), .Y(a2stg_frac1_in[33])
         );
  AOI22X1_RVT U907 ( .A1(n1027), .A2(a1stg_in1[23]), .A3(n470), .A4(
        a1stg_in1[22]), .Y(n461) );
  AO222X1_RVT U908 ( .A1(a1stg_intlngop), .A2(a1stg_in2[34]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[22]), .A5(a1stg_in2[23]), .A6(
        a1stg_norm_dbl_in2), .Y(n1088) );
  NAND2X0_RVT U909 ( .A1(n1030), .A2(n1088), .Y(n460) );
  NAND3X0_RVT U910 ( .A1(n461), .A2(n416), .A3(n460), .Y(a2stg_frac1_in[34])
         );
  AOI22X1_RVT U911 ( .A1(n1027), .A2(a1stg_in1[24]), .A3(n470), .A4(
        a1stg_in1[23]), .Y(n463) );
  AO222X1_RVT U912 ( .A1(a1stg_intlngop), .A2(a1stg_in2[35]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[23]), .A5(a1stg_in2[24]), .A6(
        a1stg_norm_dbl_in2), .Y(n1087) );
  NAND2X0_RVT U913 ( .A1(n1030), .A2(n1087), .Y(n462) );
  NAND3X0_RVT U914 ( .A1(n463), .A2(n416), .A3(n462), .Y(a2stg_frac1_in[35])
         );
  AOI22X1_RVT U915 ( .A1(n1027), .A2(a1stg_in1[25]), .A3(n470), .A4(
        a1stg_in1[24]), .Y(n465) );
  AO222X1_RVT U916 ( .A1(a1stg_intlngop), .A2(a1stg_in2[36]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[24]), .A5(a1stg_in2[25]), .A6(
        a1stg_norm_dbl_in2), .Y(n1086) );
  NAND2X0_RVT U917 ( .A1(n1030), .A2(n1086), .Y(n464) );
  NAND3X0_RVT U918 ( .A1(n465), .A2(n416), .A3(n464), .Y(a2stg_frac1_in[36])
         );
  AOI22X1_RVT U919 ( .A1(n1027), .A2(a1stg_in1[26]), .A3(n470), .A4(
        a1stg_in1[25]), .Y(n467) );
  AO222X1_RVT U920 ( .A1(a1stg_intlngop), .A2(a1stg_in2[37]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[25]), .A5(a1stg_in2[26]), .A6(
        a1stg_norm_dbl_in2), .Y(n1085) );
  NAND2X0_RVT U921 ( .A1(n1030), .A2(n1085), .Y(n466) );
  NAND3X0_RVT U922 ( .A1(n467), .A2(n416), .A3(n466), .Y(a2stg_frac1_in[37])
         );
  AOI22X1_RVT U923 ( .A1(n1027), .A2(a1stg_in1[27]), .A3(n470), .A4(
        a1stg_in1[26]), .Y(n469) );
  AO222X1_RVT U924 ( .A1(a1stg_intlngop), .A2(a1stg_in2[38]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[26]), .A5(a1stg_in2[27]), .A6(
        a1stg_norm_dbl_in2), .Y(n1084) );
  NAND2X0_RVT U925 ( .A1(n1030), .A2(n1084), .Y(n468) );
  NAND3X0_RVT U926 ( .A1(n469), .A2(n416), .A3(n468), .Y(a2stg_frac1_in[38])
         );
  AOI22X1_RVT U927 ( .A1(a1stg_in1[28]), .A2(n1027), .A3(a1stg_in1[27]), .A4(
        n470), .Y(n472) );
  AO222X1_RVT U928 ( .A1(a1stg_intlngop), .A2(a1stg_in2[39]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[27]), .A5(a1stg_in2[28]), .A6(
        a1stg_norm_dbl_in2), .Y(n1083) );
  NAND2X0_RVT U929 ( .A1(n1030), .A2(n1083), .Y(n471) );
  NAND3X0_RVT U930 ( .A1(n472), .A2(n416), .A3(n471), .Y(a2stg_frac1_in[39])
         );
  AOI22X1_RVT U931 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[0]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[11]), .Y(n475) );
  AND2X1_RVT U932 ( .A1(a5stg_to_0), .A2(a5stg_in_of), .Y(n1918) );
  INVX1_RVT U933 ( .A(n1918), .Y(n474) );
  NAND2X0_RVT U934 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[11]), .Y(n473) );
  NAND3X0_RVT U935 ( .A1(n475), .A2(n474), .A3(n473), .Y(add_frac_out[11]) );
  AOI22X1_RVT U936 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[1]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[12]), .Y(n477) );
  NAND2X0_RVT U937 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[12]), .Y(n476) );
  NAND3X0_RVT U938 ( .A1(n477), .A2(n474), .A3(n476), .Y(add_frac_out[12]) );
  AOI22X1_RVT U939 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[2]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[13]), .Y(n479) );
  NAND2X0_RVT U940 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[13]), .Y(n478) );
  NAND3X0_RVT U941 ( .A1(n479), .A2(n474), .A3(n478), .Y(add_frac_out[13]) );
  AOI22X1_RVT U942 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[3]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[14]), .Y(n481) );
  NAND2X0_RVT U943 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[14]), .Y(n480) );
  NAND3X0_RVT U944 ( .A1(n481), .A2(n474), .A3(n480), .Y(add_frac_out[14]) );
  AOI22X1_RVT U945 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[4]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[15]), .Y(n483) );
  NAND2X0_RVT U946 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[15]), .Y(n482) );
  NAND3X0_RVT U947 ( .A1(n483), .A2(n474), .A3(n482), .Y(add_frac_out[15]) );
  AOI22X1_RVT U948 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[5]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[16]), .Y(n485) );
  NAND2X0_RVT U949 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[16]), .Y(n484) );
  NAND3X0_RVT U950 ( .A1(n485), .A2(n474), .A3(n484), .Y(add_frac_out[16]) );
  AOI22X1_RVT U951 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[6]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[17]), .Y(n487) );
  NAND2X0_RVT U952 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[17]), .Y(n486) );
  NAND3X0_RVT U953 ( .A1(n487), .A2(n474), .A3(n486), .Y(add_frac_out[17]) );
  AOI22X1_RVT U954 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[7]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[18]), .Y(n489) );
  NAND2X0_RVT U955 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[18]), .Y(n488) );
  NAND3X0_RVT U956 ( .A1(n489), .A2(n474), .A3(n488), .Y(add_frac_out[18]) );
  AOI22X1_RVT U957 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[8]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[19]), .Y(n491) );
  NAND2X0_RVT U958 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[19]), .Y(n490) );
  NAND3X0_RVT U959 ( .A1(n491), .A2(n474), .A3(n490), .Y(add_frac_out[19]) );
  AOI22X1_RVT U960 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[9]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[20]), .Y(n493) );
  NAND2X0_RVT U961 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[20]), .Y(n492) );
  NAND3X0_RVT U962 ( .A1(n493), .A2(n474), .A3(n492), .Y(add_frac_out[20]) );
  AOI22X1_RVT U963 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[10]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[21]), .Y(n495) );
  NAND2X0_RVT U964 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[21]), .Y(n494) );
  NAND3X0_RVT U965 ( .A1(n495), .A2(n474), .A3(n494), .Y(add_frac_out[21]) );
  AOI22X1_RVT U966 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[11]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[22]), .Y(n497) );
  NAND2X0_RVT U967 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[22]), .Y(n496) );
  NAND3X0_RVT U968 ( .A1(n497), .A2(n474), .A3(n496), .Y(add_frac_out[22]) );
  AOI22X1_RVT U969 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[12]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[23]), .Y(n499) );
  NAND2X0_RVT U970 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[23]), .Y(n498) );
  NAND3X0_RVT U971 ( .A1(n499), .A2(n474), .A3(n498), .Y(add_frac_out[23]) );
  AOI22X1_RVT U972 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[13]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[24]), .Y(n501) );
  NAND2X0_RVT U973 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[24]), .Y(n500) );
  NAND3X0_RVT U974 ( .A1(n501), .A2(n474), .A3(n500), .Y(add_frac_out[24]) );
  AOI22X1_RVT U975 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[14]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[25]), .Y(n503) );
  NAND2X0_RVT U976 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[25]), .Y(n502) );
  NAND3X0_RVT U977 ( .A1(n503), .A2(n474), .A3(n502), .Y(add_frac_out[25]) );
  AOI22X1_RVT U978 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[15]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[26]), .Y(n505) );
  NAND2X0_RVT U979 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[26]), .Y(n504) );
  NAND3X0_RVT U980 ( .A1(n505), .A2(n474), .A3(n504), .Y(add_frac_out[26]) );
  AOI22X1_RVT U981 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[16]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[27]), .Y(n507) );
  NAND2X0_RVT U982 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[27]), .Y(n506) );
  NAND3X0_RVT U983 ( .A1(n507), .A2(n474), .A3(n506), .Y(add_frac_out[27]) );
  AOI22X1_RVT U984 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[17]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[28]), .Y(n509) );
  NAND2X0_RVT U985 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[28]), .Y(n508) );
  NAND3X0_RVT U986 ( .A1(n509), .A2(n474), .A3(n508), .Y(add_frac_out[28]) );
  AOI22X1_RVT U987 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[18]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[29]), .Y(n511) );
  NAND2X0_RVT U988 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[29]), .Y(n510) );
  NAND3X0_RVT U989 ( .A1(n511), .A2(n474), .A3(n510), .Y(add_frac_out[29]) );
  AOI22X1_RVT U990 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[19]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[30]), .Y(n513) );
  NAND2X0_RVT U991 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[30]), .Y(n512) );
  NAND3X0_RVT U992 ( .A1(n513), .A2(n474), .A3(n512), .Y(add_frac_out[30]) );
  AOI22X1_RVT U993 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[20]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[31]), .Y(n515) );
  NAND2X0_RVT U994 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[31]), .Y(n514) );
  NAND3X0_RVT U995 ( .A1(n515), .A2(n474), .A3(n514), .Y(add_frac_out[31]) );
  AOI22X1_RVT U996 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[21]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[32]), .Y(n517) );
  NAND2X0_RVT U997 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[32]), .Y(n516) );
  NAND3X0_RVT U998 ( .A1(n517), .A2(n474), .A3(n516), .Y(add_frac_out[32]) );
  AOI22X1_RVT U999 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[22]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[33]), .Y(n519) );
  NAND2X0_RVT U1000 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[33]), .Y(n518) );
  NAND3X0_RVT U1001 ( .A1(n519), .A2(n474), .A3(n518), .Y(add_frac_out[33]) );
  AOI22X1_RVT U1002 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[23]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[34]), .Y(n521) );
  NAND2X0_RVT U1003 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[34]), .Y(n520) );
  NAND3X0_RVT U1004 ( .A1(n521), .A2(n474), .A3(n520), .Y(add_frac_out[34]) );
  AOI22X1_RVT U1005 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[24]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[35]), .Y(n523) );
  NAND2X0_RVT U1006 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[35]), .Y(n522) );
  NAND3X0_RVT U1007 ( .A1(n523), .A2(n474), .A3(n522), .Y(add_frac_out[35]) );
  AOI22X1_RVT U1008 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[25]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[36]), .Y(n525) );
  NAND2X0_RVT U1009 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[36]), .Y(n524) );
  NAND3X0_RVT U1010 ( .A1(n525), .A2(n474), .A3(n524), .Y(add_frac_out[36]) );
  AOI22X1_RVT U1011 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[26]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[37]), .Y(n527) );
  NAND2X0_RVT U1012 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[37]), .Y(n526) );
  NAND3X0_RVT U1013 ( .A1(n527), .A2(n474), .A3(n526), .Y(add_frac_out[37]) );
  AOI22X1_RVT U1014 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[27]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[38]), .Y(n529) );
  NAND2X0_RVT U1015 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[38]), .Y(n528) );
  NAND3X0_RVT U1016 ( .A1(n529), .A2(n474), .A3(n528), .Y(add_frac_out[38]) );
  AOI22X1_RVT U1017 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[28]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[39]), .Y(n531) );
  NAND2X0_RVT U1018 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[39]), .Y(n530) );
  NAND3X0_RVT U1019 ( .A1(n531), .A2(n474), .A3(n530), .Y(add_frac_out[39]) );
  AOI22X1_RVT U1020 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[29]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[40]), .Y(n533) );
  NAND2X0_RVT U1021 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[40]), .Y(n532) );
  NAND3X0_RVT U1022 ( .A1(n533), .A2(n474), .A3(n532), .Y(add_frac_out[40]) );
  AOI22X1_RVT U1023 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[30]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[41]), .Y(n535) );
  NAND2X0_RVT U1024 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[41]), .Y(n534) );
  NAND3X0_RVT U1025 ( .A1(n535), .A2(n474), .A3(n534), .Y(add_frac_out[41]) );
  AOI22X1_RVT U1026 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[31]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[42]), .Y(n537) );
  NAND2X0_RVT U1027 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[42]), .Y(n536) );
  NAND3X0_RVT U1028 ( .A1(n537), .A2(n474), .A3(n536), .Y(add_frac_out[42]) );
  AOI22X1_RVT U1029 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[32]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[43]), .Y(n539) );
  NAND2X0_RVT U1030 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[43]), .Y(n538) );
  NAND3X0_RVT U1031 ( .A1(n539), .A2(n474), .A3(n538), .Y(add_frac_out[43]) );
  AOI22X1_RVT U1032 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[33]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[44]), .Y(n541) );
  NAND2X0_RVT U1033 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[44]), .Y(n540) );
  NAND3X0_RVT U1034 ( .A1(n541), .A2(n474), .A3(n540), .Y(add_frac_out[44]) );
  AOI22X1_RVT U1035 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[34]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[45]), .Y(n543) );
  NAND2X0_RVT U1036 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[45]), .Y(n542) );
  NAND3X0_RVT U1037 ( .A1(n543), .A2(n474), .A3(n542), .Y(add_frac_out[45]) );
  AOI22X1_RVT U1038 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[35]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[46]), .Y(n545) );
  NAND2X0_RVT U1039 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[46]), .Y(n544) );
  NAND3X0_RVT U1040 ( .A1(n545), .A2(n474), .A3(n544), .Y(add_frac_out[46]) );
  AOI22X1_RVT U1041 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[36]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[47]), .Y(n547) );
  NAND2X0_RVT U1042 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[47]), .Y(n546) );
  NAND3X0_RVT U1043 ( .A1(n547), .A2(n474), .A3(n546), .Y(add_frac_out[47]) );
  AOI22X1_RVT U1044 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[37]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[48]), .Y(n549) );
  NAND2X0_RVT U1045 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[48]), .Y(n548) );
  NAND3X0_RVT U1046 ( .A1(n549), .A2(n474), .A3(n548), .Y(add_frac_out[48]) );
  AOI22X1_RVT U1047 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[38]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[49]), .Y(n551) );
  NAND2X0_RVT U1048 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[49]), .Y(n550) );
  NAND3X0_RVT U1049 ( .A1(n551), .A2(n474), .A3(n550), .Y(add_frac_out[49]) );
  AOI22X1_RVT U1050 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[39]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[50]), .Y(n553) );
  NAND2X0_RVT U1051 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[50]), .Y(n552) );
  NAND3X0_RVT U1052 ( .A1(n553), .A2(n474), .A3(n552), .Y(add_frac_out[50]) );
  AOI22X1_RVT U1053 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[40]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[51]), .Y(n555) );
  NAND2X0_RVT U1054 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[51]), .Y(n554) );
  NAND3X0_RVT U1055 ( .A1(n555), .A2(n474), .A3(n554), .Y(add_frac_out[51]) );
  AOI22X1_RVT U1056 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[41]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[52]), .Y(n557) );
  NAND2X0_RVT U1057 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[52]), .Y(n556) );
  NAND3X0_RVT U1058 ( .A1(n557), .A2(n474), .A3(n556), .Y(add_frac_out[52]) );
  AOI22X1_RVT U1059 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[42]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[53]), .Y(n559) );
  NAND2X0_RVT U1060 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[53]), .Y(n558) );
  NAND3X0_RVT U1061 ( .A1(n559), .A2(n474), .A3(n558), .Y(add_frac_out[53]) );
  AOI22X1_RVT U1062 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[43]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[54]), .Y(n561) );
  NAND2X0_RVT U1063 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[54]), .Y(n560) );
  NAND3X0_RVT U1064 ( .A1(n561), .A2(n474), .A3(n560), .Y(add_frac_out[54]) );
  AOI22X1_RVT U1065 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[44]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[55]), .Y(n563) );
  NAND2X0_RVT U1066 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[55]), .Y(n562) );
  NAND3X0_RVT U1067 ( .A1(n563), .A2(n474), .A3(n562), .Y(add_frac_out[55]) );
  AOI22X1_RVT U1068 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[45]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[56]), .Y(n565) );
  NAND2X0_RVT U1069 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[56]), .Y(n564) );
  NAND3X0_RVT U1070 ( .A1(n565), .A2(n474), .A3(n564), .Y(add_frac_out[56]) );
  AOI22X1_RVT U1071 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[46]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[57]), .Y(n567) );
  NAND2X0_RVT U1072 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[57]), .Y(n566) );
  NAND3X0_RVT U1073 ( .A1(n567), .A2(n474), .A3(n566), .Y(add_frac_out[57]) );
  AOI22X1_RVT U1074 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[47]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[58]), .Y(n569) );
  NAND2X0_RVT U1075 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[58]), .Y(n568) );
  NAND3X0_RVT U1076 ( .A1(n569), .A2(n474), .A3(n568), .Y(add_frac_out[58]) );
  AOI22X1_RVT U1077 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[48]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[59]), .Y(n571) );
  NAND2X0_RVT U1078 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[59]), .Y(n570) );
  NAND3X0_RVT U1079 ( .A1(n571), .A2(n474), .A3(n570), .Y(add_frac_out[59]) );
  AOI22X1_RVT U1080 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[49]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[60]), .Y(n573) );
  NAND2X0_RVT U1081 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[60]), .Y(n572) );
  NAND3X0_RVT U1082 ( .A1(n573), .A2(n474), .A3(n572), .Y(add_frac_out[60]) );
  AOI22X1_RVT U1083 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[50]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[61]), .Y(n575) );
  NAND2X0_RVT U1084 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[61]), .Y(n574) );
  NAND3X0_RVT U1085 ( .A1(n575), .A2(n474), .A3(n574), .Y(add_frac_out[61]) );
  AOI22X1_RVT U1086 ( .A1(a5stg_frac_out_rndadd), .A2(a5stg_rndadd[51]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[62]), .Y(n577) );
  NAND2X0_RVT U1087 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[62]), .Y(n576) );
  NAND3X0_RVT U1088 ( .A1(n577), .A2(n474), .A3(n576), .Y(add_frac_out[62]) );
  OA21X1_RVT U1089 ( .A1(n579), .A2(a4stg_rnd_frac_62), .A3(n578), .Y(
        a4stg_rndadd_tmp[51]) );
  OA21X1_RVT U1090 ( .A1(n581), .A2(a4stg_rnd_frac_61), .A3(n580), .Y(
        a4stg_rndadd_tmp[50]) );
  OA21X1_RVT U1091 ( .A1(n583), .A2(a4stg_rnd_frac_60), .A3(n582), .Y(
        a4stg_rndadd_tmp[49]) );
  OA21X1_RVT U1092 ( .A1(n585), .A2(a4stg_rnd_frac_59), .A3(n584), .Y(
        a4stg_rndadd_tmp[48]) );
  OA21X1_RVT U1093 ( .A1(n587), .A2(a4stg_rnd_frac_58), .A3(n586), .Y(
        a4stg_rndadd_tmp[47]) );
  OA21X1_RVT U1094 ( .A1(n589), .A2(a4stg_rnd_frac_57), .A3(n588), .Y(
        a4stg_rndadd_tmp[46]) );
  OA21X1_RVT U1095 ( .A1(n591), .A2(a4stg_rnd_frac_56), .A3(n590), .Y(
        a4stg_rndadd_tmp[45]) );
  OA21X1_RVT U1096 ( .A1(n593), .A2(a4stg_rnd_frac_55), .A3(n592), .Y(
        a4stg_rndadd_tmp[44]) );
  OA21X1_RVT U1097 ( .A1(n595), .A2(a4stg_rnd_frac_54), .A3(n594), .Y(
        a4stg_rndadd_tmp[43]) );
  OA21X1_RVT U1098 ( .A1(n597), .A2(a4stg_rnd_frac_53), .A3(n596), .Y(
        a4stg_rndadd_tmp[42]) );
  OA21X1_RVT U1099 ( .A1(n599), .A2(a4stg_rnd_frac_52), .A3(n598), .Y(
        a4stg_rndadd_tmp[41]) );
  OA21X1_RVT U1100 ( .A1(n601), .A2(a4stg_rnd_frac_51), .A3(n600), .Y(
        a4stg_rndadd_tmp[40]) );
  OA21X1_RVT U1101 ( .A1(n603), .A2(a4stg_rnd_frac_50), .A3(n602), .Y(
        a4stg_rndadd_tmp[39]) );
  OA21X1_RVT U1102 ( .A1(n605), .A2(a4stg_rnd_frac_49), .A3(n604), .Y(
        a4stg_rndadd_tmp[38]) );
  OA21X1_RVT U1103 ( .A1(n607), .A2(a4stg_rnd_frac_48), .A3(n606), .Y(
        a4stg_rndadd_tmp[37]) );
  OA21X1_RVT U1104 ( .A1(n609), .A2(a4stg_rnd_frac_47), .A3(n608), .Y(
        a4stg_rndadd_tmp[36]) );
  OA21X1_RVT U1105 ( .A1(n611), .A2(a4stg_rnd_frac_46), .A3(n610), .Y(
        a4stg_rndadd_tmp[35]) );
  OA21X1_RVT U1106 ( .A1(n613), .A2(a4stg_rnd_frac_45), .A3(n612), .Y(
        a4stg_rndadd_tmp[34]) );
  OA21X1_RVT U1107 ( .A1(n615), .A2(a4stg_rnd_frac_44), .A3(n614), .Y(
        a4stg_rndadd_tmp[33]) );
  NAND3X0_RVT U1108 ( .A1(n620), .A2(a4stg_rnd_frac_42), .A3(a4stg_rnd_frac_41), .Y(n618) );
  OA21X1_RVT U1109 ( .A1(n617), .A2(a4stg_rnd_frac_43), .A3(n616), .Y(
        a4stg_rndadd_tmp[32]) );
  OA221X1_RVT U1110 ( .A1(a4stg_rnd_frac_42), .A2(n620), .A3(a4stg_rnd_frac_42), .A4(a4stg_rnd_frac_41), .A5(n618), .Y(a4stg_rndadd_tmp[31]) );
  NAND2X0_RVT U1111 ( .A1(n620), .A2(a4stg_rnd_frac_41), .Y(n619) );
  OA21X1_RVT U1112 ( .A1(n620), .A2(a4stg_rnd_frac_41), .A3(n619), .Y(
        a4stg_rndadd_tmp[30]) );
  FADDX1_RVT U1113 ( .A(a4stg_rnd_sng), .B(a4stg_rnd_frac_40), .CI(n621), .CO(
        n620), .S(a4stg_rndadd_tmp[29]) );
  OA21X1_RVT U1114 ( .A1(n623), .A2(a4stg_rnd_frac_39), .A3(n622), .Y(
        a4stg_rndadd_tmp[28]) );
  OA21X1_RVT U1115 ( .A1(n625), .A2(a4stg_rnd_frac[38]), .A3(n624), .Y(
        a4stg_rndadd_tmp[27]) );
  OA21X1_RVT U1116 ( .A1(n627), .A2(a4stg_rnd_frac[37]), .A3(n626), .Y(
        a4stg_rndadd_tmp[26]) );
  OA21X1_RVT U1117 ( .A1(n629), .A2(a4stg_rnd_frac[36]), .A3(n628), .Y(
        a4stg_rndadd_tmp[25]) );
  OA21X1_RVT U1118 ( .A1(n631), .A2(a4stg_rnd_frac[35]), .A3(n630), .Y(
        a4stg_rndadd_tmp[24]) );
  OA21X1_RVT U1119 ( .A1(n633), .A2(a4stg_rnd_frac[34]), .A3(n632), .Y(
        a4stg_rndadd_tmp[23]) );
  OA21X1_RVT U1120 ( .A1(n635), .A2(a4stg_rnd_frac[33]), .A3(n634), .Y(
        a4stg_rndadd_tmp[22]) );
  OA21X1_RVT U1121 ( .A1(n637), .A2(a4stg_rnd_frac[32]), .A3(n636), .Y(
        a4stg_rndadd_tmp[21]) );
  OA21X1_RVT U1122 ( .A1(n639), .A2(a4stg_rnd_frac[31]), .A3(n638), .Y(
        a4stg_rndadd_tmp[20]) );
  OA21X1_RVT U1123 ( .A1(n641), .A2(a4stg_rnd_frac[30]), .A3(n640), .Y(
        a4stg_rndadd_tmp[19]) );
  OA21X1_RVT U1124 ( .A1(n643), .A2(a4stg_rnd_frac[29]), .A3(n642), .Y(
        a4stg_rndadd_tmp[18]) );
  OA21X1_RVT U1125 ( .A1(n645), .A2(a4stg_rnd_frac[28]), .A3(n644), .Y(
        a4stg_rndadd_tmp[17]) );
  OA21X1_RVT U1126 ( .A1(n647), .A2(a4stg_rnd_frac[27]), .A3(n646), .Y(
        a4stg_rndadd_tmp[16]) );
  OA21X1_RVT U1127 ( .A1(n649), .A2(a4stg_rnd_frac[26]), .A3(n648), .Y(
        a4stg_rndadd_tmp[15]) );
  OA21X1_RVT U1128 ( .A1(n651), .A2(a4stg_rnd_frac[25]), .A3(n650), .Y(
        a4stg_rndadd_tmp[14]) );
  OA21X1_RVT U1129 ( .A1(n653), .A2(a4stg_rnd_frac[24]), .A3(n652), .Y(
        a4stg_rndadd_tmp[13]) );
  OA21X1_RVT U1130 ( .A1(n655), .A2(a4stg_rnd_frac[23]), .A3(n654), .Y(
        a4stg_rndadd_tmp[12]) );
  OA21X1_RVT U1131 ( .A1(n657), .A2(a4stg_rnd_frac[22]), .A3(n656), .Y(
        a4stg_rndadd_tmp[11]) );
  OA21X1_RVT U1132 ( .A1(n659), .A2(a4stg_rnd_frac[21]), .A3(n658), .Y(
        a4stg_rndadd_tmp[10]) );
  OA21X1_RVT U1133 ( .A1(n661), .A2(a4stg_rnd_frac[20]), .A3(n660), .Y(
        a4stg_rndadd_tmp[9]) );
  OA21X1_RVT U1134 ( .A1(n663), .A2(a4stg_rnd_frac[19]), .A3(n662), .Y(
        a4stg_rndadd_tmp[8]) );
  OA21X1_RVT U1135 ( .A1(n665), .A2(a4stg_rnd_frac[18]), .A3(n664), .Y(
        a4stg_rndadd_tmp[7]) );
  OA21X1_RVT U1136 ( .A1(n667), .A2(a4stg_rnd_frac[17]), .A3(n666), .Y(
        a4stg_rndadd_tmp[6]) );
  OA21X1_RVT U1137 ( .A1(n669), .A2(a4stg_rnd_frac[16]), .A3(n668), .Y(
        a4stg_rndadd_tmp[5]) );
  OA21X1_RVT U1138 ( .A1(n671), .A2(a4stg_rnd_frac[15]), .A3(n670), .Y(
        a4stg_rndadd_tmp[4]) );
  OA21X1_RVT U1139 ( .A1(n673), .A2(a4stg_rnd_frac[14]), .A3(n672), .Y(
        a4stg_rndadd_tmp[3]) );
  NAND3X0_RVT U1140 ( .A1(a4stg_rnd_dbl), .A2(a4stg_rnd_frac[12]), .A3(
        a4stg_rnd_frac_11), .Y(n676) );
  OA21X1_RVT U1141 ( .A1(n675), .A2(a4stg_rnd_frac[13]), .A3(n674), .Y(
        a4stg_rndadd_tmp[2]) );
  OA221X1_RVT U1142 ( .A1(a4stg_rnd_frac[12]), .A2(a4stg_rnd_dbl), .A3(
        a4stg_rnd_frac[12]), .A4(a4stg_rnd_frac_11), .A5(n676), .Y(
        a4stg_rndadd_tmp[1]) );
  NAND2X0_RVT U1143 ( .A1(a4stg_rnd_dbl), .A2(a4stg_rnd_frac_11), .Y(n677) );
  OA21X1_RVT U1144 ( .A1(a4stg_rnd_dbl), .A2(a4stg_rnd_frac_11), .A3(n677), 
        .Y(a4stg_rndadd_tmp[0]) );
  INVX1_RVT U1146 ( .A(a2stg_shr_cnt_4[4]), .Y(n715) );
  AND2X1_RVT U1147 ( .A1(a2stg_shr_cnt_5_inv[0]), .A2(n715), .Y(n2045) );
  AND2X1_RVT U1148 ( .A1(a2stg_shr_cnt_5_inv[0]), .A2(a2stg_shr_cnt_4[0]), .Y(
        n2044) );
  AOI22X1_RVT U1149 ( .A1(a2stg_frac2a[43]), .A2(n2045), .A3(a2stg_frac2a[59]), 
        .A4(n2044), .Y(n2084) );
  INVX1_RVT U1150 ( .A(a2stg_shr_cnt_3[1]), .Y(n702) );
  INVX1_RVT U1151 ( .A(a2stg_shr_cnt_3[4]), .Y(n2449) );
  NAND2X0_RVT U1152 ( .A1(a2stg_shr_cnt_5_inv[0]), .A2(a2stg_shr_cnt_4[1]), 
        .Y(n693) );
  INVX1_RVT U1153 ( .A(n693), .Y(n701) );
  NAND2X0_RVT U1154 ( .A1(a2stg_shr_cnt_5_inv[1]), .A2(n715), .Y(n694) );
  INVX1_RVT U1155 ( .A(n694), .Y(n684) );
  AOI22X1_RVT U1156 ( .A1(a2stg_frac2a[51]), .A2(n701), .A3(a2stg_frac2a[35]), 
        .A4(n684), .Y(n683) );
  OA22X1_RVT U1157 ( .A1(n2084), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n683), 
        .Y(n2192) );
  NAND2X0_RVT U1158 ( .A1(a2stg_shr_cnt_2[1]), .A2(a2stg_shr_cnt_1[1]), .Y(
        n2467) );
  AOI22X1_RVT U1159 ( .A1(a2stg_frac2a[57]), .A2(n2044), .A3(a2stg_frac2a[41]), 
        .A4(n2045), .Y(n2104) );
  INVX1_RVT U1160 ( .A(a2stg_frac2a[49]), .Y(n2103) );
  INVX1_RVT U1161 ( .A(a2stg_frac2a[33]), .Y(n708) );
  OA22X1_RVT U1162 ( .A1(n2103), .A2(n693), .A3(n708), .A4(n694), .Y(n698) );
  OA22X1_RVT U1163 ( .A1(n2104), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n698), 
        .Y(n2211) );
  NAND2X0_RVT U1164 ( .A1(a2stg_shr_cnt_1[0]), .A2(a2stg_shr_cnt_2[0]), .Y(
        n2465) );
  OA22X1_RVT U1165 ( .A1(n2192), .A2(n2467), .A3(n2211), .A4(n2465), .Y(n679)
         );
  AOI22X1_RVT U1166 ( .A1(a2stg_frac2a[45]), .A2(n2045), .A3(a2stg_frac2a[61]), 
        .A4(n2044), .Y(n2065) );
  AOI22X1_RVT U1167 ( .A1(a2stg_frac2a[53]), .A2(n701), .A3(a2stg_frac2a[37]), 
        .A4(n684), .Y(n681) );
  OA22X1_RVT U1168 ( .A1(n2065), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n681), 
        .Y(n2167) );
  NAND2X0_RVT U1169 ( .A1(a2stg_shr_cnt_1[0]), .A2(a2stg_shr_cnt_2[1]), .Y(
        n2456) );
  AO22X1_RVT U1170 ( .A1(a2stg_frac2a[55]), .A2(n701), .A3(a2stg_frac2a[39]), 
        .A4(n684), .Y(n2121) );
  AND2X1_RVT U1171 ( .A1(a2stg_shr_cnt_5[1]), .A2(n715), .Y(n682) );
  AO222X1_RVT U1172 ( .A1(a2stg_frac2a[47]), .A2(n701), .A3(a2stg_frac2a[31]), 
        .A4(n684), .A5(a2stg_frac2a[63]), .A6(n682), .Y(n2245) );
  AOI22X1_RVT U1173 ( .A1(a2stg_shr_cnt_3[1]), .A2(n2121), .A3(n2449), .A4(
        n2245), .Y(n2227) );
  AND2X1_RVT U1174 ( .A1(a2stg_shr_cnt_2[0]), .A2(a2stg_shr_cnt_1[1]), .Y(
        n2450) );
  INVX1_RVT U1175 ( .A(n2450), .Y(n2448) );
  OA22X1_RVT U1176 ( .A1(n2167), .A2(n2456), .A3(n2227), .A4(n2448), .Y(n678)
         );
  NAND2X0_RVT U1177 ( .A1(n679), .A2(n678), .Y(n2181) );
  INVX1_RVT U1178 ( .A(n2181), .Y(n2191) );
  NAND2X0_RVT U1179 ( .A1(a2stg_shr_cnt_5_inv[1]), .A2(a2stg_shr_cnt_4[2]), 
        .Y(n699) );
  INVX1_RVT U1180 ( .A(n699), .Y(n716) );
  AO22X1_RVT U1181 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[50]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[18]), .Y(n821) );
  AO22X1_RVT U1182 ( .A1(a2stg_frac2a[34]), .A2(n716), .A3(n715), .A4(n821), 
        .Y(n2491) );
  INVX1_RVT U1183 ( .A(n2491), .Y(n2375) );
  AO22X1_RVT U1184 ( .A1(a2stg_shr_cnt_5[1]), .A2(a2stg_frac2a[58]), .A3(
        a2stg_shr_cnt_5_inv[1]), .A4(a2stg_frac2a[26]), .Y(n777) );
  NAND2X0_RVT U1185 ( .A1(a2stg_shr_cnt_5_inv[3]), .A2(n715), .Y(n713) );
  INVX1_RVT U1186 ( .A(n713), .Y(n717) );
  NAND2X0_RVT U1187 ( .A1(a2stg_shr_cnt_5[3]), .A2(n715), .Y(n712) );
  INVX1_RVT U1188 ( .A(n712), .Y(n718) );
  AOI222X1_RVT U1189 ( .A1(n777), .A2(a2stg_shr_cnt_4[3]), .A3(
        a2stg_frac2a[10]), .A4(n717), .A5(a2stg_frac2a[42]), .A6(n718), .Y(
        n2441) );
  AO22X1_RVT U1190 ( .A1(a2stg_frac2a[38]), .A2(n684), .A3(a2stg_frac2a[54]), 
        .A4(n701), .Y(n725) );
  AO222X1_RVT U1191 ( .A1(a2stg_frac2a[46]), .A2(n701), .A3(a2stg_frac2a[62]), 
        .A4(n682), .A5(n684), .A6(a2stg_frac2a[30]), .Y(n2253) );
  AO22X1_RVT U1192 ( .A1(a2stg_shr_cnt_3[1]), .A2(n725), .A3(n2449), .A4(n2253), .Y(n2199) );
  INVX1_RVT U1193 ( .A(n2199), .Y(n2235) );
  NAND2X0_RVT U1194 ( .A1(a2stg_shr_cnt_3[1]), .A2(n2121), .Y(n680) );
  NAND4X0_RVT U1195 ( .A1(n2375), .A2(n2441), .A3(n2235), .A4(n680), .Y(n688)
         );
  AO22X1_RVT U1196 ( .A1(a2stg_shr_cnt_5[1]), .A2(a2stg_frac2a[57]), .A3(
        a2stg_shr_cnt_5_inv[1]), .A4(a2stg_frac2a[25]), .Y(n773) );
  AOI222X1_RVT U1197 ( .A1(n773), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[41]), .A5(n717), .A6(a2stg_frac2a[9]), .Y(n2452) );
  AO22X1_RVT U1198 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[49]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[17]), .Y(n752) );
  INVX1_RVT U1199 ( .A(n752), .Y(n707) );
  OA22X1_RVT U1200 ( .A1(a2stg_shr_cnt_4[4]), .A2(n707), .A3(n708), .A4(n699), 
        .Y(n2487) );
  AO22X1_RVT U1201 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[55]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[23]), .Y(n767) );
  AOI222X1_RVT U1202 ( .A1(n767), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[39]), .A5(n717), .A6(a2stg_frac2a[7]), .Y(n2411) );
  AO22X1_RVT U1203 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[51]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[19]), .Y(n755) );
  AO22X1_RVT U1204 ( .A1(a2stg_frac2a[35]), .A2(n716), .A3(n715), .A4(n755), 
        .Y(n2494) );
  INVX1_RVT U1205 ( .A(n2494), .Y(n2367) );
  NAND4X0_RVT U1206 ( .A1(n2452), .A2(n2487), .A3(n2411), .A4(n2367), .Y(n687)
         );
  AO22X1_RVT U1207 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[52]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[20]), .Y(n759) );
  AOI22X1_RVT U1208 ( .A1(n715), .A2(n759), .A3(a2stg_frac2a[36]), .A4(n716), 
        .Y(n2357) );
  AO22X1_RVT U1209 ( .A1(a2stg_shr_cnt_5[1]), .A2(a2stg_frac2a[56]), .A3(
        a2stg_shr_cnt_5_inv[1]), .A4(a2stg_frac2a[24]), .Y(n770) );
  AOI222X1_RVT U1210 ( .A1(n770), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[40]), .A5(n717), .A6(a2stg_frac2a[8]), .Y(n2472) );
  AO22X1_RVT U1211 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[54]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[22]), .Y(n762) );
  AO22X1_RVT U1212 ( .A1(a2stg_frac2a[38]), .A2(n716), .A3(n715), .A4(n762), 
        .Y(n2255) );
  INVX1_RVT U1213 ( .A(n2255), .Y(n2336) );
  AO22X1_RVT U1214 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[46]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[14]), .Y(n734) );
  AND2X1_RVT U1215 ( .A1(a2stg_shr_cnt_5[1]), .A2(a2stg_shr_cnt_4[2]), .Y(n700) );
  AO222X1_RVT U1216 ( .A1(n715), .A2(n734), .A3(a2stg_frac2a[62]), .A4(n700), 
        .A5(n716), .A6(a2stg_frac2a[30]), .Y(n785) );
  INVX1_RVT U1217 ( .A(n785), .Y(n2405) );
  NAND4X0_RVT U1218 ( .A1(n2357), .A2(n2472), .A3(n2336), .A4(n2405), .Y(n686)
         );
  AOI222X1_RVT U1219 ( .A1(a2stg_frac2a[45]), .A2(n701), .A3(a2stg_frac2a[29]), 
        .A4(n684), .A5(a2stg_frac2a[61]), .A6(n682), .Y(n2267) );
  OA22X1_RVT U1220 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2267), .A3(n681), .A4(n702), 
        .Y(n2244) );
  AOI222X1_RVT U1221 ( .A1(a2stg_frac2a[44]), .A2(n701), .A3(a2stg_frac2a[28]), 
        .A4(n684), .A5(a2stg_frac2a[60]), .A6(n682), .Y(n2277) );
  AOI22X1_RVT U1222 ( .A1(a2stg_frac2a[36]), .A2(n684), .A3(a2stg_frac2a[52]), 
        .A4(n701), .Y(n689) );
  OA22X1_RVT U1223 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2277), .A3(n689), .A4(n702), 
        .Y(n2256) );
  AO22X1_RVT U1224 ( .A1(a2stg_shr_cnt_5[1]), .A2(a2stg_frac2a[59]), .A3(
        a2stg_shr_cnt_5_inv[1]), .A4(a2stg_frac2a[27]), .Y(n793) );
  AOI22X1_RVT U1225 ( .A1(n701), .A2(a2stg_frac2a[43]), .A3(n715), .A4(n793), 
        .Y(n2286) );
  OA22X1_RVT U1226 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2286), .A3(n683), .A4(n702), 
        .Y(n2268) );
  AOI22X1_RVT U1227 ( .A1(n701), .A2(a2stg_frac2a[42]), .A3(n777), .A4(n715), 
        .Y(n2295) );
  AOI22X1_RVT U1228 ( .A1(a2stg_frac2a[50]), .A2(n701), .A3(a2stg_frac2a[34]), 
        .A4(n684), .Y(n690) );
  OA22X1_RVT U1229 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2295), .A3(n690), .A4(n702), 
        .Y(n2278) );
  NAND4X0_RVT U1230 ( .A1(n2244), .A2(n2256), .A3(n2268), .A4(n2278), .Y(n685)
         );
  NOR4X1_RVT U1231 ( .A1(n688), .A2(n687), .A3(n686), .A4(n685), .Y(n730) );
  NAND2X0_RVT U1232 ( .A1(n2450), .A2(n2199), .Y(n692) );
  AOI22X1_RVT U1233 ( .A1(a2stg_frac2a[44]), .A2(n2045), .A3(a2stg_frac2a[60]), 
        .A4(n2044), .Y(n2075) );
  OA22X1_RVT U1234 ( .A1(n2075), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n689), 
        .Y(n2160) );
  AOI22X1_RVT U1235 ( .A1(a2stg_frac2a[58]), .A2(n2044), .A3(a2stg_frac2a[42]), 
        .A4(n2045), .Y(n2093) );
  OA22X1_RVT U1236 ( .A1(n2093), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n690), 
        .Y(n2200) );
  OA22X1_RVT U1237 ( .A1(n2160), .A2(n2456), .A3(n2200), .A4(n2467), .Y(n691)
         );
  AND2X1_RVT U1238 ( .A1(n692), .A2(n691), .Y(n697) );
  AOI22X1_RVT U1239 ( .A1(a2stg_frac2a[56]), .A2(n2044), .A3(a2stg_frac2a[40]), 
        .A4(n2045), .Y(n2113) );
  INVX1_RVT U1240 ( .A(a2stg_frac2a[32]), .Y(n711) );
  INVX1_RVT U1241 ( .A(a2stg_frac2a[48]), .Y(n2111) );
  OA22X1_RVT U1242 ( .A1(n711), .A2(n694), .A3(n2111), .A4(n693), .Y(n703) );
  OA22X1_RVT U1243 ( .A1(n2113), .A2(n702), .A3(a2stg_shr_cnt_3[4]), .A4(n703), 
        .Y(n2220) );
  INVX1_RVT U1244 ( .A(n2465), .Y(n2345) );
  NAND2X0_RVT U1245 ( .A1(n695), .A2(n2345), .Y(n696) );
  AND2X1_RVT U1246 ( .A1(n697), .A2(n696), .Y(n2206) );
  AOI22X1_RVT U1247 ( .A1(n701), .A2(a2stg_frac2a[41]), .A3(n715), .A4(n773), 
        .Y(n2305) );
  OA22X1_RVT U1248 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2305), .A3(n698), .A4(n702), 
        .Y(n2287) );
  AO22X1_RVT U1249 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[44]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[12]), .Y(n735) );
  AO222X1_RVT U1250 ( .A1(n735), .A2(n715), .A3(n716), .A4(a2stg_frac2a[28]), 
        .A5(n700), .A6(a2stg_frac2a[60]), .Y(n782) );
  INVX1_RVT U1251 ( .A(n782), .Y(n2424) );
  AO22X1_RVT U1252 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[48]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[16]), .Y(n765) );
  INVX1_RVT U1253 ( .A(n765), .Y(n709) );
  OA22X1_RVT U1254 ( .A1(a2stg_shr_cnt_4[4]), .A2(n709), .A3(n711), .A4(n699), 
        .Y(n2398) );
  AO22X1_RVT U1255 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[47]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[15]), .Y(n733) );
  AOI222X1_RVT U1256 ( .A1(n715), .A2(n733), .A3(a2stg_frac2a[31]), .A4(n716), 
        .A5(n700), .A6(a2stg_frac2a[63]), .Y(n2410) );
  AO22X1_RVT U1257 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[45]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[13]), .Y(n731) );
  AO222X1_RVT U1258 ( .A1(n715), .A2(n731), .A3(a2stg_frac2a[61]), .A4(n700), 
        .A5(n716), .A6(a2stg_frac2a[29]), .Y(n783) );
  INVX1_RVT U1259 ( .A(n783), .Y(n2416) );
  NAND4X0_RVT U1260 ( .A1(n2424), .A2(n2398), .A3(n2410), .A4(n2416), .Y(n2489) );
  NAND4X0_RVT U1261 ( .A1(n2192), .A2(n2200), .A3(n2211), .A4(n2220), .Y(n705)
         );
  AOI22X1_RVT U1262 ( .A1(n701), .A2(a2stg_frac2a[40]), .A3(n715), .A4(n770), 
        .Y(n2313) );
  OA22X1_RVT U1263 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2313), .A3(n703), .A4(n702), 
        .Y(n2296) );
  AO21X1_RVT U1264 ( .A1(a2stg_shr_cnt_2[1]), .A2(n705), .A3(n704), .Y(n706)
         );
  NOR4X1_RVT U1265 ( .A1(n2489), .A2(n2245), .A3(n2253), .A4(n706), .Y(n724)
         );
  AO22X1_RVT U1266 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[53]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[21]), .Y(n766) );
  AOI222X1_RVT U1267 ( .A1(n766), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[37]), .A5(n717), .A6(a2stg_frac2a[5]), .Y(n2417) );
  AOI222X1_RVT U1268 ( .A1(n755), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[35]), .A5(n717), .A6(a2stg_frac2a[3]), .Y(n2433) );
  NAND4X0_RVT U1269 ( .A1(n2305), .A2(n2313), .A3(n2417), .A4(n2433), .Y(n722)
         );
  NAND4X0_RVT U1270 ( .A1(n2267), .A2(n2277), .A3(n2286), .A4(n2295), .Y(n721)
         );
  AOI222X1_RVT U1271 ( .A1(n759), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[36]), .A5(n717), .A6(a2stg_frac2a[4]), .Y(n2425) );
  AOI222X1_RVT U1272 ( .A1(n821), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[34]), .A5(n717), .A6(a2stg_frac2a[2]), .Y(n2442) );
  INVX1_RVT U1273 ( .A(a2stg_frac2a[1]), .Y(n742) );
  OA222X1_RVT U1274 ( .A1(n713), .A2(n742), .A3(n712), .A4(n708), .A5(n710), 
        .A6(n707), .Y(n2451) );
  INVX1_RVT U1275 ( .A(a2stg_frac2a[0]), .Y(n736) );
  OA222X1_RVT U1276 ( .A1(n713), .A2(n736), .A3(n712), .A4(n711), .A5(n710), 
        .A6(n709), .Y(n2470) );
  NAND4X0_RVT U1277 ( .A1(n2425), .A2(n2442), .A3(n2451), .A4(n2470), .Y(n720)
         );
  AO22X1_RVT U1278 ( .A1(a2stg_shr_cnt_5[2]), .A2(a2stg_frac2a[43]), .A3(
        a2stg_shr_cnt_5_inv[2]), .A4(a2stg_frac2a[11]), .Y(n714) );
  AOI22X1_RVT U1279 ( .A1(a2stg_shr_cnt_4[2]), .A2(n793), .A3(n715), .A4(n714), 
        .Y(n2432) );
  AOI22X1_RVT U1280 ( .A1(a2stg_frac2a[37]), .A2(n716), .A3(n715), .A4(n766), 
        .Y(n2349) );
  AO22X1_RVT U1281 ( .A1(a2stg_frac2a[39]), .A2(n716), .A3(n715), .A4(n767), 
        .Y(n2246) );
  INVX1_RVT U1282 ( .A(n2246), .Y(n2322) );
  AOI222X1_RVT U1283 ( .A1(n762), .A2(a2stg_shr_cnt_4[3]), .A3(n718), .A4(
        a2stg_frac2a[38]), .A5(n717), .A6(a2stg_frac2a[6]), .Y(n2406) );
  NAND4X0_RVT U1284 ( .A1(n2432), .A2(n2349), .A3(n2322), .A4(n2406), .Y(n719)
         );
  NOR4X1_RVT U1285 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .Y(n723) );
  AND4X1_RVT U1286 ( .A1(n2206), .A2(n2287), .A3(n724), .A4(n723), .Y(n729) );
  OA22X1_RVT U1287 ( .A1(n2160), .A2(n2467), .A3(n2220), .A4(n2448), .Y(n727)
         );
  AO22X1_RVT U1288 ( .A1(a2stg_frac2a[46]), .A2(n2045), .A3(a2stg_frac2a[62]), 
        .A4(n2044), .Y(n2053) );
  AOI22X1_RVT U1289 ( .A1(a2stg_shr_cnt_3[1]), .A2(n2053), .A3(n2449), .A4(
        n725), .Y(n2158) );
  OA22X1_RVT U1290 ( .A1(n2158), .A2(n2456), .A3(n2200), .A4(n2465), .Y(n726)
         );
  NAND2X0_RVT U1291 ( .A1(n727), .A2(n726), .Y(n2186) );
  NAND2X0_RVT U1292 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2186), .Y(n728) );
  NAND4X0_RVT U1293 ( .A1(n2191), .A2(n730), .A3(n729), .A4(n728), .Y(
        a2stg_fsdtoi_nx) );
  OR4X1_RVT U1294 ( .A1(a2stg_frac2a[10]), .A2(a2stg_frac2a[9]), .A3(
        a2stg_frac2a[11]), .A4(n731), .Y(n732) );
  OR4X1_RVT U1295 ( .A1(n735), .A2(n734), .A3(n733), .A4(n732), .Y(n751) );
  NOR4X1_RVT U1296 ( .A1(a2stg_frac2a[30]), .A2(a2stg_frac2a[25]), .A3(
        a2stg_frac2a[17]), .A4(a2stg_frac2a[23]), .Y(n749) );
  NOR4X1_RVT U1297 ( .A1(a2stg_frac2a[8]), .A2(a2stg_frac2a[16]), .A3(
        a2stg_frac2a[22]), .A4(a2stg_frac2a[14]), .Y(n748) );
  NOR3X0_RVT U1298 ( .A1(a2stg_frac2a[10]), .A2(a2stg_frac2a[9]), .A3(
        a2stg_frac2a[11]), .Y(n739) );
  NOR4X1_RVT U1299 ( .A1(a2stg_frac2a[20]), .A2(a2stg_frac2a[12]), .A3(
        a2stg_frac2a[28]), .A4(a2stg_frac2a[24]), .Y(n738) );
  NAND4X0_RVT U1300 ( .A1(n739), .A2(n738), .A3(n737), .A4(n736), .Y(n740) );
  NOR4X1_RVT U1301 ( .A1(a2stg_frac2a[26]), .A2(a2stg_frac2a[18]), .A3(
        a2stg_frac2a[5]), .A4(n740), .Y(n747) );
  NOR4X1_RVT U1302 ( .A1(a2stg_frac2a[27]), .A2(a2stg_frac2a[21]), .A3(
        a2stg_frac2a[13]), .A4(a2stg_frac2a[29]), .Y(n745) );
  NOR4X1_RVT U1303 ( .A1(a2stg_frac2a[7]), .A2(a2stg_frac2a[15]), .A3(
        a2stg_frac2a[31]), .A4(a2stg_frac2a[19]), .Y(n744) );
  AO222X1_RVT U1304 ( .A1(a2stg_shr_cnt[4]), .A2(a2stg_frac2a[42]), .A3(
        a2stg_shr_cnt[4]), .A4(a2stg_frac2a[41]), .A5(a2stg_shr_cnt[4]), .A6(
        a2stg_frac2a[43]), .Y(n741) );
  NOR4X1_RVT U1305 ( .A1(a2stg_frac2a[3]), .A2(a2stg_frac2a[2]), .A3(
        a2stg_frac2a[4]), .A4(n741), .Y(n743) );
  AND4X1_RVT U1306 ( .A1(n745), .A2(n744), .A3(n743), .A4(n742), .Y(n746) );
  NAND4X0_RVT U1307 ( .A1(n749), .A2(n748), .A3(n747), .A4(n746), .Y(n750) );
  AOI22X1_RVT U1308 ( .A1(a2stg_shr_cnt[4]), .A2(n751), .A3(a2stg_shr_cnt[5]), 
        .A4(n750), .Y(n2520) );
  AO21X1_RVT U1309 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[33]), .A3(
        a2stg_frac2a[1]), .Y(n812) );
  AO21X1_RVT U1310 ( .A1(a2stg_shr_cnt[4]), .A2(n752), .A3(n812), .Y(n826) );
  INVX1_RVT U1311 ( .A(a2stg_shr_cnt[4]), .Y(n820) );
  AO21X1_RVT U1312 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[35]), .A3(
        a2stg_frac2a[3]), .Y(n814) );
  NAND2X0_RVT U1313 ( .A1(a2stg_frac2a[34]), .A2(a2stg_shr_cnt[5]), .Y(n753)
         );
  NAND3X0_RVT U1314 ( .A1(n754), .A2(n820), .A3(n753), .Y(n819) );
  OAI22X1_RVT U1315 ( .A1(n821), .A2(n820), .A3(n814), .A4(n819), .Y(n757) );
  NAND2X0_RVT U1316 ( .A1(a2stg_shr_cnt[4]), .A2(n755), .Y(n756) );
  NAND3X0_RVT U1317 ( .A1(n758), .A2(n757), .A3(n756), .Y(n797) );
  AO21X1_RVT U1318 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[36]), .A3(
        a2stg_frac2a[4]), .Y(n811) );
  INVX1_RVT U1319 ( .A(n811), .Y(n761) );
  NAND2X0_RVT U1320 ( .A1(a2stg_shr_cnt[4]), .A2(n759), .Y(n760) );
  NAND2X0_RVT U1321 ( .A1(n761), .A2(n760), .Y(n798) );
  AO21X1_RVT U1322 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[38]), .A3(
        a2stg_frac2a[6]), .Y(n810) );
  INVX1_RVT U1323 ( .A(n810), .Y(n764) );
  NAND2X0_RVT U1324 ( .A1(a2stg_shr_cnt[4]), .A2(n762), .Y(n763) );
  NAND2X0_RVT U1325 ( .A1(n764), .A2(n763), .Y(n784) );
  AOI21X1_RVT U1326 ( .A1(a2stg_frac2a[39]), .A2(a2stg_shr_cnt[5]), .A3(
        a2stg_frac2a[7]), .Y(n818) );
  AO21X1_RVT U1327 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[32]), .A3(
        a2stg_frac2a[0]), .Y(n809) );
  OA22X1_RVT U1328 ( .A1(n820), .A2(n765), .A3(a2stg_shr_cnt[4]), .A4(n809), 
        .Y(n825) );
  INVX1_RVT U1329 ( .A(n825), .Y(n802) );
  AO21X1_RVT U1330 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[37]), .A3(
        a2stg_frac2a[5]), .Y(n808) );
  OAI22X1_RVT U1331 ( .A1(n820), .A2(n766), .A3(a2stg_shr_cnt[4]), .A4(n808), 
        .Y(n790) );
  NAND2X0_RVT U1332 ( .A1(a2stg_shr_cnt[4]), .A2(n767), .Y(n768) );
  NAND4X0_RVT U1333 ( .A1(n818), .A2(n802), .A3(n790), .A4(n768), .Y(n769) );
  NOR4X1_RVT U1334 ( .A1(n797), .A2(n798), .A3(n784), .A4(n769), .Y(n2521) );
  AO21X1_RVT U1335 ( .A1(a2stg_frac2a[40]), .A2(a2stg_shr_cnt[5]), .A3(
        a2stg_frac2a[8]), .Y(n807) );
  INVX1_RVT U1336 ( .A(n807), .Y(n772) );
  NAND2X0_RVT U1337 ( .A1(a2stg_shr_cnt[4]), .A2(n770), .Y(n771) );
  NAND2X0_RVT U1338 ( .A1(n772), .A2(n771), .Y(n2517) );
  INVX1_RVT U1339 ( .A(a2stg_shr_cnt[0]), .Y(n2503) );
  INVX1_RVT U1340 ( .A(a2stg_shr_cnt[1]), .Y(n788) );
  NAND2X0_RVT U1341 ( .A1(n2503), .A2(n788), .Y(n2504) );
  NAND2X0_RVT U1342 ( .A1(n2517), .A2(n2504), .Y(n781) );
  AO22X1_RVT U1343 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[41]), .A3(
        a2stg_shr_cnt[4]), .A4(n773), .Y(n774) );
  NOR2X0_RVT U1344 ( .A1(a2stg_frac2a[9]), .A2(n774), .Y(n2485) );
  NAND2X0_RVT U1345 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[42]), .Y(n775)
         );
  AND2X1_RVT U1346 ( .A1(n776), .A2(n775), .Y(n779) );
  NAND2X0_RVT U1347 ( .A1(a2stg_shr_cnt[4]), .A2(n777), .Y(n778) );
  AND2X1_RVT U1348 ( .A1(n779), .A2(n778), .Y(n2493) );
  AO221X1_RVT U1349 ( .A1(n2485), .A2(n2493), .A3(n2485), .A4(n2503), .A5(n788), .Y(n780) );
  NAND3X0_RVT U1350 ( .A1(n2521), .A2(n781), .A3(n780), .Y(n806) );
  AO22X1_RVT U1351 ( .A1(a2stg_shr_cnt[1]), .A2(n783), .A3(n782), .A4(n2504), 
        .Y(n804) );
  NAND2X0_RVT U1352 ( .A1(a2stg_shr_cnt[3]), .A2(n785), .Y(n786) );
  NAND2X0_RVT U1353 ( .A1(n787), .A2(n786), .Y(n2515) );
  AO221X1_RVT U1354 ( .A1(n790), .A2(n789), .A3(n790), .A4(n2503), .A5(n788), 
        .Y(n801) );
  NAND3X0_RVT U1355 ( .A1(a2stg_shr_cnt[3]), .A2(n2493), .A3(n2485), .Y(n796)
         );
  NAND2X0_RVT U1356 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[43]), .Y(n791)
         );
  AND2X1_RVT U1357 ( .A1(n792), .A2(n791), .Y(n795) );
  NAND2X0_RVT U1358 ( .A1(a2stg_shr_cnt[4]), .A2(n793), .Y(n794) );
  NAND2X0_RVT U1359 ( .A1(n795), .A2(n794), .Y(n2490) );
  OA22X1_RVT U1360 ( .A1(a2stg_shr_cnt[3]), .A2(n797), .A3(n796), .A4(n2490), 
        .Y(n2518) );
  NAND2X0_RVT U1361 ( .A1(n2504), .A2(n798), .Y(n799) );
  NAND4X0_RVT U1362 ( .A1(n802), .A2(n801), .A3(n800), .A4(n799), .Y(n803) );
  AO221X1_RVT U1363 ( .A1(a2stg_shr_cnt[3]), .A2(n2517), .A3(a2stg_shr_cnt[3]), 
        .A4(n804), .A5(n803), .Y(n805) );
  AOI22X1_RVT U1364 ( .A1(a2stg_shr_cnt[3]), .A2(n806), .A3(a2stg_shr_cnt[2]), 
        .A4(n805), .Y(n831) );
  NOR4X1_RVT U1365 ( .A1(n810), .A2(n809), .A3(n808), .A4(n807), .Y(n816) );
  AO21X1_RVT U1366 ( .A1(a2stg_shr_cnt[5]), .A2(a2stg_frac2a[34]), .A3(
        a2stg_frac2a[2]), .Y(n813) );
  NOR4X1_RVT U1367 ( .A1(n814), .A2(n813), .A3(n812), .A4(n811), .Y(n815) );
  NAND2X0_RVT U1368 ( .A1(n816), .A2(n815), .Y(n2516) );
  AO21X1_RVT U1369 ( .A1(n818), .A2(n817), .A3(n820), .Y(n830) );
  AND2X1_RVT U1370 ( .A1(n819), .A2(a2stg_shr_cnt[0]), .Y(n824) );
  NAND2X0_RVT U1371 ( .A1(a2stg_shr_cnt[4]), .A2(n822), .Y(n823) );
  AND2X1_RVT U1372 ( .A1(n824), .A2(n823), .Y(n827) );
  AO221X1_RVT U1373 ( .A1(a2stg_shr_cnt[1]), .A2(n827), .A3(a2stg_shr_cnt[1]), 
        .A4(n826), .A5(n825), .Y(n828) );
  NAND2X0_RVT U1374 ( .A1(n2504), .A2(n828), .Y(n829) );
  NAND4X0_RVT U1375 ( .A1(n2520), .A2(n831), .A3(n830), .A4(n829), .Y(
        a2stg_fsdtoix_nx) );
  AND2X1_RVT U1376 ( .A1(n1813), .A2(n1800), .Y(n1820) );
  AO22X1_RVT U1377 ( .A1(a4stg_shl_cnt_dec54_1[0]), .A2(a4stg_shl_data[47]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[63]), .Y(n840) );
  AO22X1_RVT U1378 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[31]), 
        .A3(\a4stg_shl_cnt_dec54_3[0] ), .A4(a4stg_shl_data[15]), .Y(n839) );
  AO22X1_RVT U1379 ( .A1(a4stg_shl_cnt_dec54_1[0]), .A2(a4stg_shl_data[46]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[62]), .Y(n833) );
  AO22X1_RVT U1380 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[30]), 
        .A3(\a4stg_shl_cnt_dec54_3[0] ), .A4(a4stg_shl_data[14]), .Y(n832) );
  OR2X1_RVT U1381 ( .A1(n833), .A2(n832), .Y(n1391) );
  AO22X1_RVT U1382 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[12]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[44]), .Y(n835) );
  AO22X1_RVT U1383 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[28]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[60]), .Y(n834) );
  OR2X1_RVT U1384 ( .A1(n835), .A2(n834), .Y(n1387) );
  AO22X1_RVT U1385 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[29]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[45]), .Y(n837) );
  AO22X1_RVT U1386 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[13]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[61]), .Y(n836) );
  OR2X1_RVT U1387 ( .A1(n837), .A2(n836), .Y(n1390) );
  AO22X1_RVT U1388 ( .A1(a4stg_shl_cnt[0]), .A2(n1387), .A3(n1800), .A4(n1390), 
        .Y(n1408) );
  OA222X1_RVT U1389 ( .A1(a4stg_shl_cnt[1]), .A2(a4stg_shl_cnt[0]), .A3(
        a4stg_shl_cnt[1]), .A4(n1391), .A5(n1408), .A6(n1813), .Y(n838) );
  AO221X1_RVT U1390 ( .A1(n1820), .A2(n840), .A3(n1820), .A4(n839), .A5(n838), 
        .Y(n865) );
  AO22X1_RVT U1391 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[8]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[40]), .Y(n842) );
  AO22X1_RVT U1392 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[24]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[56]), .Y(n841) );
  OR2X1_RVT U1393 ( .A1(n842), .A2(n841), .Y(n1392) );
  AO22X1_RVT U1394 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[25]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[41]), .Y(n844) );
  AO22X1_RVT U1395 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[9]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[57]), .Y(n843) );
  OR2X1_RVT U1396 ( .A1(n844), .A2(n843), .Y(n1395) );
  AO22X1_RVT U1397 ( .A1(a4stg_shl_cnt[0]), .A2(n1392), .A3(n1800), .A4(n1395), 
        .Y(n1413) );
  AO22X1_RVT U1398 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[26]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[58]), .Y(n846) );
  AO22X1_RVT U1399 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[10]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[42]), .Y(n845) );
  OR2X1_RVT U1400 ( .A1(n846), .A2(n845), .Y(n1394) );
  AO22X1_RVT U1401 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[11]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[43]), .Y(n848) );
  AO22X1_RVT U1402 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[27]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[59]), .Y(n847) );
  OR2X1_RVT U1403 ( .A1(n848), .A2(n847), .Y(n1388) );
  AO22X1_RVT U1404 ( .A1(a4stg_shl_cnt[0]), .A2(n1394), .A3(n1800), .A4(n1388), 
        .Y(n1407) );
  AO22X1_RVT U1405 ( .A1(a4stg_shl_cnt[1]), .A2(n1413), .A3(n1813), .A4(n1407), 
        .Y(n1435) );
  INVX1_RVT U1406 ( .A(a4stg_shl_cnt[3]), .Y(n1546) );
  AND2X1_RVT U1407 ( .A1(a4stg_shl_cnt[2]), .A2(n1546), .Y(n1459) );
  AO22X1_RVT U1408 ( .A1(a4stg_shl_data[32]), .A2(a4stg_shl_cnt_dec54_1[0]), 
        .A3(a4stg_shl_data[48]), .A4(a4stg_shl_cnt_dec54_0[0]), .Y(n850) );
  AO22X1_RVT U1409 ( .A1(a4stg_shl_data[16]), .A2(\a4stg_shl_cnt_dec54_2[0] ), 
        .A3(a4stg_shl_data[0]), .A4(\a4stg_shl_cnt_dec54_3[0] ), .Y(n849) );
  OR2X1_RVT U1410 ( .A1(n850), .A2(n849), .Y(n1396) );
  AO22X1_RVT U1411 ( .A1(a4stg_shl_cnt_dec54_1[0]), .A2(a4stg_shl_data[33]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[49]), .Y(n852) );
  AO22X1_RVT U1412 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[17]), 
        .A3(\a4stg_shl_cnt_dec54_3[0] ), .A4(a4stg_shl_data[1]), .Y(n851) );
  OR2X1_RVT U1413 ( .A1(n852), .A2(n851), .Y(n1398) );
  AO22X1_RVT U1414 ( .A1(a4stg_shl_cnt[0]), .A2(n1396), .A3(n1800), .A4(n1398), 
        .Y(n1410) );
  AO22X1_RVT U1415 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[2]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[34]), .Y(n854) );
  AO22X1_RVT U1416 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[18]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[50]), .Y(n853) );
  OR2X1_RVT U1417 ( .A1(n854), .A2(n853), .Y(n1397) );
  AO22X1_RVT U1418 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[3]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[35]), .Y(n856) );
  AO22X1_RVT U1419 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[19]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[51]), .Y(n855) );
  OR2X1_RVT U1420 ( .A1(n856), .A2(n855), .Y(n1400) );
  AO22X1_RVT U1421 ( .A1(a4stg_shl_cnt[0]), .A2(n1397), .A3(n1800), .A4(n1400), 
        .Y(n1412) );
  AO22X1_RVT U1422 ( .A1(a4stg_shl_cnt[1]), .A2(n1410), .A3(n1813), .A4(n1412), 
        .Y(n1434) );
  INVX1_RVT U1423 ( .A(a4stg_shl_cnt[2]), .Y(n1826) );
  AO22X1_RVT U1424 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[4]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[52]), .Y(n858) );
  AO22X1_RVT U1425 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[20]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[36]), .Y(n857) );
  OR2X1_RVT U1426 ( .A1(n858), .A2(n857), .Y(n1399) );
  AO22X1_RVT U1427 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[21]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[37]), .Y(n860) );
  AO22X1_RVT U1428 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[5]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[53]), .Y(n859) );
  OR2X1_RVT U1429 ( .A1(n860), .A2(n859), .Y(n1402) );
  AO22X1_RVT U1430 ( .A1(a4stg_shl_cnt[0]), .A2(n1399), .A3(n1800), .A4(n1402), 
        .Y(n1411) );
  AO22X1_RVT U1431 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[22]), 
        .A3(a4stg_shl_cnt_dec54_1[0]), .A4(a4stg_shl_data[38]), .Y(n862) );
  AO22X1_RVT U1432 ( .A1(\a4stg_shl_cnt_dec54_3[0] ), .A2(a4stg_shl_data[6]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[54]), .Y(n861) );
  OR2X1_RVT U1433 ( .A1(n862), .A2(n861), .Y(n1401) );
  AO22X1_RVT U1434 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[23]), 
        .A3(\a4stg_shl_cnt_dec54_3[0] ), .A4(a4stg_shl_data[7]), .Y(n864) );
  AO22X1_RVT U1435 ( .A1(a4stg_shl_cnt_dec54_1[0]), .A2(a4stg_shl_data[39]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[55]), .Y(n863) );
  OR2X1_RVT U1436 ( .A1(n864), .A2(n863), .Y(n1393) );
  AO22X1_RVT U1437 ( .A1(a4stg_shl_cnt[0]), .A2(n1401), .A3(n1800), .A4(n1393), 
        .Y(n1414) );
  AO22X1_RVT U1438 ( .A1(a4stg_shl_cnt[1]), .A2(n1411), .A3(n1813), .A4(n1414), 
        .Y(n1436) );
  AO22X1_RVT U1439 ( .A1(a4stg_shl_cnt[2]), .A2(n1434), .A3(n1826), .A4(n1436), 
        .Y(n1468) );
  AO222X1_RVT U1440 ( .A1(n865), .A2(n1874), .A3(n1435), .A4(n1459), .A5(n1468), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[63]) );
  OAI22X1_RVT U1441 ( .A1(a4stg_rnd_frac_add_inv), .A2(n2526), .A3(
        a3stg_inc_exp_inv), .A4(n866), .Y(n1877) );
  NOR2X0_RVT U1442 ( .A1(a4stg_fixtos_fxtod_inv), .A2(n2526), .Y(n1875) );
  AO22X1_RVT U1443 ( .A1(n1920), .A2(n1877), .A3(n1875), .A4(a4stg_shl[63]), 
        .Y(n868) );
  NOR2X0_RVT U1444 ( .A1(a3stg_fdtos_inv), .A2(n2526), .Y(n1870) );
  AO22X1_RVT U1445 ( .A1(n1870), .A2(n1404), .A3(n2526), .A4(a4stg_rnd_frac_63), .Y(n867) );
  OR2X1_RVT U1446 ( .A1(n868), .A2(n867), .Y(a4stg_rnd_frac_pre2_in[63]) );
  INVX1_RVT U1447 ( .A(a1stg_in2[53]), .Y(n871) );
  AOI222X1_RVT U1448 ( .A1(n870), .A2(a1stg_in1[54]), .A3(a1stg_in2[54]), .A4(
        n869), .A5(n871), .A6(a1stg_in1[53]), .Y(n892) );
  OA222X1_RVT U1449 ( .A1(a1stg_in2[52]), .A2(n873), .A3(n872), .A4(
        a1stg_in1[52]), .A5(a1stg_in1[53]), .A6(n871), .Y(n891) );
  INVX1_RVT U1450 ( .A(a1stg_in2[62]), .Y(n876) );
  INVX1_RVT U1451 ( .A(a1stg_in2[57]), .Y(n875) );
  AOI22X1_RVT U1452 ( .A1(n875), .A2(a1stg_in1[57]), .A3(n876), .A4(
        a1stg_in1[62]), .Y(n874) );
  OA221X1_RVT U1453 ( .A1(n876), .A2(a1stg_in1[62]), .A3(n875), .A4(
        a1stg_in1[57]), .A5(n874), .Y(n889) );
  INVX1_RVT U1454 ( .A(a1stg_in2[59]), .Y(n879) );
  INVX1_RVT U1455 ( .A(a1stg_in2[55]), .Y(n878) );
  AOI22X1_RVT U1456 ( .A1(n879), .A2(a1stg_in1[59]), .A3(n878), .A4(
        a1stg_in1[55]), .Y(n877) );
  OA221X1_RVT U1457 ( .A1(n879), .A2(a1stg_in1[59]), .A3(n878), .A4(
        a1stg_in1[55]), .A5(n877), .Y(n888) );
  INVX1_RVT U1458 ( .A(a1stg_in2[61]), .Y(n882) );
  INVX1_RVT U1459 ( .A(a1stg_in2[56]), .Y(n881) );
  AOI22X1_RVT U1460 ( .A1(n882), .A2(a1stg_in1[61]), .A3(n881), .A4(
        a1stg_in1[56]), .Y(n880) );
  OA221X1_RVT U1461 ( .A1(n882), .A2(a1stg_in1[61]), .A3(n881), .A4(
        a1stg_in1[56]), .A5(n880), .Y(n887) );
  INVX1_RVT U1462 ( .A(a1stg_in2[60]), .Y(n885) );
  INVX1_RVT U1463 ( .A(a1stg_in2[58]), .Y(n884) );
  AOI22X1_RVT U1464 ( .A1(n884), .A2(a1stg_in1[58]), .A3(n885), .A4(
        a1stg_in1[60]), .Y(n883) );
  OA221X1_RVT U1465 ( .A1(n885), .A2(a1stg_in1[60]), .A3(n884), .A4(
        a1stg_in1[58]), .A5(n883), .Y(n886) );
  AND4X1_RVT U1466 ( .A1(n889), .A2(n888), .A3(n887), .A4(n886), .Y(n890) );
  OA221X1_RVT U1467 ( .A1(a1stg_sngop), .A2(n892), .A3(a1stg_sngop), .A4(n891), 
        .A5(n890), .Y(a1stg_in2_eq_in1_exp) );
  AOI22X1_RVT U1468 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[54]), .A3(
        a1stg_in2[51]), .A4(a1stg_denorm_dbl_in2), .Y(n896) );
  NAND2X0_RVT U1469 ( .A1(a1stg_intlngop), .A2(a1stg_in2[63]), .Y(n893) );
  NAND4X0_RVT U1470 ( .A1(n896), .A2(n895), .A3(n894), .A4(n893), .Y(n1033) );
  AO22X1_RVT U1471 ( .A1(a1stg_in1[54]), .A2(a1stg_denorm_sng_in1), .A3(
        a1stg_in1[51]), .A4(a1stg_denorm_dbl_in1), .Y(n897) );
  AO22X1_RVT U1472 ( .A1(n1030), .A2(n1033), .A3(n1024), .A4(n1034), .Y(
        a2stg_frac1_in[63]) );
  AOI22X1_RVT U1473 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[54]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[62]), .Y(n900) );
  AOI22X1_RVT U1474 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[51]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[50]), .Y(n899) );
  NAND2X0_RVT U1475 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[53]), .Y(n898)
         );
  NAND3X0_RVT U1476 ( .A1(n900), .A2(n899), .A3(n898), .Y(n1035) );
  AO22X1_RVT U1477 ( .A1(a1stg_denorm_dbl_in1), .A2(a1stg_in1[50]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[53]), .Y(n902) );
  AO22X1_RVT U1478 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[54]), .A3(
        a1stg_norm_dbl_in1), .A4(a1stg_in1[51]), .Y(n901) );
  OR2X1_RVT U1479 ( .A1(n902), .A2(n901), .Y(n1037) );
  AO222X1_RVT U1480 ( .A1(n1035), .A2(n1030), .A3(n907), .A4(
        a2stg_frac1_in_qnan), .A5(n1024), .A6(n1037), .Y(a2stg_frac1_in[62])
         );
  AOI22X1_RVT U1481 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[52]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[50]), .Y(n904) );
  NAND2X0_RVT U1482 ( .A1(a1stg_in2[53]), .A2(a1stg_norm_sng_in2), .Y(n903) );
  NAND3X0_RVT U1483 ( .A1(n26), .A2(n904), .A3(n903), .Y(n1038) );
  AO22X1_RVT U1484 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[53]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[52]), .Y(n906) );
  AO22X1_RVT U1485 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[50]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[49]), .Y(n905) );
  OR2X1_RVT U1486 ( .A1(n906), .A2(n905), .Y(n1039) );
  AOI22X1_RVT U1487 ( .A1(n1030), .A2(n1038), .A3(n1024), .A4(n1039), .Y(n908)
         );
  NAND2X0_RVT U1488 ( .A1(a2stg_frac1_in_nv), .A2(n907), .Y(n1025) );
  NAND2X0_RVT U1489 ( .A1(n908), .A2(n1025), .Y(a2stg_frac1_in[61]) );
  AOI22X1_RVT U1490 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[51]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[49]), .Y(n910) );
  NAND2X0_RVT U1491 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[52]), .Y(n909) );
  NAND3X0_RVT U1492 ( .A1(n910), .A2(n28), .A3(n909), .Y(n1040) );
  AO22X1_RVT U1493 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[52]), .A3(
        a1stg_in1[51]), .A4(a1stg_denorm_sng_in1), .Y(n912) );
  AO22X1_RVT U1494 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[49]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[48]), .Y(n911) );
  OR2X1_RVT U1495 ( .A1(n912), .A2(n911), .Y(n1041) );
  AOI22X1_RVT U1496 ( .A1(n1030), .A2(n1040), .A3(n1024), .A4(n1041), .Y(n913)
         );
  NAND2X0_RVT U1497 ( .A1(n913), .A2(n1025), .Y(a2stg_frac1_in[60]) );
  AOI22X1_RVT U1498 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[50]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[59]), .Y(n915) );
  NAND2X0_RVT U1499 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[51]), .Y(n914) );
  NAND3X0_RVT U1500 ( .A1(n915), .A2(n29), .A3(n914), .Y(n1042) );
  AO22X1_RVT U1501 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[51]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[47]), .Y(n917) );
  AO22X1_RVT U1502 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[48]), .A3(
        a1stg_in1[50]), .A4(a1stg_denorm_sng_in1), .Y(n916) );
  OR2X1_RVT U1503 ( .A1(n917), .A2(n916), .Y(n1043) );
  AOI22X1_RVT U1504 ( .A1(n1030), .A2(n1042), .A3(n1024), .A4(n1043), .Y(n918)
         );
  NAND2X0_RVT U1505 ( .A1(n918), .A2(n1025), .Y(a2stg_frac1_in[59]) );
  AOI22X1_RVT U1506 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[49]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[58]), .Y(n920) );
  NAND2X0_RVT U1507 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[50]), .Y(n919) );
  NAND3X0_RVT U1508 ( .A1(n27), .A2(n920), .A3(n919), .Y(n1044) );
  AO22X1_RVT U1509 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[47]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[49]), .Y(n922) );
  AO22X1_RVT U1510 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[50]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[46]), .Y(n921) );
  OR2X1_RVT U1511 ( .A1(n922), .A2(n921), .Y(n1045) );
  AOI22X1_RVT U1512 ( .A1(n1030), .A2(n1044), .A3(n1024), .A4(n1045), .Y(n923)
         );
  NAND2X0_RVT U1513 ( .A1(n923), .A2(n1025), .Y(a2stg_frac1_in[58]) );
  AOI22X1_RVT U1514 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[48]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[57]), .Y(n925) );
  NAND2X0_RVT U1515 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[49]), .Y(n924) );
  NAND3X0_RVT U1516 ( .A1(n925), .A2(n30), .A3(n924), .Y(n1046) );
  AO22X1_RVT U1517 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[46]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[48]), .Y(n927) );
  AO22X1_RVT U1518 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[49]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[45]), .Y(n926) );
  OR2X1_RVT U1519 ( .A1(n927), .A2(n926), .Y(n1047) );
  AOI22X1_RVT U1520 ( .A1(n1030), .A2(n1046), .A3(n1024), .A4(n1047), .Y(n928)
         );
  NAND2X0_RVT U1521 ( .A1(n928), .A2(n1025), .Y(a2stg_frac1_in[57]) );
  AOI22X1_RVT U1522 ( .A1(a1stg_intlngop), .A2(a1stg_in2[56]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[45]), .Y(n931) );
  AOI22X1_RVT U1523 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[47]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[44]), .Y(n930) );
  NAND2X0_RVT U1524 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[48]), .Y(n929) );
  NAND3X0_RVT U1525 ( .A1(n931), .A2(n930), .A3(n929), .Y(n1048) );
  AO22X1_RVT U1526 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[45]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[47]), .Y(n933) );
  AO22X1_RVT U1527 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[48]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[44]), .Y(n932) );
  OR2X1_RVT U1528 ( .A1(n933), .A2(n932), .Y(n1049) );
  AOI22X1_RVT U1529 ( .A1(n1030), .A2(n1048), .A3(n1024), .A4(n1049), .Y(n934)
         );
  NAND2X0_RVT U1530 ( .A1(n934), .A2(n1025), .Y(a2stg_frac1_in[56]) );
  AOI22X1_RVT U1531 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[47]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[55]), .Y(n936) );
  NAND2X0_RVT U1532 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[46]), .Y(n935)
         );
  NAND3X0_RVT U1533 ( .A1(n936), .A2(n31), .A3(n935), .Y(n1050) );
  AO22X1_RVT U1534 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[47]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[43]), .Y(n938) );
  AO22X1_RVT U1535 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[44]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[46]), .Y(n937) );
  OR2X1_RVT U1536 ( .A1(n938), .A2(n937), .Y(n1051) );
  AOI22X1_RVT U1537 ( .A1(n1030), .A2(n1050), .A3(n1024), .A4(n1051), .Y(n939)
         );
  NAND2X0_RVT U1538 ( .A1(n939), .A2(n1025), .Y(a2stg_frac1_in[55]) );
  AOI22X1_RVT U1539 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[43]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[42]), .Y(n941) );
  NAND2X0_RVT U1540 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[45]), .Y(n940)
         );
  NAND3X0_RVT U1541 ( .A1(n941), .A2(n6), .A3(n940), .Y(n1052) );
  AO22X1_RVT U1542 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[43]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[45]), .Y(n943) );
  AO22X1_RVT U1543 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[46]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[42]), .Y(n942) );
  OR2X1_RVT U1544 ( .A1(n943), .A2(n942), .Y(n1053) );
  AOI22X1_RVT U1545 ( .A1(n1030), .A2(n1052), .A3(n1024), .A4(n1053), .Y(n944)
         );
  NAND2X0_RVT U1546 ( .A1(n944), .A2(n1025), .Y(a2stg_frac1_in[54]) );
  AOI22X1_RVT U1547 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[44]), .A3(
        a1stg_in2[53]), .A4(a1stg_intlngop), .Y(n947) );
  AOI22X1_RVT U1548 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[42]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[41]), .Y(n946) );
  NAND2X0_RVT U1549 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[45]), .Y(n945) );
  NAND3X0_RVT U1550 ( .A1(n947), .A2(n946), .A3(n945), .Y(n1054) );
  AO22X1_RVT U1551 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[45]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[44]), .Y(n949) );
  AO22X1_RVT U1552 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[42]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[41]), .Y(n948) );
  OR2X1_RVT U1553 ( .A1(n949), .A2(n948), .Y(n1055) );
  AOI22X1_RVT U1554 ( .A1(n1030), .A2(n1054), .A3(n1024), .A4(n1055), .Y(n950)
         );
  NAND2X0_RVT U1555 ( .A1(n950), .A2(n1025), .Y(a2stg_frac1_in[53]) );
  AOI22X1_RVT U1556 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[43]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[41]), .Y(n952) );
  NAND2X0_RVT U1557 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[44]), .Y(n951) );
  NAND3X0_RVT U1558 ( .A1(n952), .A2(n32), .A3(n951), .Y(n1056) );
  AO22X1_RVT U1559 ( .A1(a1stg_denorm_dbl_in1), .A2(a1stg_in1[40]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[43]), .Y(n954) );
  AO22X1_RVT U1560 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[44]), .A3(
        a1stg_norm_dbl_in1), .A4(a1stg_in1[41]), .Y(n953) );
  OR2X1_RVT U1561 ( .A1(n954), .A2(n953), .Y(n1057) );
  AOI22X1_RVT U1562 ( .A1(n1030), .A2(n1056), .A3(n1024), .A4(n1057), .Y(n955)
         );
  NAND2X0_RVT U1563 ( .A1(n955), .A2(n1025), .Y(a2stg_frac1_in[52]) );
  AOI22X1_RVT U1564 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[42]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[51]), .Y(n958) );
  AOI22X1_RVT U1565 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[40]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[39]), .Y(n957) );
  NAND2X0_RVT U1566 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[43]), .Y(n956) );
  NAND3X0_RVT U1567 ( .A1(n958), .A2(n957), .A3(n956), .Y(n1058) );
  AO22X1_RVT U1568 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[43]), .A3(
        a1stg_norm_dbl_in1), .A4(a1stg_in1[40]), .Y(n960) );
  AO22X1_RVT U1569 ( .A1(a1stg_denorm_dbl_in1), .A2(a1stg_in1[39]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[42]), .Y(n959) );
  OR2X1_RVT U1570 ( .A1(n960), .A2(n959), .Y(n1059) );
  AOI22X1_RVT U1571 ( .A1(n1030), .A2(n1058), .A3(n1024), .A4(n1059), .Y(n961)
         );
  NAND2X0_RVT U1572 ( .A1(n961), .A2(n1025), .Y(a2stg_frac1_in[51]) );
  AOI22X1_RVT U1573 ( .A1(a1stg_intlngop), .A2(a1stg_in2[50]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[38]), .Y(n964) );
  AOI22X1_RVT U1574 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[42]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[39]), .Y(n963) );
  NAND2X0_RVT U1575 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[41]), .Y(n962)
         );
  NAND3X0_RVT U1576 ( .A1(n964), .A2(n963), .A3(n962), .Y(n1060) );
  AO22X1_RVT U1577 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[42]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[38]), .Y(n966) );
  AO22X1_RVT U1578 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[39]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[41]), .Y(n965) );
  OR2X1_RVT U1579 ( .A1(n966), .A2(n965), .Y(n1061) );
  AOI22X1_RVT U1580 ( .A1(n1030), .A2(n1060), .A3(n1024), .A4(n1061), .Y(n967)
         );
  NAND2X0_RVT U1581 ( .A1(n967), .A2(n1025), .Y(a2stg_frac1_in[50]) );
  AOI22X1_RVT U1582 ( .A1(a1stg_intlngop), .A2(a1stg_in2[49]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[37]), .Y(n970) );
  AOI22X1_RVT U1583 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[41]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[38]), .Y(n969) );
  NAND2X0_RVT U1584 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[40]), .Y(n968)
         );
  NAND3X0_RVT U1585 ( .A1(n970), .A2(n969), .A3(n968), .Y(n1062) );
  AO22X1_RVT U1586 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[41]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[40]), .Y(n972) );
  AO22X1_RVT U1587 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[38]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[37]), .Y(n971) );
  OR2X1_RVT U1588 ( .A1(n972), .A2(n971), .Y(n1063) );
  AOI22X1_RVT U1589 ( .A1(n1030), .A2(n1062), .A3(n1024), .A4(n1063), .Y(n973)
         );
  NAND2X0_RVT U1590 ( .A1(n973), .A2(n1025), .Y(a2stg_frac1_in[49]) );
  AOI22X1_RVT U1591 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[39]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[48]), .Y(n976) );
  AOI22X1_RVT U1592 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[40]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[37]), .Y(n975) );
  NAND2X0_RVT U1593 ( .A1(a1stg_denorm_dbl_in2), .A2(a1stg_in2[36]), .Y(n974)
         );
  NAND3X0_RVT U1594 ( .A1(n976), .A2(n975), .A3(n974), .Y(n1064) );
  AO22X1_RVT U1595 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[40]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[36]), .Y(n978) );
  AO22X1_RVT U1596 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[37]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[39]), .Y(n977) );
  OR2X1_RVT U1597 ( .A1(n978), .A2(n977), .Y(n1065) );
  AOI22X1_RVT U1598 ( .A1(n1030), .A2(n1064), .A3(n1024), .A4(n1065), .Y(n979)
         );
  NAND2X0_RVT U1599 ( .A1(n979), .A2(n1025), .Y(a2stg_frac1_in[48]) );
  AOI22X1_RVT U1600 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[38]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[47]), .Y(n982) );
  AOI22X1_RVT U1601 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[39]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[36]), .Y(n981) );
  NAND2X0_RVT U1602 ( .A1(a1stg_denorm_dbl_in2), .A2(a1stg_in2[35]), .Y(n980)
         );
  NAND3X0_RVT U1603 ( .A1(n982), .A2(n981), .A3(n980), .Y(n1066) );
  AO22X1_RVT U1604 ( .A1(a1stg_denorm_dbl_in1), .A2(a1stg_in1[35]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[38]), .Y(n984) );
  AO22X1_RVT U1605 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[39]), .A3(
        a1stg_norm_dbl_in1), .A4(a1stg_in1[36]), .Y(n983) );
  OR2X1_RVT U1606 ( .A1(n984), .A2(n983), .Y(n1067) );
  AOI22X1_RVT U1607 ( .A1(n1030), .A2(n1066), .A3(n1024), .A4(n1067), .Y(n985)
         );
  NAND2X0_RVT U1608 ( .A1(n985), .A2(n1025), .Y(a2stg_frac1_in[47]) );
  AOI22X1_RVT U1609 ( .A1(a1stg_intlngop), .A2(a1stg_in2[46]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[34]), .Y(n988) );
  AOI22X1_RVT U1610 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[37]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[35]), .Y(n987) );
  NAND2X0_RVT U1611 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[38]), .Y(n986) );
  NAND3X0_RVT U1612 ( .A1(n988), .A2(n987), .A3(n986), .Y(n1068) );
  AO22X1_RVT U1613 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[38]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[34]), .Y(n990) );
  AO22X1_RVT U1614 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[35]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[37]), .Y(n989) );
  OR2X1_RVT U1615 ( .A1(n990), .A2(n989), .Y(n1069) );
  AOI22X1_RVT U1616 ( .A1(n1030), .A2(n1068), .A3(n1024), .A4(n1069), .Y(n991)
         );
  NAND2X0_RVT U1617 ( .A1(n991), .A2(n1025), .Y(a2stg_frac1_in[46]) );
  AOI22X1_RVT U1618 ( .A1(a1stg_intlngop), .A2(a1stg_in2[45]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[33]), .Y(n994) );
  AOI22X1_RVT U1619 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[36]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[34]), .Y(n993) );
  NAND2X0_RVT U1620 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[37]), .Y(n992) );
  NAND3X0_RVT U1621 ( .A1(n994), .A2(n993), .A3(n992), .Y(n1070) );
  AO22X1_RVT U1622 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[37]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[33]), .Y(n996) );
  AO22X1_RVT U1623 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[34]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[36]), .Y(n995) );
  OR2X1_RVT U1624 ( .A1(n996), .A2(n995), .Y(n1071) );
  AOI22X1_RVT U1625 ( .A1(n1030), .A2(n1070), .A3(n1024), .A4(n1071), .Y(n997)
         );
  NAND2X0_RVT U1626 ( .A1(n997), .A2(n1025), .Y(a2stg_frac1_in[45]) );
  AOI22X1_RVT U1627 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[35]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[44]), .Y(n1000) );
  AOI22X1_RVT U1628 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[33]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[32]), .Y(n999) );
  NAND2X0_RVT U1629 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[36]), .Y(n998) );
  NAND3X0_RVT U1630 ( .A1(n1000), .A2(n999), .A3(n998), .Y(n1072) );
  AO22X1_RVT U1631 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[36]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[35]), .Y(n1002) );
  AO22X1_RVT U1632 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[33]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[32]), .Y(n1001) );
  OR2X1_RVT U1633 ( .A1(n1002), .A2(n1001), .Y(n1073) );
  AOI22X1_RVT U1634 ( .A1(n1030), .A2(n1072), .A3(n1024), .A4(n1073), .Y(n1003) );
  NAND2X0_RVT U1635 ( .A1(n1003), .A2(n1025), .Y(a2stg_frac1_in[44]) );
  AOI22X1_RVT U1636 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[34]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[43]), .Y(n1006) );
  AOI22X1_RVT U1637 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[35]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[32]), .Y(n1005) );
  NAND2X0_RVT U1638 ( .A1(a1stg_denorm_dbl_in2), .A2(a1stg_in2[31]), .Y(n1004)
         );
  NAND3X0_RVT U1639 ( .A1(n1006), .A2(n1005), .A3(n1004), .Y(n1074) );
  AO22X1_RVT U1640 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[35]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[31]), .Y(n1008) );
  AO22X1_RVT U1641 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[32]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[34]), .Y(n1007) );
  OR2X1_RVT U1642 ( .A1(n1008), .A2(n1007), .Y(n1075) );
  AOI22X1_RVT U1643 ( .A1(n1030), .A2(n1074), .A3(n1024), .A4(n1075), .Y(n1009) );
  NAND2X0_RVT U1644 ( .A1(n1009), .A2(n1025), .Y(a2stg_frac1_in[43]) );
  AOI22X1_RVT U1645 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[33]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[42]), .Y(n1012) );
  AOI22X1_RVT U1646 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[34]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[31]), .Y(n1011) );
  NAND2X0_RVT U1647 ( .A1(a1stg_denorm_dbl_in2), .A2(a1stg_in2[30]), .Y(n1010)
         );
  NAND3X0_RVT U1648 ( .A1(n1012), .A2(n1011), .A3(n1010), .Y(n1076) );
  AO22X1_RVT U1649 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[34]), .A3(
        a1stg_norm_dbl_in1), .A4(a1stg_in1[31]), .Y(n1014) );
  AO22X1_RVT U1650 ( .A1(a1stg_denorm_dbl_in1), .A2(a1stg_in1[30]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[33]), .Y(n1013) );
  OR2X1_RVT U1651 ( .A1(n1014), .A2(n1013), .Y(n1077) );
  AOI22X1_RVT U1652 ( .A1(n1030), .A2(n1076), .A3(n1024), .A4(n1077), .Y(n1015) );
  NAND2X0_RVT U1653 ( .A1(n1015), .A2(n1025), .Y(a2stg_frac1_in[42]) );
  AOI22X1_RVT U1654 ( .A1(a1stg_intlngop), .A2(a1stg_in2[41]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[29]), .Y(n1018) );
  AOI22X1_RVT U1655 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[33]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[30]), .Y(n1017) );
  NAND2X0_RVT U1656 ( .A1(a1stg_denorm_sng_in2), .A2(a1stg_in2[32]), .Y(n1016)
         );
  NAND3X0_RVT U1657 ( .A1(n1018), .A2(n1017), .A3(n1016), .Y(n1078) );
  AO22X1_RVT U1658 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[33]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[29]), .Y(n1020) );
  AO22X1_RVT U1659 ( .A1(a1stg_norm_dbl_in1), .A2(a1stg_in1[30]), .A3(
        a1stg_denorm_sng_in1), .A4(a1stg_in1[32]), .Y(n1019) );
  OR2X1_RVT U1660 ( .A1(n1020), .A2(n1019), .Y(n1079) );
  AOI22X1_RVT U1661 ( .A1(n1030), .A2(n1078), .A3(n1024), .A4(n1079), .Y(n1021) );
  NAND2X0_RVT U1662 ( .A1(n1021), .A2(n1025), .Y(a2stg_frac1_in[41]) );
  AO22X1_RVT U1663 ( .A1(a1stg_norm_dbl_in2), .A2(a1stg_in2[29]), .A3(
        a1stg_denorm_dbl_in2), .A4(a1stg_in2[28]), .Y(n1023) );
  AO22X1_RVT U1664 ( .A1(a1stg_norm_sng_in2), .A2(a1stg_in2[32]), .A3(
        a1stg_intlngop), .A4(a1stg_in2[40]), .Y(n1022) );
  OR2X1_RVT U1665 ( .A1(n1023), .A2(n1022), .Y(n1080) );
  AO222X1_RVT U1666 ( .A1(a1stg_norm_sng_in1), .A2(a1stg_in1[32]), .A3(
        a1stg_denorm_dbl_in1), .A4(a1stg_in1[28]), .A5(a1stg_in1[29]), .A6(
        a1stg_norm_dbl_in1), .Y(n1081) );
  AOI22X1_RVT U1667 ( .A1(n1030), .A2(n1080), .A3(n1024), .A4(n1081), .Y(n1026) );
  NAND2X0_RVT U1668 ( .A1(n1026), .A2(n1025), .Y(a2stg_frac1_in[40]) );
  AO22X1_RVT U1669 ( .A1(a1stg_intlngop), .A2(a1stg_in2[11]), .A3(
        a1stg_norm_dbl_in2), .A4(a1stg_in2[0]), .Y(n1112) );
  AO22X1_RVT U1670 ( .A1(n1030), .A2(n1112), .A3(n1027), .A4(a1stg_in1[0]), 
        .Y(n1028) );
  OR2X1_RVT U1671 ( .A1(n1029), .A2(n1028), .Y(a2stg_frac1_in[11]) );
  AND2X1_RVT U1672 ( .A1(a1stg_intlngop), .A2(n1030), .Y(n1031) );
  AND2X1_RVT U1673 ( .A1(a1stg_in2[10]), .A2(n1031), .Y(N1198) );
  AND2X1_RVT U1674 ( .A1(a1stg_in2[9]), .A2(n1031), .Y(N1206) );
  AND2X1_RVT U1675 ( .A1(a1stg_in2[8]), .A2(n1031), .Y(N1214) );
  AND2X1_RVT U1676 ( .A1(a1stg_in2[7]), .A2(n1031), .Y(N1222) );
  AND2X1_RVT U1677 ( .A1(a1stg_in2[6]), .A2(n1031), .Y(N1230) );
  AND2X1_RVT U1678 ( .A1(a1stg_in2[5]), .A2(n1031), .Y(N1238) );
  AND2X1_RVT U1679 ( .A1(a1stg_in2[4]), .A2(n1031), .Y(N1246) );
  AND2X1_RVT U1680 ( .A1(a1stg_in2[3]), .A2(n1031), .Y(N1254) );
  AND2X1_RVT U1681 ( .A1(a1stg_in2[2]), .A2(n1031), .Y(N1262) );
  AND2X1_RVT U1682 ( .A1(a1stg_in2[1]), .A2(n1031), .Y(N1270) );
  AND2X1_RVT U1683 ( .A1(a1stg_in2[0]), .A2(n1031), .Y(N1278) );
  AND2X1_RVT U1684 ( .A1(a1stg_in2_gt_in1), .A2(a2stg_frac2_in_frac1), .Y(
        n1082) );
  AO21X1_RVT U1685 ( .A1(a2stg_frac2_in_frac1), .A2(n1032), .A3(
        a1stg_faddsubop_inv), .Y(n1114) );
  AO22X1_RVT U1686 ( .A1(n1082), .A2(n1034), .A3(n1114), .A4(n1033), .Y(
        a2stg_frac2_in[63]) );
  OR2X1_RVT U1687 ( .A1(a2stg_frac2_in_qnan), .A2(n1035), .Y(n1036) );
  AO22X1_RVT U1688 ( .A1(n1082), .A2(n1037), .A3(n1114), .A4(n1036), .Y(
        a2stg_frac2_in[62]) );
  AO22X1_RVT U1689 ( .A1(n1082), .A2(n1039), .A3(n1038), .A4(n1114), .Y(
        a2stg_frac2_in[61]) );
  AO22X1_RVT U1690 ( .A1(n1082), .A2(n1041), .A3(n1040), .A4(n1114), .Y(
        a2stg_frac2_in[60]) );
  AO22X1_RVT U1691 ( .A1(n1082), .A2(n1043), .A3(n1042), .A4(n1114), .Y(
        a2stg_frac2_in[59]) );
  AO22X1_RVT U1692 ( .A1(n1082), .A2(n1045), .A3(n1044), .A4(n1114), .Y(
        a2stg_frac2_in[58]) );
  AO22X1_RVT U1693 ( .A1(n1082), .A2(n1047), .A3(n1046), .A4(n1114), .Y(
        a2stg_frac2_in[57]) );
  AO22X1_RVT U1694 ( .A1(n1082), .A2(n1049), .A3(n1048), .A4(n1114), .Y(
        a2stg_frac2_in[56]) );
  AO22X1_RVT U1695 ( .A1(n1082), .A2(n1051), .A3(n1050), .A4(n1114), .Y(
        a2stg_frac2_in[55]) );
  AO22X1_RVT U1696 ( .A1(n1082), .A2(n1053), .A3(n1052), .A4(n1114), .Y(
        a2stg_frac2_in[54]) );
  AO22X1_RVT U1697 ( .A1(n1082), .A2(n1055), .A3(n1054), .A4(n1114), .Y(
        a2stg_frac2_in[53]) );
  AO22X1_RVT U1698 ( .A1(n1082), .A2(n1057), .A3(n1056), .A4(n1114), .Y(
        a2stg_frac2_in[52]) );
  AO22X1_RVT U1699 ( .A1(n1082), .A2(n1059), .A3(n1058), .A4(n1114), .Y(
        a2stg_frac2_in[51]) );
  AO22X1_RVT U1700 ( .A1(n1082), .A2(n1061), .A3(n1060), .A4(n1114), .Y(
        a2stg_frac2_in[50]) );
  AO22X1_RVT U1701 ( .A1(n1082), .A2(n1063), .A3(n1062), .A4(n1114), .Y(
        a2stg_frac2_in[49]) );
  AO22X1_RVT U1702 ( .A1(n1082), .A2(n1065), .A3(n1064), .A4(n1114), .Y(
        a2stg_frac2_in[48]) );
  AO22X1_RVT U1703 ( .A1(n1082), .A2(n1067), .A3(n1066), .A4(n1114), .Y(
        a2stg_frac2_in[47]) );
  AO22X1_RVT U1704 ( .A1(n1082), .A2(n1069), .A3(n1068), .A4(n1114), .Y(
        a2stg_frac2_in[46]) );
  AO22X1_RVT U1705 ( .A1(n1082), .A2(n1071), .A3(n1070), .A4(n1114), .Y(
        a2stg_frac2_in[45]) );
  AO22X1_RVT U1706 ( .A1(n1082), .A2(n1073), .A3(n1072), .A4(n1114), .Y(
        a2stg_frac2_in[44]) );
  AO22X1_RVT U1707 ( .A1(n1082), .A2(n1075), .A3(n1074), .A4(n1114), .Y(
        a2stg_frac2_in[43]) );
  AO22X1_RVT U1708 ( .A1(n1082), .A2(n1077), .A3(n1076), .A4(n1114), .Y(
        a2stg_frac2_in[42]) );
  AO22X1_RVT U1709 ( .A1(n1082), .A2(n1079), .A3(n1078), .A4(n1114), .Y(
        a2stg_frac2_in[41]) );
  AO22X1_RVT U1710 ( .A1(n1082), .A2(n1081), .A3(n1114), .A4(n1080), .Y(
        a2stg_frac2_in[40]) );
  AND2X1_RVT U1711 ( .A1(a1stg_denorm_dbl_in1), .A2(n1082), .Y(n1110) );
  AND2X1_RVT U1712 ( .A1(a1stg_norm_dbl_in1), .A2(n1082), .Y(n1113) );
  AO222X1_RVT U1713 ( .A1(n1083), .A2(n1114), .A3(n1110), .A4(a1stg_in1[27]), 
        .A5(n1113), .A6(a1stg_in1[28]), .Y(a2stg_frac2_in[39]) );
  AO222X1_RVT U1714 ( .A1(n1084), .A2(n1114), .A3(n1110), .A4(a1stg_in1[26]), 
        .A5(n1113), .A6(a1stg_in1[27]), .Y(a2stg_frac2_in[38]) );
  AO222X1_RVT U1715 ( .A1(n1085), .A2(n1114), .A3(n1110), .A4(a1stg_in1[25]), 
        .A5(n1113), .A6(a1stg_in1[26]), .Y(a2stg_frac2_in[37]) );
  AO222X1_RVT U1716 ( .A1(n1086), .A2(n1114), .A3(n1110), .A4(a1stg_in1[24]), 
        .A5(n1113), .A6(a1stg_in1[25]), .Y(a2stg_frac2_in[36]) );
  AO222X1_RVT U1717 ( .A1(n1087), .A2(n1114), .A3(n1110), .A4(a1stg_in1[23]), 
        .A5(n1113), .A6(a1stg_in1[24]), .Y(a2stg_frac2_in[35]) );
  AO222X1_RVT U1718 ( .A1(n1088), .A2(n1114), .A3(n1110), .A4(a1stg_in1[22]), 
        .A5(n1113), .A6(a1stg_in1[23]), .Y(a2stg_frac2_in[34]) );
  AO222X1_RVT U1719 ( .A1(n1089), .A2(n1114), .A3(n1110), .A4(a1stg_in1[21]), 
        .A5(n1113), .A6(a1stg_in1[22]), .Y(a2stg_frac2_in[33]) );
  AO222X1_RVT U1720 ( .A1(n1090), .A2(n1114), .A3(n1110), .A4(a1stg_in1[20]), 
        .A5(n1113), .A6(a1stg_in1[21]), .Y(a2stg_frac2_in[32]) );
  AO222X1_RVT U1721 ( .A1(n1091), .A2(n1114), .A3(n1110), .A4(a1stg_in1[19]), 
        .A5(n1113), .A6(a1stg_in1[20]), .Y(a2stg_frac2_in[31]) );
  AO222X1_RVT U1722 ( .A1(n1092), .A2(n1114), .A3(n1110), .A4(a1stg_in1[18]), 
        .A5(n1113), .A6(a1stg_in1[19]), .Y(a2stg_frac2_in[30]) );
  AO222X1_RVT U1723 ( .A1(n1093), .A2(n1114), .A3(n1110), .A4(a1stg_in1[17]), 
        .A5(n1113), .A6(a1stg_in1[18]), .Y(a2stg_frac2_in[29]) );
  AO222X1_RVT U1724 ( .A1(n1094), .A2(n1114), .A3(n1110), .A4(a1stg_in1[16]), 
        .A5(n1113), .A6(a1stg_in1[17]), .Y(a2stg_frac2_in[28]) );
  AO222X1_RVT U1725 ( .A1(n1095), .A2(n1114), .A3(n1110), .A4(a1stg_in1[15]), 
        .A5(n1113), .A6(a1stg_in1[16]), .Y(a2stg_frac2_in[27]) );
  AO222X1_RVT U1726 ( .A1(n1096), .A2(n1114), .A3(n1110), .A4(a1stg_in1[14]), 
        .A5(n1113), .A6(a1stg_in1[15]), .Y(a2stg_frac2_in[26]) );
  AO222X1_RVT U1727 ( .A1(n1097), .A2(n1114), .A3(n1110), .A4(a1stg_in1[13]), 
        .A5(n1113), .A6(a1stg_in1[14]), .Y(a2stg_frac2_in[25]) );
  AO222X1_RVT U1728 ( .A1(n1098), .A2(n1114), .A3(n1110), .A4(a1stg_in1[12]), 
        .A5(n1113), .A6(a1stg_in1[13]), .Y(a2stg_frac2_in[24]) );
  AO222X1_RVT U1729 ( .A1(n1099), .A2(n1114), .A3(n1110), .A4(a1stg_in1[11]), 
        .A5(n1113), .A6(a1stg_in1[12]), .Y(a2stg_frac2_in[23]) );
  AO222X1_RVT U1730 ( .A1(n1100), .A2(n1114), .A3(n1110), .A4(a1stg_in1[10]), 
        .A5(n1113), .A6(a1stg_in1[11]), .Y(a2stg_frac2_in[22]) );
  AO222X1_RVT U1731 ( .A1(n1101), .A2(n1114), .A3(n1110), .A4(a1stg_in1[9]), 
        .A5(n1113), .A6(a1stg_in1[10]), .Y(a2stg_frac2_in[21]) );
  AO222X1_RVT U1732 ( .A1(n1102), .A2(n1114), .A3(n1110), .A4(a1stg_in1[8]), 
        .A5(n1113), .A6(a1stg_in1[9]), .Y(a2stg_frac2_in[20]) );
  AO222X1_RVT U1733 ( .A1(n1103), .A2(n1114), .A3(n1110), .A4(a1stg_in1[7]), 
        .A5(n1113), .A6(a1stg_in1[8]), .Y(a2stg_frac2_in[19]) );
  AO222X1_RVT U1734 ( .A1(n1104), .A2(n1114), .A3(n1110), .A4(a1stg_in1[6]), 
        .A5(n1113), .A6(a1stg_in1[7]), .Y(a2stg_frac2_in[18]) );
  AO222X1_RVT U1735 ( .A1(n1105), .A2(n1114), .A3(n1110), .A4(a1stg_in1[5]), 
        .A5(n1113), .A6(a1stg_in1[6]), .Y(a2stg_frac2_in[17]) );
  AO222X1_RVT U1736 ( .A1(n1106), .A2(n1114), .A3(n1110), .A4(a1stg_in1[4]), 
        .A5(n1113), .A6(a1stg_in1[5]), .Y(a2stg_frac2_in[16]) );
  AO222X1_RVT U1737 ( .A1(n1107), .A2(n1114), .A3(n1110), .A4(a1stg_in1[3]), 
        .A5(n1113), .A6(a1stg_in1[4]), .Y(a2stg_frac2_in[15]) );
  AO222X1_RVT U1738 ( .A1(n1108), .A2(n1114), .A3(n1110), .A4(a1stg_in1[2]), 
        .A5(n1113), .A6(a1stg_in1[3]), .Y(a2stg_frac2_in[14]) );
  AO222X1_RVT U1739 ( .A1(n1109), .A2(n1114), .A3(n1110), .A4(a1stg_in1[1]), 
        .A5(n1113), .A6(a1stg_in1[2]), .Y(a2stg_frac2_in[13]) );
  AO222X1_RVT U1740 ( .A1(n1111), .A2(n1114), .A3(n1110), .A4(a1stg_in1[0]), 
        .A5(n1113), .A6(a1stg_in1[1]), .Y(a2stg_frac2_in[12]) );
  AO22X1_RVT U1741 ( .A1(a1stg_in1[0]), .A2(n1113), .A3(n1112), .A4(n1114), 
        .Y(a2stg_frac2_in[11]) );
  AND2X1_RVT U1742 ( .A1(a1stg_intlngop), .A2(n1114), .Y(n1115) );
  AND2X1_RVT U1743 ( .A1(a1stg_in2[10]), .A2(n1115), .Y(N1601) );
  AND2X1_RVT U1744 ( .A1(a1stg_in2[9]), .A2(n1115), .Y(N1607) );
  AND2X1_RVT U1745 ( .A1(a1stg_in2[8]), .A2(n1115), .Y(N1613) );
  AND2X1_RVT U1746 ( .A1(a1stg_in2[7]), .A2(n1115), .Y(N1619) );
  AND2X1_RVT U1747 ( .A1(a1stg_in2[6]), .A2(n1115), .Y(N1625) );
  AND2X1_RVT U1748 ( .A1(a1stg_in2[5]), .A2(n1115), .Y(N1631) );
  AND2X1_RVT U1749 ( .A1(a1stg_in2[4]), .A2(n1115), .Y(N1637) );
  AND2X1_RVT U1750 ( .A1(a1stg_in2[3]), .A2(n1115), .Y(N1643) );
  AND2X1_RVT U1751 ( .A1(a1stg_in2[2]), .A2(n1115), .Y(N1649) );
  AND2X1_RVT U1752 ( .A1(a1stg_in2[1]), .A2(n1115), .Y(N1655) );
  AND2X1_RVT U1753 ( .A1(a1stg_in2[0]), .A2(n1115), .Y(N1661) );
  NAND4X0_RVT U1754 ( .A1(n1119), .A2(n1118), .A3(n1117), .A4(n1116), .Y(n1120) );
  NOR4X1_RVT U1755 ( .A1(a2stg_frac2[62]), .A2(a2stg_frac2[32]), .A3(
        a2stg_frac2[33]), .A4(n1120), .Y(n1152) );
  AND4X1_RVT U1756 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .Y(n1151)
         );
  AND4X1_RVT U1757 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), .Y(n1150)
         );
  AND4X1_RVT U1758 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .Y(n1148)
         );
  AND4X1_RVT U1759 ( .A1(n1136), .A2(n1135), .A3(n1134), .A4(n1133), .Y(n1147)
         );
  AND4X1_RVT U1760 ( .A1(n1140), .A2(n1139), .A3(n1138), .A4(n1137), .Y(n1146)
         );
  AND4X1_RVT U1761 ( .A1(n1144), .A2(n1143), .A3(n1142), .A4(n1141), .Y(n1145)
         );
  AND4X1_RVT U1762 ( .A1(n1148), .A2(n1147), .A3(n1146), .A4(n1145), .Y(n1149)
         );
  NAND4X0_RVT U1763 ( .A1(n1152), .A2(n1151), .A3(n1150), .A4(n1149), .Y(
        a2stg_frac2hi_neq_0) );
  AND4X1_RVT U1764 ( .A1(n1156), .A2(n1155), .A3(n1154), .A4(n1153), .Y(n1179)
         );
  AND4X1_RVT U1765 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .Y(n1178)
         );
  AND4X1_RVT U1766 ( .A1(n1164), .A2(n1163), .A3(n1162), .A4(n1161), .Y(n1176)
         );
  AND4X1_RVT U1767 ( .A1(n1168), .A2(n1167), .A3(n1166), .A4(n1165), .Y(n1175)
         );
  AND4X1_RVT U1768 ( .A1(n1172), .A2(n1171), .A3(n1170), .A4(n1169), .Y(n1174)
         );
  AND4X1_RVT U1769 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), .Y(n1177)
         );
  NAND3X0_RVT U1770 ( .A1(n1179), .A2(n1178), .A3(n1177), .Y(
        a2stg_frac2lo_neq_0) );
  INVX1_RVT U1771 ( .A(a2stg_exp[1]), .Y(n1182) );
  INVX1_RVT U1772 ( .A(a2stg_exp[2]), .Y(n1181) );
  INVX1_RVT U1773 ( .A(a2stg_exp[3]), .Y(n1180) );
  INVX1_RVT U1774 ( .A(a2stg_exp[0]), .Y(n1183) );
  AND4X1_RVT U1775 ( .A1(n1182), .A2(n1181), .A3(n1180), .A4(n1183), .Y(n1199)
         );
  INVX1_RVT U1776 ( .A(a2stg_exp[5]), .Y(n1185) );
  INVX1_RVT U1777 ( .A(a2stg_exp[4]), .Y(n1187) );
  AND3X1_RVT U1778 ( .A1(a2stg_expdec_neq_0), .A2(n1185), .A3(n1187), .Y(n1184) );
  AND2X1_RVT U1779 ( .A1(n1199), .A2(n1184), .Y(a2stg_expdec[53]) );
  AND4X1_RVT U1780 ( .A1(a2stg_exp[0]), .A2(n1182), .A3(n1181), .A4(n1180), 
        .Y(n1200) );
  AND2X1_RVT U1781 ( .A1(n1184), .A2(n1200), .Y(a2stg_expdec[52]) );
  AND4X1_RVT U1782 ( .A1(a2stg_exp[1]), .A2(n1180), .A3(n1181), .A4(n1183), 
        .Y(n1201) );
  AND2X1_RVT U1783 ( .A1(n1184), .A2(n1201), .Y(a2stg_expdec[51]) );
  AND4X1_RVT U1784 ( .A1(a2stg_exp[1]), .A2(a2stg_exp[0]), .A3(n1180), .A4(
        n1181), .Y(n1202) );
  AND2X1_RVT U1785 ( .A1(n1184), .A2(n1202), .Y(a2stg_expdec[50]) );
  AND4X1_RVT U1786 ( .A1(a2stg_exp[2]), .A2(n1182), .A3(n1180), .A4(n1183), 
        .Y(n1203) );
  AND2X1_RVT U1787 ( .A1(n1184), .A2(n1203), .Y(a2stg_expdec[49]) );
  AND4X1_RVT U1788 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[0]), .A3(n1182), .A4(
        n1180), .Y(n1205) );
  AND2X1_RVT U1789 ( .A1(n1184), .A2(n1205), .Y(a2stg_expdec[48]) );
  AND4X1_RVT U1790 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[1]), .A3(n1180), .A4(
        n1183), .Y(n1188) );
  AND2X1_RVT U1791 ( .A1(n1184), .A2(n1188), .Y(a2stg_expdec[47]) );
  AND4X1_RVT U1792 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[1]), .A3(a2stg_exp[0]), 
        .A4(n1180), .Y(n1189) );
  AND2X1_RVT U1793 ( .A1(n1184), .A2(n1189), .Y(a2stg_expdec[46]) );
  AND4X1_RVT U1794 ( .A1(a2stg_exp[3]), .A2(n1182), .A3(n1181), .A4(n1183), 
        .Y(n1190) );
  AND2X1_RVT U1795 ( .A1(n1184), .A2(n1190), .Y(a2stg_expdec[45]) );
  AND4X1_RVT U1796 ( .A1(a2stg_exp[3]), .A2(a2stg_exp[0]), .A3(n1182), .A4(
        n1181), .Y(n1191) );
  AND2X1_RVT U1797 ( .A1(n1184), .A2(n1191), .Y(a2stg_expdec[44]) );
  AND4X1_RVT U1798 ( .A1(a2stg_exp[1]), .A2(a2stg_exp[3]), .A3(n1181), .A4(
        n1183), .Y(n1192) );
  AND2X1_RVT U1799 ( .A1(n1184), .A2(n1192), .Y(a2stg_expdec[43]) );
  AND4X1_RVT U1800 ( .A1(a2stg_exp[1]), .A2(a2stg_exp[3]), .A3(a2stg_exp[0]), 
        .A4(n1181), .Y(n1193) );
  AND2X1_RVT U1801 ( .A1(n1184), .A2(n1193), .Y(a2stg_expdec[42]) );
  AND4X1_RVT U1802 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[3]), .A3(n1182), .A4(
        n1183), .Y(n1194) );
  AND2X1_RVT U1803 ( .A1(n1184), .A2(n1194), .Y(a2stg_expdec[41]) );
  AND4X1_RVT U1804 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[3]), .A3(a2stg_exp[0]), 
        .A4(n1182), .Y(n1195) );
  AND2X1_RVT U1805 ( .A1(n1184), .A2(n1195), .Y(a2stg_expdec[40]) );
  AND4X1_RVT U1806 ( .A1(a2stg_exp[2]), .A2(a2stg_exp[1]), .A3(a2stg_exp[3]), 
        .A4(n1183), .Y(n1196) );
  AND2X1_RVT U1807 ( .A1(n1184), .A2(n1196), .Y(a2stg_expdec[39]) );
  AND4X1_RVT U1808 ( .A1(a2stg_exp[1]), .A2(a2stg_exp[2]), .A3(a2stg_exp[3]), 
        .A4(a2stg_exp[0]), .Y(n1198) );
  AND2X1_RVT U1809 ( .A1(n1184), .A2(n1198), .Y(a2stg_expdec[38]) );
  AND3X1_RVT U1810 ( .A1(a2stg_expdec_neq_0), .A2(a2stg_exp[4]), .A3(n1185), 
        .Y(n1186) );
  AND2X1_RVT U1811 ( .A1(n1199), .A2(n1186), .Y(a2stg_expdec[37]) );
  AND2X1_RVT U1812 ( .A1(n1200), .A2(n1186), .Y(a2stg_expdec[36]) );
  AND2X1_RVT U1813 ( .A1(n1201), .A2(n1186), .Y(a2stg_expdec[35]) );
  AND2X1_RVT U1814 ( .A1(n1202), .A2(n1186), .Y(a2stg_expdec[34]) );
  AND2X1_RVT U1815 ( .A1(n1203), .A2(n1186), .Y(a2stg_expdec[33]) );
  AND2X1_RVT U1816 ( .A1(n1205), .A2(n1186), .Y(a2stg_expdec[32]) );
  AND2X1_RVT U1817 ( .A1(n1188), .A2(n1186), .Y(a2stg_expdec[31]) );
  AND2X1_RVT U1818 ( .A1(n1189), .A2(n1186), .Y(a2stg_expdec[30]) );
  AND2X1_RVT U1819 ( .A1(n1190), .A2(n1186), .Y(a2stg_expdec[29]) );
  AND2X1_RVT U1820 ( .A1(n1191), .A2(n1186), .Y(a2stg_expdec[28]) );
  AND2X1_RVT U1821 ( .A1(n1192), .A2(n1186), .Y(a2stg_expdec[27]) );
  AND2X1_RVT U1822 ( .A1(n1193), .A2(n1186), .Y(a2stg_expdec[26]) );
  AND2X1_RVT U1823 ( .A1(n1194), .A2(n1186), .Y(a2stg_expdec[25]) );
  AND2X1_RVT U1824 ( .A1(n1195), .A2(n1186), .Y(a2stg_expdec[24]) );
  AND2X1_RVT U1825 ( .A1(n1196), .A2(n1186), .Y(a2stg_expdec[23]) );
  AND2X1_RVT U1826 ( .A1(n1198), .A2(n1186), .Y(a2stg_expdec[22]) );
  AND3X1_RVT U1827 ( .A1(a2stg_expdec_neq_0), .A2(a2stg_exp[5]), .A3(n1187), 
        .Y(n1197) );
  AND2X1_RVT U1828 ( .A1(n1199), .A2(n1197), .Y(a2stg_expdec[21]) );
  AND2X1_RVT U1829 ( .A1(n1200), .A2(n1197), .Y(a2stg_expdec[20]) );
  AND2X1_RVT U1830 ( .A1(n1201), .A2(n1197), .Y(a2stg_expdec[19]) );
  AND2X1_RVT U1831 ( .A1(n1202), .A2(n1197), .Y(a2stg_expdec[18]) );
  AND2X1_RVT U1832 ( .A1(n1203), .A2(n1197), .Y(a2stg_expdec[17]) );
  AND2X1_RVT U1833 ( .A1(n1205), .A2(n1197), .Y(a2stg_expdec[16]) );
  AND2X1_RVT U1834 ( .A1(n1188), .A2(n1197), .Y(a2stg_expdec[15]) );
  AND2X1_RVT U1835 ( .A1(n1189), .A2(n1197), .Y(a2stg_expdec[14]) );
  AND2X1_RVT U1836 ( .A1(n1190), .A2(n1197), .Y(a2stg_expdec[13]) );
  AND2X1_RVT U1837 ( .A1(n1191), .A2(n1197), .Y(a2stg_expdec[12]) );
  AND2X1_RVT U1838 ( .A1(n1192), .A2(n1197), .Y(a2stg_expdec[11]) );
  AND2X1_RVT U1839 ( .A1(n1193), .A2(n1197), .Y(a2stg_expdec[10]) );
  AND2X1_RVT U1840 ( .A1(n1194), .A2(n1197), .Y(a2stg_expdec[9]) );
  AND2X1_RVT U1841 ( .A1(n1195), .A2(n1197), .Y(a2stg_expdec[8]) );
  AND2X1_RVT U1842 ( .A1(n1196), .A2(n1197), .Y(a2stg_expdec[7]) );
  AND2X1_RVT U1843 ( .A1(n1198), .A2(n1197), .Y(a2stg_expdec[6]) );
  AND3X1_RVT U1844 ( .A1(a2stg_exp[5]), .A2(a2stg_expdec_neq_0), .A3(
        a2stg_exp[4]), .Y(n1204) );
  AND2X1_RVT U1845 ( .A1(n1199), .A2(n1204), .Y(a2stg_expdec[5]) );
  AND2X1_RVT U1846 ( .A1(n1200), .A2(n1204), .Y(a2stg_expdec[4]) );
  AND2X1_RVT U1847 ( .A1(n1201), .A2(n1204), .Y(a2stg_expdec[3]) );
  AND2X1_RVT U1848 ( .A1(n1202), .A2(n1204), .Y(a2stg_expdec[2]) );
  AND2X1_RVT U1849 ( .A1(n1203), .A2(n1204), .Y(a2stg_expdec[1]) );
  AND2X1_RVT U1850 ( .A1(n1205), .A2(n1204), .Y(a2stg_expdec[0]) );
  NOR4X1_RVT U1851 ( .A1(a3stg_ld0_frac[1]), .A2(a3stg_ld0_frac[0]), .A3(
        a3stg_ld0_frac[2]), .A4(a3stg_ld0_frac[3]), .Y(n1209) );
  NOR4X1_RVT U1852 ( .A1(a3stg_ld0_frac[6]), .A2(a3stg_ld0_frac[7]), .A3(
        a3stg_ld0_frac[8]), .A4(a3stg_ld0_frac[9]), .Y(n1208) );
  NAND4X0_RVT U1853 ( .A1(n1209), .A2(n1208), .A3(n1207), .A4(n1206), .Y(n1210) );
  AO21X1_RVT U1854 ( .A1(n1211), .A2(n1210), .A3(a3stg_ld0_frac[10]), .Y(
        a3stg_ld0_dnrm_10) );
  FADDX1_RVT U1855 ( .A(a3stg_frac1[60]), .B(a3stg_frac2[60]), .CI(n1212), 
        .CO(n410), .S(n1429) );
  AND2X1_RVT U1856 ( .A1(n1429), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[62]) );
  FADDX1_RVT U1857 ( .A(a3stg_frac1[59]), .B(a3stg_frac2[59]), .CI(n1213), 
        .CO(n1212), .S(n1437) );
  AND2X1_RVT U1858 ( .A1(n1437), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[61]) );
  FADDX1_RVT U1859 ( .A(a3stg_frac1[58]), .B(a3stg_frac2[58]), .CI(n1214), 
        .CO(n1213), .S(n1445) );
  AND2X1_RVT U1860 ( .A1(n1445), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[60]) );
  FADDX1_RVT U1861 ( .A(a3stg_frac1[57]), .B(a3stg_frac2[57]), .CI(n1215), 
        .CO(n1214), .S(n1453) );
  AND2X1_RVT U1862 ( .A1(n1453), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[59]) );
  FADDX1_RVT U1863 ( .A(a3stg_frac1[56]), .B(a3stg_frac2[56]), .CI(n1216), 
        .CO(n1215), .S(n1462) );
  AND2X1_RVT U1864 ( .A1(n1462), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[58]) );
  FADDX1_RVT U1865 ( .A(a3stg_frac1[55]), .B(a3stg_frac2[55]), .CI(n1217), 
        .CO(n1216), .S(n1469) );
  AND2X1_RVT U1866 ( .A1(n1469), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[57]) );
  FADDX1_RVT U1867 ( .A(a3stg_frac1[54]), .B(a3stg_frac2[54]), .CI(n1218), 
        .CO(n1217), .S(n1476) );
  AND2X1_RVT U1868 ( .A1(n1476), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[56]) );
  FADDX1_RVT U1869 ( .A(a3stg_frac1[53]), .B(a3stg_frac2[53]), .CI(n1219), 
        .CO(n1218), .S(n1483) );
  AND2X1_RVT U1870 ( .A1(n1483), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[55]) );
  FADDX1_RVT U1871 ( .A(a3stg_frac1[52]), .B(a3stg_frac2[52]), .CI(n1220), 
        .CO(n1219), .S(n1490) );
  AND2X1_RVT U1872 ( .A1(n1490), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[54]) );
  FADDX1_RVT U1873 ( .A(a3stg_frac1[51]), .B(a3stg_frac2[51]), .CI(n1221), 
        .CO(n1220), .S(n1497) );
  AND2X1_RVT U1874 ( .A1(n1497), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[53]) );
  FADDX1_RVT U1875 ( .A(a3stg_frac1[50]), .B(a3stg_frac2[50]), .CI(n1222), 
        .CO(n1221), .S(n1504) );
  AND2X1_RVT U1876 ( .A1(n1504), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[52]) );
  FADDX1_RVT U1877 ( .A(a3stg_frac1[49]), .B(a3stg_frac2[49]), .CI(n1223), 
        .CO(n1222), .S(n1511) );
  AND2X1_RVT U1878 ( .A1(n1511), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[51]) );
  FADDX1_RVT U1879 ( .A(a3stg_frac1[48]), .B(a3stg_frac2[48]), .CI(n1224), 
        .CO(n1223), .S(n1518) );
  AND2X1_RVT U1880 ( .A1(n1518), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[50]) );
  FADDX1_RVT U1881 ( .A(a3stg_frac1[47]), .B(a3stg_frac2[47]), .CI(n1225), 
        .CO(n1224), .S(n1525) );
  AND2X1_RVT U1882 ( .A1(n1525), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[49]) );
  FADDX1_RVT U1883 ( .A(a3stg_frac1[46]), .B(a3stg_frac2[46]), .CI(n1226), 
        .CO(n1225), .S(n1532) );
  AND2X1_RVT U1884 ( .A1(n1532), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[48]) );
  FADDX1_RVT U1885 ( .A(a3stg_frac1[45]), .B(a3stg_frac2[45]), .CI(n1227), 
        .CO(n1226), .S(n1539) );
  AND2X1_RVT U1886 ( .A1(n1539), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[47]) );
  FADDX1_RVT U1887 ( .A(a3stg_frac1[44]), .B(a3stg_frac2[44]), .CI(n1228), 
        .CO(n1227), .S(n1547) );
  AND2X1_RVT U1888 ( .A1(n1547), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[46]) );
  FADDX1_RVT U1889 ( .A(a3stg_frac1[43]), .B(a3stg_frac2[43]), .CI(n1229), 
        .CO(n1228), .S(n1554) );
  AND2X1_RVT U1890 ( .A1(n1554), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[45]) );
  FADDX1_RVT U1891 ( .A(a3stg_frac1[42]), .B(a3stg_frac2[42]), .CI(n1230), 
        .CO(n1229), .S(n1561) );
  AND2X1_RVT U1892 ( .A1(n1561), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[44]) );
  FADDX1_RVT U1893 ( .A(a3stg_frac1[41]), .B(a3stg_frac2[41]), .CI(n1231), 
        .CO(n1230), .S(n1568) );
  AND2X1_RVT U1894 ( .A1(n1568), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[43]) );
  FADDX1_RVT U1895 ( .A(a3stg_frac1[40]), .B(a3stg_frac2[40]), .CI(n1232), 
        .CO(n1231), .S(n1575) );
  AND2X1_RVT U1896 ( .A1(n1575), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[42]) );
  FADDX1_RVT U1897 ( .A(a3stg_frac1[39]), .B(a3stg_frac2[39]), .CI(n1233), 
        .CO(n1232), .S(n1582) );
  AND2X1_RVT U1898 ( .A1(n1582), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[41]) );
  FADDX1_RVT U1899 ( .A(a3stg_frac1[38]), .B(a3stg_frac2[38]), .CI(n1234), 
        .CO(n1233), .S(n1589) );
  AND2X1_RVT U1900 ( .A1(n1589), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[40]) );
  FADDX1_RVT U1901 ( .A(a3stg_frac1[37]), .B(a3stg_frac2[37]), .CI(n1235), 
        .CO(n1234), .S(n1596) );
  AND2X1_RVT U1902 ( .A1(n1596), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[39]) );
  FADDX1_RVT U1903 ( .A(a3stg_frac1[36]), .B(a3stg_frac2[36]), .CI(n1236), 
        .CO(n1235), .S(n1603) );
  AND2X1_RVT U1904 ( .A1(n1603), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[38]) );
  FADDX1_RVT U1905 ( .A(a3stg_frac1[35]), .B(a3stg_frac2[35]), .CI(n1237), 
        .CO(n1236), .S(n1610) );
  AND2X1_RVT U1906 ( .A1(n1610), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[37]) );
  FADDX1_RVT U1907 ( .A(a3stg_frac1[34]), .B(a3stg_frac2[34]), .CI(n1238), 
        .CO(n1237), .S(n1617) );
  AND2X1_RVT U1908 ( .A1(n1617), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[36]) );
  FADDX1_RVT U1909 ( .A(a3stg_frac1[33]), .B(a3stg_frac2[33]), .CI(n1239), 
        .CO(n1238), .S(n1624) );
  AND2X1_RVT U1910 ( .A1(n1624), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[35]) );
  FADDX1_RVT U1911 ( .A(a3stg_frac1[32]), .B(a3stg_frac2[32]), .CI(n1240), 
        .CO(n1239), .S(n1631) );
  AND2X1_RVT U1912 ( .A1(n1631), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[34]) );
  FADDX1_RVT U1913 ( .A(a3stg_frac1[31]), .B(a3stg_frac2[31]), .CI(n1241), 
        .CO(n1240), .S(n1638) );
  AND2X1_RVT U1914 ( .A1(n1638), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[33]) );
  FADDX1_RVT U1915 ( .A(a3stg_frac1[30]), .B(a3stg_frac2[30]), .CI(n1242), 
        .CO(n1241), .S(n1645) );
  AND2X1_RVT U1916 ( .A1(n1645), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[32]) );
  FADDX1_RVT U1917 ( .A(a3stg_frac1[29]), .B(a3stg_frac2[29]), .CI(n1243), 
        .CO(n1242), .S(n1651) );
  AND2X1_RVT U1918 ( .A1(n1651), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[31]) );
  FADDX1_RVT U1919 ( .A(a3stg_frac1[28]), .B(a3stg_frac2[28]), .CI(n1244), 
        .CO(n1243), .S(n1657) );
  AND2X1_RVT U1920 ( .A1(n1657), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[30]) );
  FADDX1_RVT U1921 ( .A(a3stg_frac1[27]), .B(a3stg_frac2[27]), .CI(n1245), 
        .CO(n1244), .S(n1663) );
  AND2X1_RVT U1922 ( .A1(n1663), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[29]) );
  FADDX1_RVT U1923 ( .A(a3stg_frac1[26]), .B(a3stg_frac2[26]), .CI(n1246), 
        .CO(n1245), .S(n1734) );
  AND2X1_RVT U1924 ( .A1(n1734), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[28]) );
  FADDX1_RVT U1925 ( .A(a3stg_frac1[25]), .B(a3stg_frac2[25]), .CI(n1247), 
        .CO(n1246), .S(n1742) );
  AND2X1_RVT U1926 ( .A1(n1742), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[27]) );
  FADDX1_RVT U1927 ( .A(a3stg_frac1[24]), .B(a3stg_frac2[24]), .CI(n1248), 
        .CO(n1247), .S(n1748) );
  AND2X1_RVT U1928 ( .A1(n1748), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[26]) );
  FADDX1_RVT U1929 ( .A(a3stg_frac1[23]), .B(a3stg_frac2[23]), .CI(n1249), 
        .CO(n1248), .S(n1754) );
  AND2X1_RVT U1930 ( .A1(n1754), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[25]) );
  FADDX1_RVT U1931 ( .A(a3stg_frac1[22]), .B(a3stg_frac2[22]), .CI(n1250), 
        .CO(n1249), .S(n1760) );
  AND2X1_RVT U1932 ( .A1(n1760), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[24]) );
  AOI21X1_RVT U1933 ( .A1(n1253), .A2(n1291), .A3(n1252), .Y(n1256) );
  NAND2X0_RVT U1934 ( .A1(n3), .A2(n1254), .Y(n1255) );
  XOR2X1_RVT U1935 ( .A1(n1256), .A2(n1255), .Y(n1766) );
  AND2X1_RVT U1936 ( .A1(n1766), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[23]) );
  AOI21X1_RVT U1937 ( .A1(n1260), .A2(n1291), .A3(n1259), .Y(n1268) );
  OAI21X1_RVT U1938 ( .A1(n1261), .A2(n1268), .A3(n1265), .Y(n1264) );
  NAND2X0_RVT U1939 ( .A1(n4), .A2(n1262), .Y(n1263) );
  XNOR2X1_RVT U1940 ( .A1(n1264), .A2(n1263), .Y(n1772) );
  AND2X1_RVT U1941 ( .A1(n1772), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[22]) );
  NAND2X0_RVT U1942 ( .A1(n1266), .A2(n1265), .Y(n1267) );
  XOR2X1_RVT U1943 ( .A1(n1268), .A2(n1267), .Y(n1778) );
  AND2X1_RVT U1944 ( .A1(n1778), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[21]) );
  AOI21X1_RVT U1945 ( .A1(n1270), .A2(n1291), .A3(n1269), .Y(n1280) );
  OAI21X1_RVT U1946 ( .A1(n1276), .A2(n1280), .A3(n1277), .Y(n1275) );
  NAND2X0_RVT U1947 ( .A1(n1273), .A2(n1272), .Y(n1274) );
  XNOR2X1_RVT U1948 ( .A1(n1275), .A2(n1274), .Y(n1784) );
  AND2X1_RVT U1949 ( .A1(n1784), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[20]) );
  NAND2X0_RVT U1950 ( .A1(n1278), .A2(n1277), .Y(n1279) );
  XOR2X1_RVT U1951 ( .A1(n1280), .A2(n1279), .Y(n1790) );
  AND2X1_RVT U1952 ( .A1(n1790), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[19]) );
  AOI21X1_RVT U1953 ( .A1(n1289), .A2(n1291), .A3(n1282), .Y(n1287) );
  NAND2X0_RVT U1954 ( .A1(n1285), .A2(n1284), .Y(n1286) );
  XOR2X1_RVT U1955 ( .A1(n1287), .A2(n1286), .Y(n1797) );
  AND2X1_RVT U1956 ( .A1(n1797), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[18]) );
  NAND2X0_RVT U1957 ( .A1(n1289), .A2(n1288), .Y(n1290) );
  XNOR2X1_RVT U1958 ( .A1(n1291), .A2(n1290), .Y(n1804) );
  AND2X1_RVT U1959 ( .A1(n1804), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[17]) );
  OAI21X1_RVT U1960 ( .A1(n1296), .A2(n1346), .A3(n1295), .Y(n1312) );
  INVX1_RVT U1961 ( .A(n1312), .Y(n1321) );
  OAI21X1_RVT U1962 ( .A1(n1299), .A2(n1321), .A3(n1298), .Y(n1309) );
  AOI21X1_RVT U1963 ( .A1(n1307), .A2(n1309), .A3(n1300), .Y(n1305) );
  NAND2X0_RVT U1964 ( .A1(n1303), .A2(n1302), .Y(n1304) );
  XOR2X1_RVT U1965 ( .A1(n1305), .A2(n1304), .Y(n1809) );
  AND2X1_RVT U1966 ( .A1(n1809), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[16]) );
  NAND2X0_RVT U1967 ( .A1(n1307), .A2(n1306), .Y(n1308) );
  XNOR2X1_RVT U1968 ( .A1(n1309), .A2(n1308), .Y(n1816) );
  AND2X1_RVT U1969 ( .A1(n1816), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[15]) );
  AOI21X1_RVT U1970 ( .A1(n1319), .A2(n1312), .A3(n1311), .Y(n1317) );
  NAND2X0_RVT U1971 ( .A1(n1315), .A2(n1314), .Y(n1316) );
  XOR2X1_RVT U1972 ( .A1(n1317), .A2(n1316), .Y(n1823) );
  AND2X1_RVT U1973 ( .A1(n1823), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[14]) );
  NAND2X0_RVT U1974 ( .A1(n1319), .A2(n1318), .Y(n1320) );
  XOR2X1_RVT U1975 ( .A1(n1321), .A2(n1320), .Y(n1828) );
  AND2X1_RVT U1976 ( .A1(n1828), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[13]) );
  OAI21X1_RVT U1977 ( .A1(n1326), .A2(n1346), .A3(n1325), .Y(n1336) );
  AOI21X1_RVT U1978 ( .A1(n1334), .A2(n1336), .A3(n1327), .Y(n1332) );
  NAND2X0_RVT U1979 ( .A1(n1330), .A2(n1329), .Y(n1331) );
  XOR2X1_RVT U1980 ( .A1(n1332), .A2(n1331), .Y(n1833) );
  AND2X1_RVT U1981 ( .A1(n1833), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[12]) );
  NAND2X0_RVT U1982 ( .A1(n1334), .A2(n1333), .Y(n1335) );
  XNOR2X1_RVT U1983 ( .A1(n1336), .A2(n1335), .Y(n1837) );
  AND2X1_RVT U1984 ( .A1(n1837), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[11]) );
  OAI21X1_RVT U1985 ( .A1(n1342), .A2(n1346), .A3(n1343), .Y(n1341) );
  NAND2X0_RVT U1986 ( .A1(n1339), .A2(n1338), .Y(n1340) );
  XNOR2X1_RVT U1987 ( .A1(n1341), .A2(n1340), .Y(n1842) );
  AND2X1_RVT U1988 ( .A1(n1842), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[10]) );
  NAND2X0_RVT U1989 ( .A1(n1344), .A2(n1343), .Y(n1345) );
  XOR2X1_RVT U1990 ( .A1(n1346), .A2(n1345), .Y(n1846) );
  AND2X1_RVT U1991 ( .A1(n1846), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[9]) );
  AOI21X1_RVT U1992 ( .A1(n1349), .A2(n1370), .A3(n1348), .Y(n1359) );
  OAI21X1_RVT U1993 ( .A1(n1355), .A2(n1359), .A3(n1356), .Y(n1354) );
  NAND2X0_RVT U1994 ( .A1(n1352), .A2(n1351), .Y(n1353) );
  XNOR2X1_RVT U1995 ( .A1(n1354), .A2(n1353), .Y(n1850) );
  AND2X1_RVT U1996 ( .A1(n1850), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[8]) );
  NAND2X0_RVT U1997 ( .A1(n1357), .A2(n1356), .Y(n1358) );
  XOR2X1_RVT U1998 ( .A1(n1359), .A2(n1358), .Y(n1854) );
  AND2X1_RVT U1999 ( .A1(n1854), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[7]) );
  AOI21X1_RVT U2000 ( .A1(n1368), .A2(n1370), .A3(n1361), .Y(n1366) );
  NAND2X0_RVT U2001 ( .A1(n1364), .A2(n1363), .Y(n1365) );
  XOR2X1_RVT U2002 ( .A1(n1366), .A2(n1365), .Y(n1858) );
  AND2X1_RVT U2003 ( .A1(n1858), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[6]) );
  NAND2X0_RVT U2004 ( .A1(n1368), .A2(n1367), .Y(n1369) );
  XNOR2X1_RVT U2005 ( .A1(n1370), .A2(n1369), .Y(n1862) );
  AND2X1_RVT U2006 ( .A1(n1862), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[5]) );
  INVX1_RVT U2007 ( .A(n1371), .Y(n1381) );
  OAI21X1_RVT U2008 ( .A1(n1377), .A2(n1381), .A3(n1378), .Y(n1376) );
  NAND2X0_RVT U2009 ( .A1(n1374), .A2(n1373), .Y(n1375) );
  XNOR2X1_RVT U2010 ( .A1(n1376), .A2(n1375), .Y(n1865) );
  AND2X1_RVT U2011 ( .A1(n1865), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[4]) );
  NAND2X0_RVT U2012 ( .A1(n1379), .A2(n1378), .Y(n1380) );
  XOR2X1_RVT U2013 ( .A1(n1381), .A2(n1380), .Y(n1869) );
  AND2X1_RVT U2014 ( .A1(n1869), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[3]) );
  NAND2X0_RVT U2015 ( .A1(n1384), .A2(n1383), .Y(n1385) );
  XNOR2X1_RVT U2016 ( .A1(n1385), .A2(a3stg_frac2[0]), .Y(n1876) );
  AND2X1_RVT U2017 ( .A1(n1876), .A2(n2542), .Y(a4stg_rnd_frac_pre1_in[2]) );
  AND2X1_RVT U2018 ( .A1(n1919), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[62]) );
  AND2X1_RVT U2019 ( .A1(n1429), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[61]) );
  AND2X1_RVT U2020 ( .A1(n1437), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[60]) );
  AND2X1_RVT U2021 ( .A1(n1445), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[59]) );
  AND2X1_RVT U2022 ( .A1(n1453), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[58]) );
  AND2X1_RVT U2023 ( .A1(n1462), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[57]) );
  AND2X1_RVT U2024 ( .A1(n1469), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[56]) );
  AND2X1_RVT U2025 ( .A1(n1476), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[55]) );
  AND2X1_RVT U2026 ( .A1(n1483), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[54]) );
  AND2X1_RVT U2027 ( .A1(n1490), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[53]) );
  AND2X1_RVT U2028 ( .A1(n1497), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[52]) );
  AND2X1_RVT U2029 ( .A1(n1504), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[51]) );
  AND2X1_RVT U2030 ( .A1(n1511), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[50]) );
  AND2X1_RVT U2031 ( .A1(n1518), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[49]) );
  AND2X1_RVT U2032 ( .A1(n1525), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[48]) );
  AND2X1_RVT U2033 ( .A1(n1532), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[47]) );
  AND2X1_RVT U2034 ( .A1(n1539), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[46]) );
  AND2X1_RVT U2035 ( .A1(n1547), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[45]) );
  AND2X1_RVT U2036 ( .A1(n1554), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[44]) );
  AND2X1_RVT U2037 ( .A1(n1561), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[43]) );
  AND2X1_RVT U2038 ( .A1(n1568), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[42]) );
  AND2X1_RVT U2039 ( .A1(n1575), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[41]) );
  AND2X1_RVT U2040 ( .A1(n1582), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[40]) );
  AND2X1_RVT U2041 ( .A1(n1589), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[39]) );
  AND2X1_RVT U2042 ( .A1(n1596), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[38]) );
  AND2X1_RVT U2043 ( .A1(n1603), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[37]) );
  AND2X1_RVT U2044 ( .A1(n1610), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[36]) );
  AND2X1_RVT U2045 ( .A1(n1617), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[35]) );
  AND2X1_RVT U2046 ( .A1(n1624), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[34]) );
  AND2X1_RVT U2047 ( .A1(n1631), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[33]) );
  AND2X1_RVT U2048 ( .A1(n1638), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[32]) );
  AND2X1_RVT U2049 ( .A1(n1645), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[31]) );
  AND2X1_RVT U2050 ( .A1(n1651), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[30]) );
  AND2X1_RVT U2051 ( .A1(n1657), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[29]) );
  AND2X1_RVT U2052 ( .A1(n1663), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[28]) );
  AND2X1_RVT U2053 ( .A1(n1734), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[27]) );
  AND2X1_RVT U2054 ( .A1(n1742), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[26]) );
  AND2X1_RVT U2055 ( .A1(n1748), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[25]) );
  AND2X1_RVT U2056 ( .A1(n1754), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[24]) );
  AND2X1_RVT U2057 ( .A1(n1760), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[23]) );
  AND2X1_RVT U2058 ( .A1(n1766), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[22]) );
  AND2X1_RVT U2059 ( .A1(n1772), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[21]) );
  AND2X1_RVT U2060 ( .A1(n1778), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[20]) );
  AND2X1_RVT U2061 ( .A1(n1784), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[19]) );
  AND2X1_RVT U2062 ( .A1(n1790), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[18]) );
  AND2X1_RVT U2063 ( .A1(n1797), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[17]) );
  AND2X1_RVT U2064 ( .A1(n1804), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[16]) );
  AND2X1_RVT U2065 ( .A1(n1809), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[15]) );
  AND2X1_RVT U2066 ( .A1(n1816), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[14]) );
  AND2X1_RVT U2067 ( .A1(n1823), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[13]) );
  AND2X1_RVT U2068 ( .A1(n1828), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[12]) );
  AND2X1_RVT U2069 ( .A1(n1833), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[11]) );
  AND2X1_RVT U2070 ( .A1(n1837), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[10]) );
  AND2X1_RVT U2071 ( .A1(n1842), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[9]) );
  AND2X1_RVT U2072 ( .A1(n1846), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[8]) );
  AND2X1_RVT U2073 ( .A1(n1850), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[7]) );
  AND2X1_RVT U2074 ( .A1(n1854), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[6]) );
  AND2X1_RVT U2075 ( .A1(n1858), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[5]) );
  AND2X1_RVT U2076 ( .A1(n1862), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[4]) );
  AND2X1_RVT U2077 ( .A1(n1865), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[3]) );
  AND2X1_RVT U2078 ( .A1(n1869), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[2]) );
  AND2X1_RVT U2079 ( .A1(n1876), .A2(n1), .Y(a4stg_rnd_frac_pre3_in[1]) );
  AND2X1_RVT U2080 ( .A1(a4stg_shl_cnt[0]), .A2(n1813), .Y(n1389) );
  AO22X1_RVT U2081 ( .A1(a4stg_shl_cnt[0]), .A2(n1388), .A3(n1800), .A4(n1387), 
        .Y(n1420) );
  AO222X1_RVT U2082 ( .A1(n1391), .A2(n1820), .A3(n1390), .A4(n1389), .A5(
        n1420), .A6(a4stg_shl_cnt[1]), .Y(n1403) );
  AO22X1_RVT U2083 ( .A1(a4stg_shl_cnt[0]), .A2(n1393), .A3(n1800), .A4(n1392), 
        .Y(n1425) );
  AO22X1_RVT U2084 ( .A1(a4stg_shl_cnt[0]), .A2(n1395), .A3(n1800), .A4(n1394), 
        .Y(n1419) );
  AO22X1_RVT U2085 ( .A1(a4stg_shl_cnt[1]), .A2(n1425), .A3(n1813), .A4(n1419), 
        .Y(n1444) );
  AO222X1_RVT U2086 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[15]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[47]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[31]), .Y(n1409) );
  AO22X1_RVT U2087 ( .A1(a4stg_shl_cnt[0]), .A2(n1409), .A3(n1800), .A4(n1396), 
        .Y(n1422) );
  AO22X1_RVT U2088 ( .A1(a4stg_shl_cnt[0]), .A2(n1398), .A3(n1800), .A4(n1397), 
        .Y(n1424) );
  AO22X1_RVT U2089 ( .A1(a4stg_shl_cnt[1]), .A2(n1422), .A3(n1813), .A4(n1424), 
        .Y(n1442) );
  AO22X1_RVT U2090 ( .A1(a4stg_shl_cnt[0]), .A2(n1400), .A3(n1800), .A4(n1399), 
        .Y(n1423) );
  AO22X1_RVT U2091 ( .A1(a4stg_shl_cnt[0]), .A2(n1402), .A3(n1800), .A4(n1401), 
        .Y(n1426) );
  AO22X1_RVT U2092 ( .A1(a4stg_shl_cnt[1]), .A2(n1423), .A3(n1813), .A4(n1426), 
        .Y(n1443) );
  AO22X1_RVT U2093 ( .A1(a4stg_shl_cnt[2]), .A2(n1442), .A3(n1826), .A4(n1443), 
        .Y(n1475) );
  AO222X1_RVT U2094 ( .A1(n1403), .A2(n1874), .A3(n1444), .A4(n1459), .A5(
        n1475), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[62]) );
  AO22X1_RVT U2095 ( .A1(n1404), .A2(n1877), .A3(n1875), .A4(a4stg_shl[62]), 
        .Y(n1406) );
  AO22X1_RVT U2096 ( .A1(n1919), .A2(n1870), .A3(a4stg_rnd_frac_62), .A4(n2526), .Y(n1405) );
  OR2X1_RVT U2097 ( .A1(n1406), .A2(n1405), .Y(a4stg_rnd_frac_pre2_in[62]) );
  OA221X1_RVT U2098 ( .A1(a4stg_shl_cnt[1]), .A2(n1408), .A3(n1813), .A4(n1407), .A5(n1874), .Y(n1416) );
  AO222X1_RVT U2099 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[14]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[46]), .A5(
        a4stg_shl_data[30]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1421) );
  AO22X1_RVT U2100 ( .A1(a4stg_shl_cnt[0]), .A2(n1421), .A3(n1800), .A4(n1409), 
        .Y(n1433) );
  AO22X1_RVT U2101 ( .A1(a4stg_shl_cnt[1]), .A2(n1433), .A3(n1813), .A4(n1410), 
        .Y(n1450) );
  AO22X1_RVT U2102 ( .A1(a4stg_shl_cnt[1]), .A2(n1412), .A3(n1813), .A4(n1411), 
        .Y(n1451) );
  AO22X1_RVT U2103 ( .A1(a4stg_shl_cnt[2]), .A2(n1450), .A3(n1826), .A4(n1451), 
        .Y(n1482) );
  AO22X1_RVT U2104 ( .A1(a4stg_shl_cnt[1]), .A2(n1414), .A3(n1813), .A4(n1413), 
        .Y(n1452) );
  AO22X1_RVT U2105 ( .A1(a4stg_shl_cnt[3]), .A2(n1482), .A3(n1459), .A4(n1452), 
        .Y(n1415) );
  OR2X1_RVT U2106 ( .A1(n1416), .A2(n1415), .Y(a4stg_shl[61]) );
  AO22X1_RVT U2107 ( .A1(n1875), .A2(a4stg_shl[61]), .A3(n1919), .A4(n1877), 
        .Y(n1418) );
  AO22X1_RVT U2108 ( .A1(n1429), .A2(n1870), .A3(a4stg_rnd_frac_61), .A4(n2526), .Y(n1417) );
  OR2X1_RVT U2109 ( .A1(n1418), .A2(n1417), .Y(a4stg_rnd_frac_pre2_in[61]) );
  OA221X1_RVT U2110 ( .A1(a4stg_shl_cnt[1]), .A2(n1420), .A3(n1813), .A4(n1419), .A5(n1874), .Y(n1428) );
  AO222X1_RVT U2111 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[13]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[45]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[29]), .Y(n1432) );
  AO22X1_RVT U2112 ( .A1(a4stg_shl_cnt[0]), .A2(n1432), .A3(n1800), .A4(n1421), 
        .Y(n1441) );
  AO22X1_RVT U2113 ( .A1(a4stg_shl_cnt[1]), .A2(n1441), .A3(n1813), .A4(n1422), 
        .Y(n1458) );
  AO22X1_RVT U2114 ( .A1(a4stg_shl_cnt[1]), .A2(n1424), .A3(n1813), .A4(n1423), 
        .Y(n1460) );
  AO22X1_RVT U2115 ( .A1(a4stg_shl_cnt[2]), .A2(n1458), .A3(n1826), .A4(n1460), 
        .Y(n1489) );
  AO22X1_RVT U2116 ( .A1(a4stg_shl_cnt[1]), .A2(n1426), .A3(n1813), .A4(n1425), 
        .Y(n1461) );
  AO22X1_RVT U2117 ( .A1(a4stg_shl_cnt[3]), .A2(n1489), .A3(n1459), .A4(n1461), 
        .Y(n1427) );
  OR2X1_RVT U2118 ( .A1(n1428), .A2(n1427), .Y(a4stg_shl[60]) );
  AO22X1_RVT U2119 ( .A1(n1875), .A2(a4stg_shl[60]), .A3(n1429), .A4(n1877), 
        .Y(n1431) );
  AO22X1_RVT U2120 ( .A1(n1437), .A2(n1870), .A3(a4stg_rnd_frac_60), .A4(n2526), .Y(n1430) );
  OR2X1_RVT U2121 ( .A1(n1431), .A2(n1430), .Y(a4stg_rnd_frac_pre2_in[60]) );
  AO222X1_RVT U2122 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[12]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[44]), .A5(
        a4stg_shl_data[28]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1440) );
  AO22X1_RVT U2123 ( .A1(a4stg_shl_cnt[0]), .A2(n1440), .A3(n1800), .A4(n1432), 
        .Y(n1449) );
  AO22X1_RVT U2124 ( .A1(a4stg_shl_cnt[1]), .A2(n1449), .A3(n1813), .A4(n1433), 
        .Y(n1467) );
  AO22X1_RVT U2125 ( .A1(a4stg_shl_cnt[2]), .A2(n1467), .A3(n1826), .A4(n1434), 
        .Y(n1496) );
  AO222X1_RVT U2126 ( .A1(n1436), .A2(n1459), .A3(n1435), .A4(n1874), .A5(
        n1496), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[59]) );
  AO22X1_RVT U2127 ( .A1(n1875), .A2(a4stg_shl[59]), .A3(n1437), .A4(n1877), 
        .Y(n1439) );
  AO22X1_RVT U2128 ( .A1(n1445), .A2(n1870), .A3(a4stg_rnd_frac_59), .A4(n2526), .Y(n1438) );
  OR2X1_RVT U2129 ( .A1(n1439), .A2(n1438), .Y(a4stg_rnd_frac_pre2_in[59]) );
  AO222X1_RVT U2130 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[11]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[43]), .A5(
        a4stg_shl_data[27]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1448) );
  AO22X1_RVT U2131 ( .A1(a4stg_shl_cnt[0]), .A2(n1448), .A3(n1800), .A4(n1440), 
        .Y(n1457) );
  AO22X1_RVT U2132 ( .A1(a4stg_shl_cnt[1]), .A2(n1457), .A3(n1813), .A4(n1441), 
        .Y(n1474) );
  AO22X1_RVT U2133 ( .A1(a4stg_shl_cnt[2]), .A2(n1474), .A3(n1826), .A4(n1442), 
        .Y(n1503) );
  AO222X1_RVT U2134 ( .A1(n1444), .A2(n1874), .A3(n1443), .A4(n1459), .A5(
        n1503), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[58]) );
  AO22X1_RVT U2135 ( .A1(n1875), .A2(a4stg_shl[58]), .A3(n1445), .A4(n1877), 
        .Y(n1447) );
  AO22X1_RVT U2136 ( .A1(n1453), .A2(n1870), .A3(a4stg_rnd_frac_58), .A4(n2526), .Y(n1446) );
  OR2X1_RVT U2137 ( .A1(n1447), .A2(n1446), .Y(a4stg_rnd_frac_pre2_in[58]) );
  AO222X1_RVT U2138 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[10]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[42]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[26]), .Y(n1456) );
  AO22X1_RVT U2139 ( .A1(a4stg_shl_cnt[0]), .A2(n1456), .A3(n1800), .A4(n1448), 
        .Y(n1466) );
  AO22X1_RVT U2140 ( .A1(a4stg_shl_cnt[1]), .A2(n1466), .A3(n1813), .A4(n1449), 
        .Y(n1481) );
  AO22X1_RVT U2141 ( .A1(a4stg_shl_cnt[2]), .A2(n1481), .A3(n1826), .A4(n1450), 
        .Y(n1510) );
  AO222X1_RVT U2142 ( .A1(n1452), .A2(n1874), .A3(n1451), .A4(n1459), .A5(
        n1510), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[57]) );
  AO22X1_RVT U2143 ( .A1(n1875), .A2(a4stg_shl[57]), .A3(n1453), .A4(n1877), 
        .Y(n1455) );
  AO22X1_RVT U2144 ( .A1(n1462), .A2(n1870), .A3(a4stg_rnd_frac_57), .A4(n2526), .Y(n1454) );
  OR2X1_RVT U2145 ( .A1(n1455), .A2(n1454), .Y(a4stg_rnd_frac_pre2_in[57]) );
  AO222X1_RVT U2146 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[9]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[41]), .A5(
        a4stg_shl_data[25]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1465) );
  AO22X1_RVT U2147 ( .A1(a4stg_shl_cnt[0]), .A2(n1465), .A3(n1800), .A4(n1456), 
        .Y(n1473) );
  AO22X1_RVT U2148 ( .A1(a4stg_shl_cnt[1]), .A2(n1473), .A3(n1813), .A4(n1457), 
        .Y(n1488) );
  AO22X1_RVT U2149 ( .A1(a4stg_shl_cnt[2]), .A2(n1488), .A3(n1826), .A4(n1458), 
        .Y(n1517) );
  AO222X1_RVT U2150 ( .A1(n1461), .A2(n1874), .A3(n1460), .A4(n1459), .A5(
        n1517), .A6(a4stg_shl_cnt[3]), .Y(a4stg_shl[56]) );
  AO22X1_RVT U2151 ( .A1(n1875), .A2(a4stg_shl[56]), .A3(n1462), .A4(n1877), 
        .Y(n1464) );
  AO22X1_RVT U2152 ( .A1(n1469), .A2(n1870), .A3(a4stg_rnd_frac_56), .A4(n2526), .Y(n1463) );
  OR2X1_RVT U2153 ( .A1(n1464), .A2(n1463), .Y(a4stg_rnd_frac_pre2_in[56]) );
  AO222X1_RVT U2154 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[8]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[40]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[24]), .Y(n1472) );
  AO22X1_RVT U2155 ( .A1(a4stg_shl_cnt[0]), .A2(n1472), .A3(n1800), .A4(n1465), 
        .Y(n1480) );
  AO22X1_RVT U2156 ( .A1(a4stg_shl_cnt[1]), .A2(n1480), .A3(n1813), .A4(n1466), 
        .Y(n1495) );
  AO22X1_RVT U2157 ( .A1(a4stg_shl_cnt[2]), .A2(n1495), .A3(n1826), .A4(n1467), 
        .Y(n1524) );
  AO22X1_RVT U2158 ( .A1(a4stg_shl_cnt[3]), .A2(n1524), .A3(n1546), .A4(n1468), 
        .Y(a4stg_shl[55]) );
  AO22X1_RVT U2159 ( .A1(n1875), .A2(a4stg_shl[55]), .A3(n1469), .A4(n1877), 
        .Y(n1471) );
  AO22X1_RVT U2160 ( .A1(n1476), .A2(n1870), .A3(a4stg_rnd_frac_55), .A4(n2526), .Y(n1470) );
  OR2X1_RVT U2161 ( .A1(n1471), .A2(n1470), .Y(a4stg_rnd_frac_pre2_in[55]) );
  AO222X1_RVT U2162 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[7]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[39]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[23]), .Y(n1479) );
  AO22X1_RVT U2163 ( .A1(a4stg_shl_cnt[0]), .A2(n1479), .A3(n1800), .A4(n1472), 
        .Y(n1487) );
  AO22X1_RVT U2164 ( .A1(a4stg_shl_cnt[1]), .A2(n1487), .A3(n1813), .A4(n1473), 
        .Y(n1502) );
  AO22X1_RVT U2165 ( .A1(a4stg_shl_cnt[2]), .A2(n1502), .A3(n1826), .A4(n1474), 
        .Y(n1531) );
  AO22X1_RVT U2166 ( .A1(a4stg_shl_cnt[3]), .A2(n1531), .A3(n1546), .A4(n1475), 
        .Y(a4stg_shl[54]) );
  AO22X1_RVT U2167 ( .A1(n1875), .A2(a4stg_shl[54]), .A3(n1476), .A4(n1877), 
        .Y(n1478) );
  AO22X1_RVT U2168 ( .A1(n1483), .A2(n1870), .A3(a4stg_rnd_frac_54), .A4(n2526), .Y(n1477) );
  OR2X1_RVT U2169 ( .A1(n1478), .A2(n1477), .Y(a4stg_rnd_frac_pre2_in[54]) );
  AO222X1_RVT U2170 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[6]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[38]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[22]), .Y(n1486) );
  AO22X1_RVT U2171 ( .A1(a4stg_shl_cnt[0]), .A2(n1486), .A3(n1800), .A4(n1479), 
        .Y(n1494) );
  AO22X1_RVT U2172 ( .A1(a4stg_shl_cnt[1]), .A2(n1494), .A3(n1813), .A4(n1480), 
        .Y(n1509) );
  AO22X1_RVT U2173 ( .A1(a4stg_shl_cnt[2]), .A2(n1509), .A3(n1826), .A4(n1481), 
        .Y(n1538) );
  AO22X1_RVT U2174 ( .A1(a4stg_shl_cnt[3]), .A2(n1538), .A3(n1546), .A4(n1482), 
        .Y(a4stg_shl[53]) );
  AO22X1_RVT U2175 ( .A1(n1875), .A2(a4stg_shl[53]), .A3(n1483), .A4(n1877), 
        .Y(n1485) );
  AO22X1_RVT U2176 ( .A1(n1490), .A2(n1870), .A3(a4stg_rnd_frac_53), .A4(n2526), .Y(n1484) );
  OR2X1_RVT U2177 ( .A1(n1485), .A2(n1484), .Y(a4stg_rnd_frac_pre2_in[53]) );
  AO222X1_RVT U2178 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[5]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[37]), .A5(
        a4stg_shl_data[21]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1493) );
  AO22X1_RVT U2179 ( .A1(a4stg_shl_cnt[0]), .A2(n1493), .A3(n1800), .A4(n1486), 
        .Y(n1501) );
  AO22X1_RVT U2180 ( .A1(a4stg_shl_cnt[1]), .A2(n1501), .A3(n1813), .A4(n1487), 
        .Y(n1516) );
  AO22X1_RVT U2181 ( .A1(a4stg_shl_cnt[2]), .A2(n1516), .A3(n1826), .A4(n1488), 
        .Y(n1545) );
  AO22X1_RVT U2182 ( .A1(a4stg_shl_cnt[3]), .A2(n1545), .A3(n1546), .A4(n1489), 
        .Y(a4stg_shl[52]) );
  AO22X1_RVT U2183 ( .A1(n1875), .A2(a4stg_shl[52]), .A3(n1490), .A4(n1877), 
        .Y(n1492) );
  AO22X1_RVT U2184 ( .A1(n1497), .A2(n1870), .A3(a4stg_rnd_frac_52), .A4(n2526), .Y(n1491) );
  OR2X1_RVT U2185 ( .A1(n1492), .A2(n1491), .Y(a4stg_rnd_frac_pre2_in[52]) );
  AO222X1_RVT U2186 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[4]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[36]), .A5(
        a4stg_shl_data[20]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1500) );
  AO22X1_RVT U2187 ( .A1(a4stg_shl_cnt[0]), .A2(n1500), .A3(n1800), .A4(n1493), 
        .Y(n1508) );
  AO22X1_RVT U2188 ( .A1(a4stg_shl_cnt[1]), .A2(n1508), .A3(n1813), .A4(n1494), 
        .Y(n1523) );
  AO22X1_RVT U2189 ( .A1(a4stg_shl_cnt[2]), .A2(n1523), .A3(n1826), .A4(n1495), 
        .Y(n1553) );
  AO22X1_RVT U2190 ( .A1(a4stg_shl_cnt[3]), .A2(n1553), .A3(n1546), .A4(n1496), 
        .Y(a4stg_shl[51]) );
  AO22X1_RVT U2191 ( .A1(n1875), .A2(a4stg_shl[51]), .A3(n1497), .A4(n1877), 
        .Y(n1499) );
  AO22X1_RVT U2192 ( .A1(n1504), .A2(n1870), .A3(a4stg_rnd_frac_51), .A4(n2526), .Y(n1498) );
  OR2X1_RVT U2193 ( .A1(n1499), .A2(n1498), .Y(a4stg_rnd_frac_pre2_in[51]) );
  AO222X1_RVT U2194 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[3]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[35]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[19]), .Y(n1507) );
  AO22X1_RVT U2195 ( .A1(a4stg_shl_cnt[0]), .A2(n1507), .A3(n1800), .A4(n1500), 
        .Y(n1515) );
  AO22X1_RVT U2196 ( .A1(a4stg_shl_cnt[1]), .A2(n1515), .A3(n1813), .A4(n1501), 
        .Y(n1530) );
  AO22X1_RVT U2197 ( .A1(a4stg_shl_cnt[2]), .A2(n1530), .A3(n1826), .A4(n1502), 
        .Y(n1560) );
  AO22X1_RVT U2198 ( .A1(a4stg_shl_cnt[3]), .A2(n1560), .A3(n1546), .A4(n1503), 
        .Y(a4stg_shl[50]) );
  AO22X1_RVT U2199 ( .A1(n1875), .A2(a4stg_shl[50]), .A3(n1504), .A4(n1877), 
        .Y(n1506) );
  AO22X1_RVT U2200 ( .A1(n1511), .A2(n1870), .A3(a4stg_rnd_frac_50), .A4(n2526), .Y(n1505) );
  OR2X1_RVT U2201 ( .A1(n1506), .A2(n1505), .Y(a4stg_rnd_frac_pre2_in[50]) );
  AO222X1_RVT U2202 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[2]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[34]), .A5(
        a4stg_shl_cnt_dec54_1[0]), .A6(a4stg_shl_data[18]), .Y(n1514) );
  AO22X1_RVT U2203 ( .A1(a4stg_shl_cnt[0]), .A2(n1514), .A3(n1800), .A4(n1507), 
        .Y(n1522) );
  AO22X1_RVT U2204 ( .A1(a4stg_shl_cnt[1]), .A2(n1522), .A3(n1813), .A4(n1508), 
        .Y(n1537) );
  AO22X1_RVT U2205 ( .A1(a4stg_shl_cnt[2]), .A2(n1537), .A3(n1826), .A4(n1509), 
        .Y(n1567) );
  AO22X1_RVT U2206 ( .A1(a4stg_shl_cnt[3]), .A2(n1567), .A3(n1546), .A4(n1510), 
        .Y(a4stg_shl[49]) );
  AO22X1_RVT U2207 ( .A1(n1875), .A2(a4stg_shl[49]), .A3(n1511), .A4(n1877), 
        .Y(n1513) );
  AO22X1_RVT U2208 ( .A1(n1518), .A2(n1870), .A3(a4stg_rnd_frac_49), .A4(n2526), .Y(n1512) );
  OR2X1_RVT U2209 ( .A1(n1513), .A2(n1512), .Y(a4stg_rnd_frac_pre2_in[49]) );
  AO222X1_RVT U2210 ( .A1(\a4stg_shl_cnt_dec54_2[0] ), .A2(a4stg_shl_data[1]), 
        .A3(a4stg_shl_cnt_dec54_0[0]), .A4(a4stg_shl_data[33]), .A5(
        a4stg_shl_data[17]), .A6(a4stg_shl_cnt_dec54_1[0]), .Y(n1521) );
  AO22X1_RVT U2211 ( .A1(a4stg_shl_cnt[0]), .A2(n1521), .A3(n1800), .A4(n1514), 
        .Y(n1529) );
  AO22X1_RVT U2212 ( .A1(a4stg_shl_cnt[1]), .A2(n1529), .A3(n1813), .A4(n1515), 
        .Y(n1544) );
  AO22X1_RVT U2213 ( .A1(a4stg_shl_cnt[2]), .A2(n1544), .A3(n1826), .A4(n1516), 
        .Y(n1574) );
  AO22X1_RVT U2214 ( .A1(a4stg_shl_cnt[3]), .A2(n1574), .A3(n1546), .A4(n1517), 
        .Y(a4stg_shl[48]) );
  AO22X1_RVT U2215 ( .A1(n1875), .A2(a4stg_shl[48]), .A3(n1518), .A4(n1877), 
        .Y(n1520) );
  AO22X1_RVT U2216 ( .A1(n1525), .A2(n1870), .A3(a4stg_rnd_frac_48), .A4(n2526), .Y(n1519) );
  OR2X1_RVT U2217 ( .A1(n1520), .A2(n1519), .Y(a4stg_rnd_frac_pre2_in[48]) );
  AO222X1_RVT U2218 ( .A1(a4stg_shl_data[16]), .A2(a4stg_shl_cnt_dec54_1[0]), 
        .A3(a4stg_shl_data[0]), .A4(\a4stg_shl_cnt_dec54_2[0] ), .A5(
        a4stg_shl_data[32]), .A6(a4stg_shl_cnt_dec54_0[0]), .Y(n1528) );
  AO22X1_RVT U2219 ( .A1(a4stg_shl_cnt[0]), .A2(n1528), .A3(n1800), .A4(n1521), 
        .Y(n1536) );
  AO22X1_RVT U2220 ( .A1(a4stg_shl_cnt[1]), .A2(n1536), .A3(n1813), .A4(n1522), 
        .Y(n1552) );
  AO22X1_RVT U2221 ( .A1(a4stg_shl_cnt[2]), .A2(n1552), .A3(n1826), .A4(n1523), 
        .Y(n1581) );
  AO22X1_RVT U2222 ( .A1(a4stg_shl_cnt[3]), .A2(n1581), .A3(n1546), .A4(n1524), 
        .Y(a4stg_shl[47]) );
  AO22X1_RVT U2223 ( .A1(n1875), .A2(a4stg_shl[47]), .A3(n1525), .A4(n1877), 
        .Y(n1527) );
  AO22X1_RVT U2224 ( .A1(n1532), .A2(n1870), .A3(a4stg_rnd_frac_47), .A4(n2526), .Y(n1526) );
  OR2X1_RVT U2225 ( .A1(n1527), .A2(n1526), .Y(a4stg_rnd_frac_pre2_in[47]) );
  AO22X1_RVT U2226 ( .A1(a4stg_shl_data[31]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[15]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1535) );
  AO22X1_RVT U2227 ( .A1(a4stg_shl_cnt[0]), .A2(n1535), .A3(n1800), .A4(n1528), 
        .Y(n1543) );
  AO22X1_RVT U2228 ( .A1(a4stg_shl_cnt[1]), .A2(n1543), .A3(n1813), .A4(n1529), 
        .Y(n1559) );
  AO22X1_RVT U2229 ( .A1(a4stg_shl_cnt[2]), .A2(n1559), .A3(n1826), .A4(n1530), 
        .Y(n1588) );
  AO22X1_RVT U2230 ( .A1(a4stg_shl_cnt[3]), .A2(n1588), .A3(n1546), .A4(n1531), 
        .Y(a4stg_shl[46]) );
  AO22X1_RVT U2231 ( .A1(n1875), .A2(a4stg_shl[46]), .A3(n1532), .A4(n1877), 
        .Y(n1534) );
  AO22X1_RVT U2232 ( .A1(n1539), .A2(n1870), .A3(a4stg_rnd_frac_46), .A4(n2526), .Y(n1533) );
  OR2X1_RVT U2233 ( .A1(n1534), .A2(n1533), .Y(a4stg_rnd_frac_pre2_in[46]) );
  AO22X1_RVT U2234 ( .A1(a4stg_shl_data[14]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[30]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1542) );
  AO22X1_RVT U2235 ( .A1(a4stg_shl_cnt[0]), .A2(n1542), .A3(n1800), .A4(n1535), 
        .Y(n1551) );
  AO22X1_RVT U2236 ( .A1(a4stg_shl_cnt[1]), .A2(n1551), .A3(n1813), .A4(n1536), 
        .Y(n1566) );
  AO22X1_RVT U2237 ( .A1(a4stg_shl_cnt[2]), .A2(n1566), .A3(n1826), .A4(n1537), 
        .Y(n1595) );
  AO22X1_RVT U2238 ( .A1(a4stg_shl_cnt[3]), .A2(n1595), .A3(n1546), .A4(n1538), 
        .Y(a4stg_shl[45]) );
  AO22X1_RVT U2239 ( .A1(n1875), .A2(a4stg_shl[45]), .A3(n1539), .A4(n1877), 
        .Y(n1541) );
  AO22X1_RVT U2240 ( .A1(n1547), .A2(n1870), .A3(a4stg_rnd_frac_45), .A4(n2526), .Y(n1540) );
  OR2X1_RVT U2241 ( .A1(n1541), .A2(n1540), .Y(a4stg_rnd_frac_pre2_in[45]) );
  AO22X1_RVT U2242 ( .A1(a4stg_shl_data[13]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[29]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1550) );
  AO22X1_RVT U2243 ( .A1(a4stg_shl_cnt[0]), .A2(n1550), .A3(n1800), .A4(n1542), 
        .Y(n1558) );
  AO22X1_RVT U2244 ( .A1(a4stg_shl_cnt[1]), .A2(n1558), .A3(n1813), .A4(n1543), 
        .Y(n1573) );
  AO22X1_RVT U2245 ( .A1(a4stg_shl_cnt[2]), .A2(n1573), .A3(n1826), .A4(n1544), 
        .Y(n1602) );
  AO22X1_RVT U2246 ( .A1(a4stg_shl_cnt[3]), .A2(n1602), .A3(n1546), .A4(n1545), 
        .Y(a4stg_shl[44]) );
  AO22X1_RVT U2247 ( .A1(n1875), .A2(a4stg_shl[44]), .A3(n1547), .A4(n1877), 
        .Y(n1549) );
  AO22X1_RVT U2248 ( .A1(n1554), .A2(n1870), .A3(a4stg_rnd_frac_44), .A4(n2526), .Y(n1548) );
  OR2X1_RVT U2249 ( .A1(n1549), .A2(n1548), .Y(a4stg_rnd_frac_pre2_in[44]) );
  AO22X1_RVT U2250 ( .A1(a4stg_shl_data[28]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[12]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1557) );
  AO22X1_RVT U2251 ( .A1(a4stg_shl_cnt[0]), .A2(n1557), .A3(n1800), .A4(n1550), 
        .Y(n1565) );
  AO22X1_RVT U2252 ( .A1(a4stg_shl_cnt[1]), .A2(n1565), .A3(n1813), .A4(n1551), 
        .Y(n1580) );
  AO22X1_RVT U2253 ( .A1(a4stg_shl_cnt[2]), .A2(n1580), .A3(n1826), .A4(n1552), 
        .Y(n1609) );
  AO22X1_RVT U2254 ( .A1(a4stg_shl_cnt[3]), .A2(n1609), .A3(n1546), .A4(n1553), 
        .Y(a4stg_shl[43]) );
  AO22X1_RVT U2255 ( .A1(n1875), .A2(a4stg_shl[43]), .A3(n1554), .A4(n1877), 
        .Y(n1556) );
  AO22X1_RVT U2256 ( .A1(n1561), .A2(n1870), .A3(a4stg_rnd_frac_43), .A4(n2526), .Y(n1555) );
  OR2X1_RVT U2257 ( .A1(n1556), .A2(n1555), .Y(a4stg_rnd_frac_pre2_in[43]) );
  AO22X1_RVT U2258 ( .A1(a4stg_shl_data[27]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[11]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1564) );
  AO22X1_RVT U2259 ( .A1(a4stg_shl_cnt[0]), .A2(n1564), .A3(n1800), .A4(n1557), 
        .Y(n1572) );
  AO22X1_RVT U2260 ( .A1(a4stg_shl_cnt[1]), .A2(n1572), .A3(n1813), .A4(n1558), 
        .Y(n1587) );
  AO22X1_RVT U2261 ( .A1(a4stg_shl_cnt[2]), .A2(n1587), .A3(n1826), .A4(n1559), 
        .Y(n1616) );
  AO22X1_RVT U2262 ( .A1(a4stg_shl_cnt[3]), .A2(n1616), .A3(n1546), .A4(n1560), 
        .Y(a4stg_shl[42]) );
  AO22X1_RVT U2263 ( .A1(n1875), .A2(a4stg_shl[42]), .A3(n1561), .A4(n1877), 
        .Y(n1563) );
  AO22X1_RVT U2264 ( .A1(n1568), .A2(n1870), .A3(a4stg_rnd_frac_42), .A4(n2526), .Y(n1562) );
  OR2X1_RVT U2265 ( .A1(n1563), .A2(n1562), .Y(a4stg_rnd_frac_pre2_in[42]) );
  AO22X1_RVT U2266 ( .A1(a4stg_shl_data[10]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[26]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1571) );
  AO22X1_RVT U2267 ( .A1(a4stg_shl_cnt[0]), .A2(n1571), .A3(n1800), .A4(n1564), 
        .Y(n1579) );
  AO22X1_RVT U2268 ( .A1(a4stg_shl_cnt[1]), .A2(n1579), .A3(n1813), .A4(n1565), 
        .Y(n1594) );
  AO22X1_RVT U2269 ( .A1(a4stg_shl_cnt[2]), .A2(n1594), .A3(n1826), .A4(n1566), 
        .Y(n1623) );
  AO22X1_RVT U2270 ( .A1(a4stg_shl_cnt[3]), .A2(n1623), .A3(n1546), .A4(n1567), 
        .Y(a4stg_shl[41]) );
  AO22X1_RVT U2271 ( .A1(n1875), .A2(a4stg_shl[41]), .A3(n1568), .A4(n1877), 
        .Y(n1570) );
  AO22X1_RVT U2272 ( .A1(n1575), .A2(n1870), .A3(a4stg_rnd_frac_41), .A4(n2526), .Y(n1569) );
  OR2X1_RVT U2273 ( .A1(n1570), .A2(n1569), .Y(a4stg_rnd_frac_pre2_in[41]) );
  AO22X1_RVT U2274 ( .A1(a4stg_shl_data[9]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[25]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1578) );
  AO22X1_RVT U2275 ( .A1(a4stg_shl_cnt[0]), .A2(n1578), .A3(n1800), .A4(n1571), 
        .Y(n1586) );
  AO22X1_RVT U2276 ( .A1(a4stg_shl_cnt[1]), .A2(n1586), .A3(n1813), .A4(n1572), 
        .Y(n1601) );
  AO22X1_RVT U2277 ( .A1(a4stg_shl_cnt[2]), .A2(n1601), .A3(n1826), .A4(n1573), 
        .Y(n1630) );
  AO22X1_RVT U2278 ( .A1(a4stg_shl_cnt[3]), .A2(n1630), .A3(n1546), .A4(n1574), 
        .Y(a4stg_shl[40]) );
  AO22X1_RVT U2279 ( .A1(n1875), .A2(a4stg_shl[40]), .A3(n1575), .A4(n1877), 
        .Y(n1577) );
  AO22X1_RVT U2280 ( .A1(n1582), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_40), .Y(n1576) );
  OR2X1_RVT U2281 ( .A1(n1577), .A2(n1576), .Y(a4stg_rnd_frac_pre2_in[40]) );
  AO22X1_RVT U2282 ( .A1(a4stg_shl_data[24]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[8]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1585) );
  AO22X1_RVT U2283 ( .A1(a4stg_shl_cnt[0]), .A2(n1585), .A3(n1800), .A4(n1578), 
        .Y(n1593) );
  AO22X1_RVT U2284 ( .A1(a4stg_shl_cnt[1]), .A2(n1593), .A3(n1813), .A4(n1579), 
        .Y(n1608) );
  AO22X1_RVT U2285 ( .A1(a4stg_shl_cnt[2]), .A2(n1608), .A3(n1826), .A4(n1580), 
        .Y(n1637) );
  AO22X1_RVT U2286 ( .A1(a4stg_shl_cnt[3]), .A2(n1637), .A3(n1546), .A4(n1581), 
        .Y(a4stg_shl[39]) );
  AO22X1_RVT U2287 ( .A1(n1875), .A2(a4stg_shl[39]), .A3(n1582), .A4(n1877), 
        .Y(n1584) );
  AO22X1_RVT U2288 ( .A1(n1589), .A2(n1870), .A3(a4stg_rnd_frac_39), .A4(n2526), .Y(n1583) );
  OR2X1_RVT U2289 ( .A1(n1584), .A2(n1583), .Y(a4stg_rnd_frac_pre2_in[39]) );
  AO22X1_RVT U2290 ( .A1(a4stg_shl_data[7]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[23]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1592) );
  AO22X1_RVT U2291 ( .A1(a4stg_shl_cnt[0]), .A2(n1592), .A3(n1800), .A4(n1585), 
        .Y(n1600) );
  AO22X1_RVT U2292 ( .A1(a4stg_shl_cnt[1]), .A2(n1600), .A3(n1813), .A4(n1586), 
        .Y(n1615) );
  AO22X1_RVT U2293 ( .A1(a4stg_shl_cnt[2]), .A2(n1615), .A3(n1826), .A4(n1587), 
        .Y(n1644) );
  AO22X1_RVT U2294 ( .A1(a4stg_shl_cnt[3]), .A2(n1644), .A3(n1546), .A4(n1588), 
        .Y(a4stg_shl[38]) );
  AO22X1_RVT U2295 ( .A1(n1875), .A2(a4stg_shl[38]), .A3(n1589), .A4(n1877), 
        .Y(n1591) );
  AO22X1_RVT U2296 ( .A1(n1596), .A2(n1870), .A3(a4stg_rnd_frac[38]), .A4(
        n2526), .Y(n1590) );
  OR2X1_RVT U2297 ( .A1(n1591), .A2(n1590), .Y(a4stg_rnd_frac_pre2_in[38]) );
  AO22X1_RVT U2298 ( .A1(a4stg_shl_data[6]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[22]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1599) );
  AO22X1_RVT U2299 ( .A1(a4stg_shl_cnt[0]), .A2(n1599), .A3(n1800), .A4(n1592), 
        .Y(n1607) );
  AO22X1_RVT U2300 ( .A1(a4stg_shl_cnt[1]), .A2(n1607), .A3(n1813), .A4(n1593), 
        .Y(n1622) );
  AO22X1_RVT U2301 ( .A1(a4stg_shl_cnt[2]), .A2(n1622), .A3(n1826), .A4(n1594), 
        .Y(n1650) );
  AO22X1_RVT U2302 ( .A1(a4stg_shl_cnt[3]), .A2(n1650), .A3(n1546), .A4(n1595), 
        .Y(a4stg_shl[37]) );
  AO22X1_RVT U2303 ( .A1(n1875), .A2(a4stg_shl[37]), .A3(n1596), .A4(n1877), 
        .Y(n1598) );
  AO22X1_RVT U2304 ( .A1(n1603), .A2(n1870), .A3(a4stg_rnd_frac[37]), .A4(
        n2526), .Y(n1597) );
  OR2X1_RVT U2305 ( .A1(n1598), .A2(n1597), .Y(a4stg_rnd_frac_pre2_in[37]) );
  AO22X1_RVT U2306 ( .A1(a4stg_shl_data[5]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[21]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1606) );
  AO22X1_RVT U2307 ( .A1(a4stg_shl_cnt[0]), .A2(n1606), .A3(n1800), .A4(n1599), 
        .Y(n1614) );
  AO22X1_RVT U2308 ( .A1(a4stg_shl_cnt[1]), .A2(n1614), .A3(n1813), .A4(n1600), 
        .Y(n1629) );
  AO22X1_RVT U2309 ( .A1(a4stg_shl_cnt[2]), .A2(n1629), .A3(n1826), .A4(n1601), 
        .Y(n1656) );
  AO22X1_RVT U2310 ( .A1(a4stg_shl_cnt[3]), .A2(n1656), .A3(n1546), .A4(n1602), 
        .Y(a4stg_shl[36]) );
  AO22X1_RVT U2311 ( .A1(n1875), .A2(a4stg_shl[36]), .A3(n1603), .A4(n1877), 
        .Y(n1605) );
  AO22X1_RVT U2312 ( .A1(n1610), .A2(n1870), .A3(a4stg_rnd_frac[36]), .A4(
        n2526), .Y(n1604) );
  OR2X1_RVT U2313 ( .A1(n1605), .A2(n1604), .Y(a4stg_rnd_frac_pre2_in[36]) );
  AO22X1_RVT U2314 ( .A1(a4stg_shl_data[20]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[4]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1613) );
  AO22X1_RVT U2315 ( .A1(a4stg_shl_cnt[0]), .A2(n1613), .A3(n1800), .A4(n1606), 
        .Y(n1621) );
  AO22X1_RVT U2316 ( .A1(a4stg_shl_cnt[1]), .A2(n1621), .A3(n1813), .A4(n1607), 
        .Y(n1636) );
  AO22X1_RVT U2317 ( .A1(a4stg_shl_cnt[2]), .A2(n1636), .A3(n1826), .A4(n1608), 
        .Y(n1662) );
  AO22X1_RVT U2318 ( .A1(a4stg_shl_cnt[3]), .A2(n1662), .A3(n1546), .A4(n1609), 
        .Y(a4stg_shl[35]) );
  AO22X1_RVT U2319 ( .A1(n1875), .A2(a4stg_shl[35]), .A3(n1610), .A4(n1877), 
        .Y(n1612) );
  AO22X1_RVT U2320 ( .A1(n1617), .A2(n1870), .A3(a4stg_rnd_frac[35]), .A4(
        n2526), .Y(n1611) );
  OR2X1_RVT U2321 ( .A1(n1612), .A2(n1611), .Y(a4stg_rnd_frac_pre2_in[35]) );
  AO22X1_RVT U2322 ( .A1(a4stg_shl_data[19]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[3]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1620) );
  AO22X1_RVT U2323 ( .A1(a4stg_shl_cnt[0]), .A2(n1620), .A3(n1800), .A4(n1613), 
        .Y(n1628) );
  AO22X1_RVT U2324 ( .A1(a4stg_shl_cnt[1]), .A2(n1628), .A3(n1813), .A4(n1614), 
        .Y(n1643) );
  AO22X1_RVT U2325 ( .A1(a4stg_shl_cnt[2]), .A2(n1643), .A3(n1826), .A4(n1615), 
        .Y(n1733) );
  AO22X1_RVT U2326 ( .A1(a4stg_shl_cnt[3]), .A2(n1733), .A3(n1546), .A4(n1616), 
        .Y(a4stg_shl[34]) );
  AO22X1_RVT U2327 ( .A1(n1875), .A2(a4stg_shl[34]), .A3(n1617), .A4(n1877), 
        .Y(n1619) );
  AO22X1_RVT U2328 ( .A1(n1624), .A2(n1870), .A3(a4stg_rnd_frac[34]), .A4(
        n2526), .Y(n1618) );
  OR2X1_RVT U2329 ( .A1(n1619), .A2(n1618), .Y(a4stg_rnd_frac_pre2_in[34]) );
  AO22X1_RVT U2330 ( .A1(a4stg_shl_data[18]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[2]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1627) );
  AO22X1_RVT U2331 ( .A1(a4stg_shl_cnt[0]), .A2(n1627), .A3(n1800), .A4(n1620), 
        .Y(n1635) );
  AO22X1_RVT U2332 ( .A1(a4stg_shl_cnt[1]), .A2(n1635), .A3(n1813), .A4(n1621), 
        .Y(n1649) );
  AO22X1_RVT U2333 ( .A1(a4stg_shl_cnt[2]), .A2(n1649), .A3(n1826), .A4(n1622), 
        .Y(n1741) );
  AO22X1_RVT U2334 ( .A1(a4stg_shl_cnt[3]), .A2(n1741), .A3(n1546), .A4(n1623), 
        .Y(a4stg_shl[33]) );
  AO22X1_RVT U2335 ( .A1(n1875), .A2(a4stg_shl[33]), .A3(n1624), .A4(n1877), 
        .Y(n1626) );
  AO22X1_RVT U2336 ( .A1(n1631), .A2(n1870), .A3(a4stg_rnd_frac[33]), .A4(
        n2526), .Y(n1625) );
  OR2X1_RVT U2337 ( .A1(n1626), .A2(n1625), .Y(a4stg_rnd_frac_pre2_in[33]) );
  AO22X1_RVT U2338 ( .A1(a4stg_shl_data[1]), .A2(a4stg_shl_cnt_dec54_1[1]), 
        .A3(a4stg_shl_data[17]), .A4(a4stg_shl_cnt_dec54_0[1]), .Y(n1634) );
  AO22X1_RVT U2339 ( .A1(a4stg_shl_cnt[0]), .A2(n1634), .A3(n1800), .A4(n1627), 
        .Y(n1642) );
  AO22X1_RVT U2340 ( .A1(a4stg_shl_cnt[1]), .A2(n1642), .A3(n1813), .A4(n1628), 
        .Y(n1655) );
  AO22X1_RVT U2341 ( .A1(a4stg_shl_cnt[2]), .A2(n1655), .A3(n1826), .A4(n1629), 
        .Y(n1747) );
  AO22X1_RVT U2342 ( .A1(a4stg_shl_cnt[3]), .A2(n1747), .A3(n1546), .A4(n1630), 
        .Y(a4stg_shl[32]) );
  AO22X1_RVT U2343 ( .A1(n1875), .A2(a4stg_shl[32]), .A3(n1631), .A4(n1877), 
        .Y(n1633) );
  AO22X1_RVT U2344 ( .A1(n1638), .A2(n1870), .A3(a4stg_rnd_frac[32]), .A4(
        n2526), .Y(n1632) );
  OR2X1_RVT U2345 ( .A1(n1633), .A2(n1632), .Y(a4stg_rnd_frac_pre2_in[32]) );
  AO22X1_RVT U2346 ( .A1(a4stg_shl_data[16]), .A2(a4stg_shl_cnt_dec54_0[1]), 
        .A3(a4stg_shl_data[0]), .A4(a4stg_shl_cnt_dec54_1[1]), .Y(n1641) );
  AO22X1_RVT U2347 ( .A1(a4stg_shl_cnt[0]), .A2(n1641), .A3(n1800), .A4(n1634), 
        .Y(n1648) );
  AO22X1_RVT U2348 ( .A1(a4stg_shl_cnt[1]), .A2(n1648), .A3(n1813), .A4(n1635), 
        .Y(n1661) );
  AO22X1_RVT U2349 ( .A1(a4stg_shl_cnt[2]), .A2(n1661), .A3(n1826), .A4(n1636), 
        .Y(n1753) );
  AO22X1_RVT U2350 ( .A1(a4stg_shl_cnt[3]), .A2(n1753), .A3(n1546), .A4(n1637), 
        .Y(a4stg_shl[31]) );
  AO22X1_RVT U2351 ( .A1(n1875), .A2(a4stg_shl[31]), .A3(n1638), .A4(n1877), 
        .Y(n1640) );
  AO22X1_RVT U2352 ( .A1(n1645), .A2(n1870), .A3(a4stg_rnd_frac[31]), .A4(
        n2526), .Y(n1639) );
  OR2X1_RVT U2353 ( .A1(n1640), .A2(n1639), .Y(a4stg_rnd_frac_pre2_in[31]) );
  AND2X1_RVT U2354 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_cnt_dec54_0[1]), .Y(
        n1666) );
  AO22X1_RVT U2355 ( .A1(n1666), .A2(a4stg_shl_data[15]), .A3(n1800), .A4(
        n1641), .Y(n1654) );
  AO22X1_RVT U2356 ( .A1(a4stg_shl_cnt[1]), .A2(n1654), .A3(n1813), .A4(n1642), 
        .Y(n1732) );
  AO22X1_RVT U2357 ( .A1(a4stg_shl_cnt[2]), .A2(n1732), .A3(n1826), .A4(n1643), 
        .Y(n1759) );
  AO22X1_RVT U2358 ( .A1(a4stg_shl_cnt[3]), .A2(n1759), .A3(n1546), .A4(n1644), 
        .Y(a4stg_shl[30]) );
  AO22X1_RVT U2359 ( .A1(n1875), .A2(a4stg_shl[30]), .A3(n1645), .A4(n1877), 
        .Y(n1647) );
  AO22X1_RVT U2360 ( .A1(n1651), .A2(n1870), .A3(a4stg_rnd_frac[30]), .A4(
        n2526), .Y(n1646) );
  OR2X1_RVT U2361 ( .A1(n1647), .A2(n1646), .Y(a4stg_rnd_frac_pre2_in[30]) );
  AND2X1_RVT U2362 ( .A1(a4stg_shl_cnt_dec54_0[1]), .A2(n1800), .Y(n1737) );
  AO22X1_RVT U2363 ( .A1(a4stg_shl_data[14]), .A2(n1666), .A3(
        a4stg_shl_data[15]), .A4(n1737), .Y(n1660) );
  AO22X1_RVT U2364 ( .A1(a4stg_shl_cnt[1]), .A2(n1660), .A3(n1813), .A4(n1648), 
        .Y(n1740) );
  AO22X1_RVT U2365 ( .A1(a4stg_shl_cnt[2]), .A2(n1740), .A3(n1826), .A4(n1649), 
        .Y(n1765) );
  AO22X1_RVT U2366 ( .A1(a4stg_shl_cnt[3]), .A2(n1765), .A3(n1546), .A4(n1650), 
        .Y(a4stg_shl[29]) );
  AO22X1_RVT U2367 ( .A1(n1875), .A2(a4stg_shl[29]), .A3(n1651), .A4(n1877), 
        .Y(n1653) );
  AO22X1_RVT U2368 ( .A1(n1657), .A2(n1870), .A3(a4stg_rnd_frac[29]), .A4(
        n2526), .Y(n1652) );
  OR2X1_RVT U2369 ( .A1(n1653), .A2(n1652), .Y(a4stg_rnd_frac_pre2_in[29]) );
  AO22X1_RVT U2370 ( .A1(a4stg_shl_data[13]), .A2(n1666), .A3(
        a4stg_shl_data[14]), .A4(n1737), .Y(n1667) );
  AO22X1_RVT U2371 ( .A1(a4stg_shl_cnt[1]), .A2(n1667), .A3(n1813), .A4(n1654), 
        .Y(n1746) );
  AO22X1_RVT U2372 ( .A1(a4stg_shl_cnt[2]), .A2(n1746), .A3(n1826), .A4(n1655), 
        .Y(n1771) );
  AO22X1_RVT U2373 ( .A1(a4stg_shl_cnt[3]), .A2(n1771), .A3(n1546), .A4(n1656), 
        .Y(a4stg_shl[28]) );
  AO22X1_RVT U2374 ( .A1(n1875), .A2(a4stg_shl[28]), .A3(n1657), .A4(n1877), 
        .Y(n1659) );
  AO22X1_RVT U2375 ( .A1(n1663), .A2(n1870), .A3(a4stg_rnd_frac[28]), .A4(
        n2526), .Y(n1658) );
  OR2X1_RVT U2376 ( .A1(n1659), .A2(n1658), .Y(a4stg_rnd_frac_pre2_in[28]) );
  AO22X1_RVT U2377 ( .A1(a4stg_shl_data[12]), .A2(n1666), .A3(
        a4stg_shl_data[13]), .A4(n1737), .Y(n1739) );
  AO22X1_RVT U2378 ( .A1(a4stg_shl_cnt[1]), .A2(n1739), .A3(n1813), .A4(n1660), 
        .Y(n1752) );
  AO22X1_RVT U2379 ( .A1(a4stg_shl_cnt[2]), .A2(n1752), .A3(n1826), .A4(n1661), 
        .Y(n1777) );
  AO22X1_RVT U2380 ( .A1(a4stg_shl_cnt[3]), .A2(n1777), .A3(n1546), .A4(n1662), 
        .Y(a4stg_shl[27]) );
  AO22X1_RVT U2381 ( .A1(n1875), .A2(a4stg_shl[27]), .A3(n1663), .A4(n1877), 
        .Y(n1665) );
  AO22X1_RVT U2382 ( .A1(n1734), .A2(n1870), .A3(a4stg_rnd_frac[27]), .A4(
        n2526), .Y(n1664) );
  OR2X1_RVT U2383 ( .A1(n1665), .A2(n1664), .Y(a4stg_rnd_frac_pre2_in[27]) );
  AO22X1_RVT U2384 ( .A1(a4stg_shl_data[12]), .A2(n1737), .A3(
        a4stg_shl_data[11]), .A4(n1666), .Y(n1745) );
  AO22X1_RVT U2385 ( .A1(a4stg_shl_cnt[1]), .A2(n1745), .A3(n1813), .A4(n1667), 
        .Y(n1758) );
  AO22X1_RVT U2386 ( .A1(a4stg_shl_cnt[2]), .A2(n1758), .A3(n1826), .A4(n1732), 
        .Y(n1783) );
  AO22X1_RVT U2387 ( .A1(a4stg_shl_cnt[3]), .A2(n1783), .A3(n1546), .A4(n1733), 
        .Y(a4stg_shl[26]) );
  AO22X1_RVT U2388 ( .A1(n1875), .A2(a4stg_shl[26]), .A3(n1734), .A4(n1877), 
        .Y(n1736) );
  AO22X1_RVT U2389 ( .A1(n1742), .A2(n1870), .A3(a4stg_rnd_frac[26]), .A4(
        n2526), .Y(n1735) );
  OR2X1_RVT U2390 ( .A1(n1736), .A2(n1735), .Y(a4stg_rnd_frac_pre2_in[26]) );
  AND2X1_RVT U2391 ( .A1(a4stg_shl_data[10]), .A2(a4stg_shl_cnt_dec54_0[2]), 
        .Y(n1738) );
  AO22X1_RVT U2392 ( .A1(a4stg_shl_cnt[0]), .A2(n1738), .A3(a4stg_shl_data[11]), .A4(n1737), .Y(n1751) );
  AO22X1_RVT U2393 ( .A1(a4stg_shl_cnt[1]), .A2(n1751), .A3(n1813), .A4(n1739), 
        .Y(n1764) );
  AO22X1_RVT U2394 ( .A1(a4stg_shl_cnt[2]), .A2(n1764), .A3(n1826), .A4(n1740), 
        .Y(n1789) );
  AO22X1_RVT U2395 ( .A1(a4stg_shl_cnt[3]), .A2(n1789), .A3(n1546), .A4(n1741), 
        .Y(a4stg_shl[25]) );
  AO22X1_RVT U2396 ( .A1(n1875), .A2(a4stg_shl[25]), .A3(n1742), .A4(n1877), 
        .Y(n1744) );
  AO22X1_RVT U2397 ( .A1(n1748), .A2(n1870), .A3(a4stg_rnd_frac[25]), .A4(
        n2526), .Y(n1743) );
  OR2X1_RVT U2398 ( .A1(n1744), .A2(n1743), .Y(a4stg_rnd_frac_pre2_in[25]) );
  OA221X1_RVT U2399 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[10]), .A3(
        n1800), .A4(a4stg_shl_data[9]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(
        n1757) );
  AO22X1_RVT U2400 ( .A1(a4stg_shl_cnt[1]), .A2(n1757), .A3(n1813), .A4(n1745), 
        .Y(n1770) );
  AO22X1_RVT U2401 ( .A1(a4stg_shl_cnt[2]), .A2(n1770), .A3(n1826), .A4(n1746), 
        .Y(n1796) );
  AO22X1_RVT U2402 ( .A1(a4stg_shl_cnt[3]), .A2(n1796), .A3(n1546), .A4(n1747), 
        .Y(a4stg_shl[24]) );
  AO22X1_RVT U2403 ( .A1(n1875), .A2(a4stg_shl[24]), .A3(n1748), .A4(n1877), 
        .Y(n1750) );
  AO22X1_RVT U2404 ( .A1(n1754), .A2(n1870), .A3(a4stg_rnd_frac[24]), .A4(
        n2526), .Y(n1749) );
  OR2X1_RVT U2405 ( .A1(n1750), .A2(n1749), .Y(a4stg_rnd_frac_pre2_in[24]) );
  OA221X1_RVT U2406 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[9]), .A3(n1800), .A4(a4stg_shl_data[8]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1763) );
  AO22X1_RVT U2407 ( .A1(a4stg_shl_cnt[1]), .A2(n1763), .A3(n1813), .A4(n1751), 
        .Y(n1776) );
  AO22X1_RVT U2408 ( .A1(a4stg_shl_cnt[2]), .A2(n1776), .A3(n1826), .A4(n1752), 
        .Y(n1803) );
  AO22X1_RVT U2409 ( .A1(a4stg_shl_cnt[3]), .A2(n1803), .A3(n1546), .A4(n1753), 
        .Y(a4stg_shl[23]) );
  AO22X1_RVT U2410 ( .A1(n1875), .A2(a4stg_shl[23]), .A3(n1754), .A4(n1877), 
        .Y(n1756) );
  AO22X1_RVT U2411 ( .A1(n1760), .A2(n1870), .A3(a4stg_rnd_frac[23]), .A4(
        n2526), .Y(n1755) );
  OR2X1_RVT U2412 ( .A1(n1756), .A2(n1755), .Y(a4stg_rnd_frac_pre2_in[23]) );
  OA221X1_RVT U2413 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[8]), .A3(n1800), .A4(a4stg_shl_data[7]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1769) );
  AO22X1_RVT U2414 ( .A1(a4stg_shl_cnt[1]), .A2(n1769), .A3(n1813), .A4(n1757), 
        .Y(n1782) );
  AO22X1_RVT U2415 ( .A1(a4stg_shl_cnt[2]), .A2(n1782), .A3(n1826), .A4(n1758), 
        .Y(n1808) );
  AO22X1_RVT U2416 ( .A1(a4stg_shl_cnt[3]), .A2(n1808), .A3(n1546), .A4(n1759), 
        .Y(a4stg_shl[22]) );
  AO22X1_RVT U2417 ( .A1(n1875), .A2(a4stg_shl[22]), .A3(n1760), .A4(n1877), 
        .Y(n1762) );
  AO22X1_RVT U2418 ( .A1(n1766), .A2(n1870), .A3(a4stg_rnd_frac[22]), .A4(
        n2526), .Y(n1761) );
  OR2X1_RVT U2419 ( .A1(n1762), .A2(n1761), .Y(a4stg_rnd_frac_pre2_in[22]) );
  OA221X1_RVT U2420 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[7]), .A3(n1800), .A4(a4stg_shl_data[6]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1775) );
  AO22X1_RVT U2421 ( .A1(a4stg_shl_cnt[1]), .A2(n1775), .A3(n1813), .A4(n1763), 
        .Y(n1788) );
  AO22X1_RVT U2422 ( .A1(a4stg_shl_cnt[2]), .A2(n1788), .A3(n1826), .A4(n1764), 
        .Y(n1815) );
  AO22X1_RVT U2423 ( .A1(a4stg_shl_cnt[3]), .A2(n1815), .A3(n1546), .A4(n1765), 
        .Y(a4stg_shl[21]) );
  AO22X1_RVT U2424 ( .A1(n1875), .A2(a4stg_shl[21]), .A3(n1766), .A4(n1877), 
        .Y(n1768) );
  AO22X1_RVT U2425 ( .A1(n1772), .A2(n1870), .A3(a4stg_rnd_frac[21]), .A4(
        n2526), .Y(n1767) );
  OR2X1_RVT U2426 ( .A1(n1768), .A2(n1767), .Y(a4stg_rnd_frac_pre2_in[21]) );
  OA221X1_RVT U2427 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[6]), .A3(n1800), .A4(a4stg_shl_data[5]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1781) );
  AO22X1_RVT U2428 ( .A1(a4stg_shl_cnt[1]), .A2(n1781), .A3(n1813), .A4(n1769), 
        .Y(n1795) );
  AO22X1_RVT U2429 ( .A1(a4stg_shl_cnt[2]), .A2(n1795), .A3(n1826), .A4(n1770), 
        .Y(n1822) );
  AO22X1_RVT U2430 ( .A1(a4stg_shl_cnt[3]), .A2(n1822), .A3(n1546), .A4(n1771), 
        .Y(a4stg_shl[20]) );
  AO22X1_RVT U2431 ( .A1(n1875), .A2(a4stg_shl[20]), .A3(n1772), .A4(n1877), 
        .Y(n1774) );
  AO22X1_RVT U2432 ( .A1(n1778), .A2(n1870), .A3(a4stg_rnd_frac[20]), .A4(
        n2526), .Y(n1773) );
  OR2X1_RVT U2433 ( .A1(n1774), .A2(n1773), .Y(a4stg_rnd_frac_pre2_in[20]) );
  OA221X1_RVT U2434 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[5]), .A3(n1800), .A4(a4stg_shl_data[4]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1787) );
  AO22X1_RVT U2435 ( .A1(a4stg_shl_cnt[1]), .A2(n1787), .A3(n1813), .A4(n1775), 
        .Y(n1802) );
  AO22X1_RVT U2436 ( .A1(a4stg_shl_cnt[2]), .A2(n1802), .A3(n1826), .A4(n1776), 
        .Y(n1827) );
  AO22X1_RVT U2437 ( .A1(a4stg_shl_cnt[3]), .A2(n1827), .A3(n1546), .A4(n1777), 
        .Y(a4stg_shl[19]) );
  AO22X1_RVT U2438 ( .A1(n1875), .A2(a4stg_shl[19]), .A3(n1778), .A4(n1877), 
        .Y(n1780) );
  AO22X1_RVT U2439 ( .A1(n1784), .A2(n1870), .A3(a4stg_rnd_frac[19]), .A4(
        n2526), .Y(n1779) );
  OR2X1_RVT U2440 ( .A1(n1780), .A2(n1779), .Y(a4stg_rnd_frac_pre2_in[19]) );
  OA221X1_RVT U2441 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[4]), .A3(n1800), .A4(a4stg_shl_data[3]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1793) );
  AO22X1_RVT U2442 ( .A1(a4stg_shl_cnt[1]), .A2(n1793), .A3(n1813), .A4(n1781), 
        .Y(n1807) );
  AO22X1_RVT U2443 ( .A1(a4stg_shl_cnt[2]), .A2(n1807), .A3(n1826), .A4(n1782), 
        .Y(n1831) );
  AO22X1_RVT U2444 ( .A1(a4stg_shl_cnt[3]), .A2(n1831), .A3(n1546), .A4(n1783), 
        .Y(a4stg_shl[18]) );
  AO22X1_RVT U2445 ( .A1(n1875), .A2(a4stg_shl[18]), .A3(n1784), .A4(n1877), 
        .Y(n1786) );
  AO22X1_RVT U2446 ( .A1(n1790), .A2(n1870), .A3(a4stg_rnd_frac[18]), .A4(
        n2526), .Y(n1785) );
  OR2X1_RVT U2447 ( .A1(n1786), .A2(n1785), .Y(a4stg_rnd_frac_pre2_in[18]) );
  OA221X1_RVT U2448 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[3]), .A3(n1800), .A4(a4stg_shl_data[2]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1801) );
  AO22X1_RVT U2449 ( .A1(a4stg_shl_cnt[1]), .A2(n1801), .A3(n1813), .A4(n1787), 
        .Y(n1814) );
  AO22X1_RVT U2450 ( .A1(a4stg_shl_cnt[2]), .A2(n1814), .A3(n1826), .A4(n1788), 
        .Y(n1836) );
  AO22X1_RVT U2451 ( .A1(a4stg_shl_cnt[3]), .A2(n1836), .A3(n1546), .A4(n1789), 
        .Y(a4stg_shl[17]) );
  AO22X1_RVT U2452 ( .A1(n1875), .A2(a4stg_shl[17]), .A3(n1790), .A4(n1877), 
        .Y(n1792) );
  AO22X1_RVT U2453 ( .A1(n1797), .A2(n1870), .A3(a4stg_rnd_frac[17]), .A4(
        n2526), .Y(n1791) );
  OR2X1_RVT U2454 ( .A1(n1792), .A2(n1791), .Y(a4stg_rnd_frac_pre2_in[17]) );
  AO22X1_RVT U2455 ( .A1(a4stg_shl_cnt[1]), .A2(n1794), .A3(n1813), .A4(n1793), 
        .Y(n1821) );
  AO22X1_RVT U2456 ( .A1(a4stg_shl_cnt[2]), .A2(n1821), .A3(n1826), .A4(n1795), 
        .Y(n1840) );
  AO22X1_RVT U2457 ( .A1(a4stg_shl_cnt[3]), .A2(n1840), .A3(n1546), .A4(n1796), 
        .Y(a4stg_shl[16]) );
  AO22X1_RVT U2458 ( .A1(n1875), .A2(a4stg_shl[16]), .A3(n1797), .A4(n1877), 
        .Y(n1799) );
  AO22X1_RVT U2459 ( .A1(n1804), .A2(n1870), .A3(a4stg_rnd_frac[16]), .A4(
        n2526), .Y(n1798) );
  OR2X1_RVT U2460 ( .A1(n1799), .A2(n1798), .Y(a4stg_rnd_frac_pre2_in[16]) );
  OA221X1_RVT U2461 ( .A1(a4stg_shl_cnt[0]), .A2(a4stg_shl_data[1]), .A3(n1800), .A4(a4stg_shl_data[0]), .A5(a4stg_shl_cnt_dec54_0[2]), .Y(n1812) );
  AO22X1_RVT U2462 ( .A1(a4stg_shl_cnt[1]), .A2(n1812), .A3(n1813), .A4(n1801), 
        .Y(n1861) );
  AO22X1_RVT U2463 ( .A1(a4stg_shl_cnt[2]), .A2(n1861), .A3(n1826), .A4(n1802), 
        .Y(n1845) );
  AO22X1_RVT U2464 ( .A1(a4stg_shl_cnt[3]), .A2(n1845), .A3(n1546), .A4(n1803), 
        .Y(a4stg_shl[15]) );
  AO22X1_RVT U2465 ( .A1(n1875), .A2(a4stg_shl[15]), .A3(n1804), .A4(n1877), 
        .Y(n1806) );
  AO22X1_RVT U2466 ( .A1(n1809), .A2(n1870), .A3(a4stg_rnd_frac[15]), .A4(
        n2526), .Y(n1805) );
  OR2X1_RVT U2467 ( .A1(n1806), .A2(n1805), .Y(a4stg_rnd_frac_pre2_in[15]) );
  AO22X1_RVT U2468 ( .A1(a4stg_shl_cnt[2]), .A2(n1832), .A3(n1826), .A4(n1807), 
        .Y(n1849) );
  AO22X1_RVT U2469 ( .A1(a4stg_shl_cnt[3]), .A2(n1849), .A3(n1546), .A4(n1808), 
        .Y(a4stg_shl[14]) );
  AO22X1_RVT U2470 ( .A1(n1875), .A2(a4stg_shl[14]), .A3(n1809), .A4(n1877), 
        .Y(n1811) );
  AO22X1_RVT U2471 ( .A1(n1816), .A2(n1870), .A3(a4stg_rnd_frac[14]), .A4(
        n2526), .Y(n1810) );
  OR2X1_RVT U2472 ( .A1(n1811), .A2(n1810), .Y(a4stg_rnd_frac_pre2_in[14]) );
  AND2X1_RVT U2473 ( .A1(n1813), .A2(n1812), .Y(n1868) );
  AO22X1_RVT U2474 ( .A1(a4stg_shl_cnt[2]), .A2(n1868), .A3(n1826), .A4(n1814), 
        .Y(n1853) );
  AO22X1_RVT U2475 ( .A1(a4stg_shl_cnt[3]), .A2(n1853), .A3(n1546), .A4(n1815), 
        .Y(a4stg_shl[13]) );
  AO22X1_RVT U2476 ( .A1(n1875), .A2(a4stg_shl[13]), .A3(n1816), .A4(n1877), 
        .Y(n1818) );
  AO22X1_RVT U2477 ( .A1(n1823), .A2(n1870), .A3(a4stg_rnd_frac[13]), .A4(
        n2526), .Y(n1817) );
  OR2X1_RVT U2478 ( .A1(n1818), .A2(n1817), .Y(a4stg_rnd_frac_pre2_in[13]) );
  AND2X1_RVT U2479 ( .A1(n1820), .A2(n1819), .Y(n1873) );
  AO22X1_RVT U2480 ( .A1(a4stg_shl_cnt[2]), .A2(n1873), .A3(n1826), .A4(n1821), 
        .Y(n1857) );
  AO22X1_RVT U2481 ( .A1(a4stg_shl_cnt[3]), .A2(n1857), .A3(n1546), .A4(n1822), 
        .Y(a4stg_shl[12]) );
  AO22X1_RVT U2482 ( .A1(n1875), .A2(a4stg_shl[12]), .A3(n1823), .A4(n1877), 
        .Y(n1825) );
  AO22X1_RVT U2483 ( .A1(n1828), .A2(n1870), .A3(a4stg_rnd_frac[12]), .A4(
        n2526), .Y(n1824) );
  OR2X1_RVT U2484 ( .A1(n1825), .A2(n1824), .Y(a4stg_rnd_frac_pre2_in[12]) );
  AND2X1_RVT U2485 ( .A1(a4stg_shl_cnt[3]), .A2(n1826), .Y(n1841) );
  AO22X1_RVT U2486 ( .A1(n1841), .A2(n1861), .A3(n1546), .A4(n1827), .Y(
        a4stg_shl[11]) );
  AO22X1_RVT U2487 ( .A1(n1875), .A2(a4stg_shl[11]), .A3(n1828), .A4(n1877), 
        .Y(n1830) );
  AO22X1_RVT U2488 ( .A1(n1833), .A2(n1870), .A3(a4stg_rnd_frac_11), .A4(n2526), .Y(n1829) );
  OR2X1_RVT U2489 ( .A1(n1830), .A2(n1829), .Y(a4stg_rnd_frac_pre2_in[11]) );
  AO22X1_RVT U2490 ( .A1(n1841), .A2(n1832), .A3(n1546), .A4(n1831), .Y(
        a4stg_shl[10]) );
  AO22X1_RVT U2491 ( .A1(n1875), .A2(a4stg_shl[10]), .A3(n1833), .A4(n1877), 
        .Y(n1835) );
  AO22X1_RVT U2492 ( .A1(n1837), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_10), .Y(n1834) );
  OR2X1_RVT U2493 ( .A1(n1835), .A2(n1834), .Y(a4stg_rnd_frac_pre2_in[10]) );
  AO22X1_RVT U2494 ( .A1(n1841), .A2(n1868), .A3(n1546), .A4(n1836), .Y(
        a4stg_shl[9]) );
  AO22X1_RVT U2495 ( .A1(n1875), .A2(a4stg_shl[9]), .A3(n1837), .A4(n1877), 
        .Y(n1839) );
  AO22X1_RVT U2496 ( .A1(n1842), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_9), 
        .Y(n1838) );
  OR2X1_RVT U2497 ( .A1(n1839), .A2(n1838), .Y(a4stg_rnd_frac_pre2_in[9]) );
  AO22X1_RVT U2498 ( .A1(n1841), .A2(n1873), .A3(n1546), .A4(n1840), .Y(
        a4stg_shl[8]) );
  AO22X1_RVT U2499 ( .A1(n1875), .A2(a4stg_shl[8]), .A3(n1842), .A4(n1877), 
        .Y(n1844) );
  AO22X1_RVT U2500 ( .A1(n1846), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_8), 
        .Y(n1843) );
  OR2X1_RVT U2501 ( .A1(n1844), .A2(n1843), .Y(a4stg_rnd_frac_pre2_in[8]) );
  AND2X1_RVT U2502 ( .A1(n1546), .A2(n1845), .Y(a4stg_shl[7]) );
  AO22X1_RVT U2503 ( .A1(a4stg_shl[7]), .A2(n1875), .A3(n1846), .A4(n1877), 
        .Y(n1848) );
  AO22X1_RVT U2504 ( .A1(n1850), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_7), 
        .Y(n1847) );
  OR2X1_RVT U2505 ( .A1(n1848), .A2(n1847), .Y(a4stg_rnd_frac_pre2_in[7]) );
  AND2X1_RVT U2506 ( .A1(n1546), .A2(n1849), .Y(a4stg_shl[6]) );
  AO22X1_RVT U2507 ( .A1(a4stg_shl[6]), .A2(n1875), .A3(n1850), .A4(n1877), 
        .Y(n1852) );
  AO22X1_RVT U2508 ( .A1(n1854), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_6), 
        .Y(n1851) );
  OR2X1_RVT U2509 ( .A1(n1852), .A2(n1851), .Y(a4stg_rnd_frac_pre2_in[6]) );
  AND2X1_RVT U2510 ( .A1(n1546), .A2(n1853), .Y(a4stg_shl[5]) );
  AO22X1_RVT U2511 ( .A1(a4stg_shl[5]), .A2(n1875), .A3(n1854), .A4(n1877), 
        .Y(n1856) );
  AO22X1_RVT U2512 ( .A1(n1858), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_5), 
        .Y(n1855) );
  OR2X1_RVT U2513 ( .A1(n1856), .A2(n1855), .Y(a4stg_rnd_frac_pre2_in[5]) );
  AND2X1_RVT U2514 ( .A1(n1546), .A2(n1857), .Y(a4stg_shl[4]) );
  AO22X1_RVT U2515 ( .A1(a4stg_shl[4]), .A2(n1875), .A3(n1858), .A4(n1877), 
        .Y(n1860) );
  AO22X1_RVT U2516 ( .A1(n1862), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_4), 
        .Y(n1859) );
  OR2X1_RVT U2517 ( .A1(n1860), .A2(n1859), .Y(a4stg_rnd_frac_pre2_in[4]) );
  AND2X1_RVT U2518 ( .A1(n1874), .A2(n1861), .Y(a4stg_shl[3]) );
  AO22X1_RVT U2519 ( .A1(a4stg_shl[3]), .A2(n1875), .A3(n1862), .A4(n1877), 
        .Y(n1864) );
  AO22X1_RVT U2520 ( .A1(n1865), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_3), 
        .Y(n1863) );
  OR2X1_RVT U2521 ( .A1(n1864), .A2(n1863), .Y(a4stg_rnd_frac_pre2_in[3]) );
  AO22X1_RVT U2522 ( .A1(n1870), .A2(n1869), .A3(n1865), .A4(n1877), .Y(n1867)
         );
  AO22X1_RVT U2523 ( .A1(a4stg_shl[2]), .A2(n1875), .A3(n2526), .A4(
        a4stg_rnd_frac_2), .Y(n1866) );
  OR2X1_RVT U2524 ( .A1(n1867), .A2(n1866), .Y(a4stg_rnd_frac_pre2_in[2]) );
  AND2X1_RVT U2525 ( .A1(n1874), .A2(n1868), .Y(a4stg_shl[1]) );
  AO22X1_RVT U2526 ( .A1(a4stg_shl[1]), .A2(n1875), .A3(n1869), .A4(n1877), 
        .Y(n1872) );
  AO22X1_RVT U2527 ( .A1(n1876), .A2(n1870), .A3(n2526), .A4(a4stg_rnd_frac_1), 
        .Y(n1871) );
  OR2X1_RVT U2528 ( .A1(n1872), .A2(n1871), .Y(a4stg_rnd_frac_pre2_in[1]) );
  AND2X1_RVT U2529 ( .A1(n1874), .A2(n1873), .Y(a4stg_shl[0]) );
  AO222X1_RVT U2530 ( .A1(n2526), .A2(a4stg_rnd_frac_pre2[0]), .A3(n1877), 
        .A4(n1876), .A5(n1875), .A6(a4stg_shl[0]), .Y(
        a4stg_rnd_frac_pre2_in[0]) );
  AND2X1_RVT U2531 ( .A1(a3stg_ld0_frac[63]), .A2(a3stg_denorm_inva), .Y(
        a4stg_shl_data_in[63]) );
  AO22X1_RVT U2532 ( .A1(n5), .A2(a3stg_ld0_frac[63]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[62]), .Y(a4stg_shl_data_in[62]) );
  AO22X1_RVT U2533 ( .A1(n5), .A2(a3stg_ld0_frac[62]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[61]), .Y(a4stg_shl_data_in[61]) );
  AO22X1_RVT U2534 ( .A1(n5), .A2(a3stg_ld0_frac[61]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[60]), .Y(a4stg_shl_data_in[60]) );
  AO22X1_RVT U2535 ( .A1(n5), .A2(a3stg_ld0_frac[60]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[59]), .Y(a4stg_shl_data_in[59]) );
  AO22X1_RVT U2536 ( .A1(n5), .A2(a3stg_ld0_frac[59]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[58]), .Y(a4stg_shl_data_in[58]) );
  AO22X1_RVT U2537 ( .A1(n5), .A2(a3stg_ld0_frac[58]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[57]), .Y(a4stg_shl_data_in[57]) );
  AO22X1_RVT U2538 ( .A1(n5), .A2(a3stg_ld0_frac[57]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[56]), .Y(a4stg_shl_data_in[56]) );
  AO22X1_RVT U2539 ( .A1(n5), .A2(a3stg_ld0_frac[56]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[55]), .Y(a4stg_shl_data_in[55]) );
  AO22X1_RVT U2540 ( .A1(n5), .A2(a3stg_ld0_frac[55]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[54]), .Y(a4stg_shl_data_in[54]) );
  AO22X1_RVT U2541 ( .A1(n5), .A2(a3stg_ld0_frac[54]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[53]), .Y(a4stg_shl_data_in[53]) );
  AO22X1_RVT U2542 ( .A1(n5), .A2(a3stg_ld0_frac[53]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[52]), .Y(a4stg_shl_data_in[52]) );
  AO22X1_RVT U2543 ( .A1(n5), .A2(a3stg_ld0_frac[52]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[51]), .Y(a4stg_shl_data_in[51]) );
  AO22X1_RVT U2544 ( .A1(n5), .A2(a3stg_ld0_frac[51]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[50]), .Y(a4stg_shl_data_in[50]) );
  AO22X1_RVT U2545 ( .A1(n5), .A2(a3stg_ld0_frac[50]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[49]), .Y(a4stg_shl_data_in[49]) );
  AO22X1_RVT U2546 ( .A1(n5), .A2(a3stg_ld0_frac[49]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[48]), .Y(a4stg_shl_data_in[48]) );
  AO22X1_RVT U2547 ( .A1(n5), .A2(a3stg_ld0_frac[48]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[47]), .Y(a4stg_shl_data_in[47]) );
  AO22X1_RVT U2548 ( .A1(n5), .A2(a3stg_ld0_frac[47]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[46]), .Y(a4stg_shl_data_in[46]) );
  AO22X1_RVT U2549 ( .A1(n5), .A2(a3stg_ld0_frac[46]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[45]), .Y(a4stg_shl_data_in[45]) );
  AO22X1_RVT U2550 ( .A1(n5), .A2(a3stg_ld0_frac[45]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[44]), .Y(a4stg_shl_data_in[44]) );
  AO22X1_RVT U2551 ( .A1(n5), .A2(a3stg_ld0_frac[44]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[43]), .Y(a4stg_shl_data_in[43]) );
  AO22X1_RVT U2552 ( .A1(n5), .A2(a3stg_ld0_frac[43]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[42]), .Y(a4stg_shl_data_in[42]) );
  AO22X1_RVT U2553 ( .A1(n5), .A2(a3stg_ld0_frac[42]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[41]), .Y(a4stg_shl_data_in[41]) );
  AO22X1_RVT U2554 ( .A1(n5), .A2(a3stg_ld0_frac[41]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[40]), .Y(a4stg_shl_data_in[40]) );
  AO22X1_RVT U2555 ( .A1(n5), .A2(a3stg_ld0_frac[40]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[39]), .Y(a4stg_shl_data_in[39]) );
  AO22X1_RVT U2556 ( .A1(n5), .A2(a3stg_ld0_frac[39]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[38]), .Y(a4stg_shl_data_in[38]) );
  AO22X1_RVT U2557 ( .A1(n5), .A2(a3stg_ld0_frac[38]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[37]), .Y(a4stg_shl_data_in[37]) );
  AO22X1_RVT U2558 ( .A1(n5), .A2(a3stg_ld0_frac[37]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[36]), .Y(a4stg_shl_data_in[36]) );
  AO22X1_RVT U2559 ( .A1(n5), .A2(a3stg_ld0_frac[36]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[35]), .Y(a4stg_shl_data_in[35]) );
  AO22X1_RVT U2560 ( .A1(n5), .A2(a3stg_ld0_frac[35]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[34]), .Y(a4stg_shl_data_in[34]) );
  AO22X1_RVT U2561 ( .A1(n5), .A2(a3stg_ld0_frac[34]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[33]), .Y(a4stg_shl_data_in[33]) );
  AO22X1_RVT U2562 ( .A1(n5), .A2(a3stg_ld0_frac[33]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[32]), .Y(a4stg_shl_data_in[32]) );
  AO22X1_RVT U2563 ( .A1(n5), .A2(a3stg_ld0_frac[32]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[31]), .Y(a4stg_shl_data_in[31]) );
  AO22X1_RVT U2564 ( .A1(n5), .A2(a3stg_ld0_frac[31]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[30]), .Y(a4stg_shl_data_in[30]) );
  AO22X1_RVT U2565 ( .A1(n5), .A2(a3stg_ld0_frac[30]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[29]), .Y(a4stg_shl_data_in[29]) );
  AO22X1_RVT U2566 ( .A1(n5), .A2(a3stg_ld0_frac[29]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[28]), .Y(a4stg_shl_data_in[28]) );
  AO22X1_RVT U2567 ( .A1(n5), .A2(a3stg_ld0_frac[28]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[27]), .Y(a4stg_shl_data_in[27]) );
  AO22X1_RVT U2568 ( .A1(n5), .A2(a3stg_ld0_frac[27]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[26]), .Y(a4stg_shl_data_in[26]) );
  AO22X1_RVT U2569 ( .A1(n5), .A2(a3stg_ld0_frac[26]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[25]), .Y(a4stg_shl_data_in[25]) );
  AO22X1_RVT U2570 ( .A1(n5), .A2(a3stg_ld0_frac[25]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[24]), .Y(a4stg_shl_data_in[24]) );
  AO22X1_RVT U2571 ( .A1(n5), .A2(a3stg_ld0_frac[24]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[23]), .Y(a4stg_shl_data_in[23]) );
  AO22X1_RVT U2572 ( .A1(n5), .A2(a3stg_ld0_frac[23]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[22]), .Y(a4stg_shl_data_in[22]) );
  AO22X1_RVT U2573 ( .A1(n5), .A2(a3stg_ld0_frac[22]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[21]), .Y(a4stg_shl_data_in[21]) );
  AO22X1_RVT U2574 ( .A1(n5), .A2(a3stg_ld0_frac[21]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[20]), .Y(a4stg_shl_data_in[20]) );
  AO22X1_RVT U2575 ( .A1(n5), .A2(a3stg_ld0_frac[20]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[19]), .Y(a4stg_shl_data_in[19]) );
  AO22X1_RVT U2576 ( .A1(n5), .A2(a3stg_ld0_frac[19]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[18]), .Y(a4stg_shl_data_in[18]) );
  AO22X1_RVT U2577 ( .A1(n5), .A2(a3stg_ld0_frac[18]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[17]), .Y(a4stg_shl_data_in[17]) );
  AO22X1_RVT U2578 ( .A1(n5), .A2(a3stg_ld0_frac[17]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[16]), .Y(a4stg_shl_data_in[16]) );
  AO22X1_RVT U2579 ( .A1(n5), .A2(a3stg_ld0_frac[16]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[15]), .Y(a4stg_shl_data_in[15]) );
  AO22X1_RVT U2580 ( .A1(n5), .A2(a3stg_ld0_frac[15]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[14]), .Y(a4stg_shl_data_in[14]) );
  AO22X1_RVT U2581 ( .A1(n5), .A2(a3stg_ld0_frac[14]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[13]), .Y(a4stg_shl_data_in[13]) );
  AO22X1_RVT U2582 ( .A1(n5), .A2(a3stg_ld0_frac[13]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[12]), .Y(a4stg_shl_data_in[12]) );
  AO22X1_RVT U2583 ( .A1(n5), .A2(a3stg_ld0_frac[12]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[11]), .Y(a4stg_shl_data_in[11]) );
  AO22X1_RVT U2584 ( .A1(n5), .A2(a3stg_ld0_frac[11]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[10]), .Y(a4stg_shl_data_in[10]) );
  AO22X1_RVT U2585 ( .A1(n5), .A2(a3stg_ld0_frac[10]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[9]), .Y(a4stg_shl_data_in[9]) );
  AO22X1_RVT U2586 ( .A1(n5), .A2(a3stg_ld0_frac[9]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[8]), .Y(a4stg_shl_data_in[8]) );
  AO22X1_RVT U2587 ( .A1(n5), .A2(a3stg_ld0_frac[8]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[7]), .Y(a4stg_shl_data_in[7]) );
  AO22X1_RVT U2588 ( .A1(n5), .A2(a3stg_ld0_frac[7]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[6]), .Y(a4stg_shl_data_in[6]) );
  AO22X1_RVT U2589 ( .A1(n5), .A2(a3stg_ld0_frac[6]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[5]), .Y(a4stg_shl_data_in[5]) );
  AO22X1_RVT U2590 ( .A1(n5), .A2(a3stg_ld0_frac[5]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[4]), .Y(a4stg_shl_data_in[4]) );
  AO22X1_RVT U2591 ( .A1(n5), .A2(a3stg_ld0_frac[4]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[3]), .Y(a4stg_shl_data_in[3]) );
  AO22X1_RVT U2592 ( .A1(n5), .A2(a3stg_ld0_frac[3]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[2]), .Y(a4stg_shl_data_in[2]) );
  AO22X1_RVT U2593 ( .A1(n5), .A2(a3stg_ld0_frac[2]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[1]), .Y(a4stg_shl_data_in[1]) );
  AO22X1_RVT U2594 ( .A1(n5), .A2(a3stg_ld0_frac[1]), .A3(a3stg_denorm_inva), 
        .A4(a3stg_ld0_frac[0]), .Y(a4stg_shl_data_in[0]) );
  NOR4X1_RVT U2595 ( .A1(a4stg_rnd_frac_47), .A2(a4stg_rnd_frac_45), .A3(
        a4stg_rnd_frac_44), .A4(a4stg_rnd_frac_42), .Y(n1884) );
  NOR4X1_RVT U2596 ( .A1(a4stg_rnd_frac_43), .A2(a4stg_rnd_frac_41), .A3(
        a4stg_rnd_frac_63), .A4(a4stg_rnd_frac_40), .Y(n1883) );
  NOR4X1_RVT U2597 ( .A1(a4stg_rnd_frac_54), .A2(a4stg_rnd_frac_53), .A3(
        a4stg_rnd_frac_52), .A4(a4stg_rnd_frac_51), .Y(n1881) );
  NOR4X1_RVT U2598 ( .A1(a4stg_rnd_frac_50), .A2(a4stg_rnd_frac_49), .A3(
        a4stg_rnd_frac_48), .A4(a4stg_rnd_frac_46), .Y(n1880) );
  NOR4X1_RVT U2599 ( .A1(a4stg_rnd_frac_62), .A2(a4stg_rnd_frac_61), .A3(
        a4stg_rnd_frac_60), .A4(a4stg_rnd_frac_57), .Y(n1879) );
  NOR4X1_RVT U2600 ( .A1(a4stg_rnd_frac_59), .A2(a4stg_rnd_frac_58), .A3(
        a4stg_rnd_frac_56), .A4(a4stg_rnd_frac_55), .Y(n1878) );
  AND4X1_RVT U2601 ( .A1(n1881), .A2(n1880), .A3(n1879), .A4(n1878), .Y(n1882)
         );
  NAND4X0_RVT U2602 ( .A1(n1885), .A2(n1884), .A3(n1883), .A4(n1882), .Y(
        a4stg_frac_neq_0) );
  NOR4X1_RVT U2603 ( .A1(a4stg_shl_data[31]), .A2(a4stg_shl_data[15]), .A3(
        a4stg_shl_data[47]), .A4(a4stg_shl_data[63]), .Y(n1889) );
  NOR4X1_RVT U2604 ( .A1(a4stg_shl_data[14]), .A2(a4stg_shl_data[30]), .A3(
        a4stg_shl_data[62]), .A4(a4stg_shl_data[46]), .Y(n1888) );
  NOR4X1_RVT U2605 ( .A1(a4stg_shl_data[61]), .A2(a4stg_shl_data[13]), .A3(
        a4stg_shl_data[45]), .A4(a4stg_shl_data[29]), .Y(n1887) );
  NOR4X1_RVT U2606 ( .A1(a4stg_shl_data[60]), .A2(a4stg_shl_data[28]), .A3(
        a4stg_shl_data[44]), .A4(a4stg_shl_data[12]), .Y(n1886) );
  NAND4X0_RVT U2607 ( .A1(n1889), .A2(n1888), .A3(n1887), .A4(n1886), .Y(n1905) );
  NOR4X1_RVT U2608 ( .A1(a4stg_shl_data[27]), .A2(a4stg_shl_data[59]), .A3(
        a4stg_shl_data[43]), .A4(a4stg_shl_data[11]), .Y(n1893) );
  NOR4X1_RVT U2609 ( .A1(a4stg_shl_data[10]), .A2(a4stg_shl_data[42]), .A3(
        a4stg_shl_data[26]), .A4(a4stg_shl_data[58]), .Y(n1892) );
  NOR4X1_RVT U2610 ( .A1(a4stg_shl_data[57]), .A2(a4stg_shl_data[9]), .A3(
        a4stg_shl_data[25]), .A4(a4stg_shl_data[41]), .Y(n1891) );
  NOR4X1_RVT U2611 ( .A1(a4stg_shl_data[24]), .A2(a4stg_shl_data[56]), .A3(
        a4stg_shl_data[8]), .A4(a4stg_shl_data[40]), .Y(n1890) );
  NAND4X0_RVT U2612 ( .A1(n1893), .A2(n1892), .A3(n1891), .A4(n1890), .Y(n1904) );
  NOR4X1_RVT U2613 ( .A1(a4stg_shl_data[55]), .A2(a4stg_shl_data[39]), .A3(
        a4stg_shl_data[7]), .A4(a4stg_shl_data[23]), .Y(n1897) );
  NOR4X1_RVT U2614 ( .A1(a4stg_shl_data[54]), .A2(a4stg_shl_data[6]), .A3(
        a4stg_shl_data[38]), .A4(a4stg_shl_data[22]), .Y(n1896) );
  NOR4X1_RVT U2615 ( .A1(a4stg_shl_data[53]), .A2(a4stg_shl_data[5]), .A3(
        a4stg_shl_data[21]), .A4(a4stg_shl_data[37]), .Y(n1895) );
  NOR4X1_RVT U2616 ( .A1(a4stg_shl_data[36]), .A2(a4stg_shl_data[20]), .A3(
        a4stg_shl_data[52]), .A4(a4stg_shl_data[4]), .Y(n1894) );
  NAND4X0_RVT U2617 ( .A1(n1897), .A2(n1896), .A3(n1895), .A4(n1894), .Y(n1903) );
  NOR4X1_RVT U2618 ( .A1(a4stg_shl_data[51]), .A2(a4stg_shl_data[19]), .A3(
        a4stg_shl_data[3]), .A4(a4stg_shl_data[35]), .Y(n1901) );
  NOR4X1_RVT U2619 ( .A1(a4stg_shl_data[18]), .A2(a4stg_shl_data[50]), .A3(
        a4stg_shl_data[2]), .A4(a4stg_shl_data[34]), .Y(n1900) );
  NOR4X1_RVT U2620 ( .A1(a4stg_shl_data[1]), .A2(a4stg_shl_data[17]), .A3(
        a4stg_shl_data[49]), .A4(a4stg_shl_data[33]), .Y(n1899) );
  NOR4X1_RVT U2621 ( .A1(a4stg_shl_data[16]), .A2(a4stg_shl_data[0]), .A3(
        a4stg_shl_data[32]), .A4(a4stg_shl_data[48]), .Y(n1898) );
  NAND4X0_RVT U2622 ( .A1(n1901), .A2(n1900), .A3(n1899), .A4(n1898), .Y(n1902) );
  OR4X1_RVT U2623 ( .A1(n1905), .A2(n1904), .A3(n1903), .A4(n1902), .Y(
        a4stg_shl_data_neq_0) );
  AO22X1_RVT U2624 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[63]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[63]), .Y(n1906) );
  OR2X1_RVT U2625 ( .A1(n1918), .A2(n1906), .Y(add_frac_out[63]) );
  AO22X1_RVT U2626 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[10]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[10]), .Y(n1907) );
  OR2X1_RVT U2627 ( .A1(n1918), .A2(n1907), .Y(add_frac_out[10]) );
  AO22X1_RVT U2628 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[9]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[9]), .Y(n1908) );
  OR2X1_RVT U2629 ( .A1(n1918), .A2(n1908), .Y(add_frac_out[9]) );
  AO22X1_RVT U2630 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[8]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[8]), .Y(n1909) );
  OR2X1_RVT U2631 ( .A1(n1918), .A2(n1909), .Y(add_frac_out[8]) );
  AO22X1_RVT U2632 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[7]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[7]), .Y(n1910) );
  OR2X1_RVT U2633 ( .A1(n1918), .A2(n1910), .Y(add_frac_out[7]) );
  AO22X1_RVT U2634 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[6]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[6]), .Y(n1911) );
  OR2X1_RVT U2635 ( .A1(n1918), .A2(n1911), .Y(add_frac_out[6]) );
  AO22X1_RVT U2636 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[5]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[5]), .Y(n1912) );
  OR2X1_RVT U2637 ( .A1(n1918), .A2(n1912), .Y(add_frac_out[5]) );
  AO22X1_RVT U2638 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[4]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[4]), .Y(n1913) );
  OR2X1_RVT U2639 ( .A1(n1918), .A2(n1913), .Y(add_frac_out[4]) );
  AO22X1_RVT U2640 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[3]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[3]), .Y(n1914) );
  OR2X1_RVT U2641 ( .A1(n1918), .A2(n1914), .Y(add_frac_out[3]) );
  AO22X1_RVT U2642 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[2]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[2]), .Y(n1915) );
  OR2X1_RVT U2643 ( .A1(n1918), .A2(n1915), .Y(add_frac_out[2]) );
  AO22X1_RVT U2644 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[1]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[1]), .Y(n1916) );
  OR2X1_RVT U2645 ( .A1(n1918), .A2(n1916), .Y(add_frac_out[1]) );
  AO22X1_RVT U2646 ( .A1(a5stg_frac_out_shl), .A2(a5stg_shl[0]), .A3(
        a5stg_frac_out_rnd_frac), .A4(a5stg_rnd_frac[0]), .Y(n1917) );
  OR2X1_RVT U2647 ( .A1(n1918), .A2(n1917), .Y(add_frac_out[0]) );
  NAND4X0_RVT U2648 ( .A1(n1919), .A2(n1922), .A3(a3stg_inc_exp_inv), .A4(
        n1921), .Y(a3stg_dec_exp_inv) );
  AO21X1_RVT U2649 ( .A1(n1922), .A2(n1921), .A3(n1920), .Y(a3stg_same_exp_inv) );
  NAND2X0_RVT U2650 ( .A1(n2045), .A2(n2449), .Y(n2035) );
  INVX1_RVT U2651 ( .A(n2035), .Y(n1982) );
  NAND2X0_RVT U2652 ( .A1(n2450), .A2(n1982), .Y(n1948) );
  INVX1_RVT U2653 ( .A(n1948), .Y(n1925) );
  NAND3X0_RVT U2654 ( .A1(a2stg_frac2a[63]), .A2(a2stg_shr_cnt_0[0]), .A3(
        n1925), .Y(n1927) );
  OA21X1_RVT U2655 ( .A1(a2stg_shr_frac2_shr_dbl), .A2(a2stg_shr_frac2_shr_sng), .A3(a2stg_expadd_11), .Y(n2176) );
  AO22X1_RVT U2656 ( .A1(n1923), .A2(n2176), .A3(\DP_OP_16J2_123_4718/n1 ), 
        .A4(n2526), .Y(n1924) );
  HADDX1_RVT U2657 ( .A0(a2stg_sub_step), .B0(n1924), .SO(n1731) );
  INVX1_RVT U2658 ( .A(a2stg_frac2a[62]), .Y(n1947) );
  NAND2X0_RVT U2659 ( .A1(a2stg_shr_cnt_0[0]), .A2(n1925), .Y(n1926) );
  INVX1_RVT U2660 ( .A(a2stg_frac2a[63]), .Y(n1954) );
  NAND2X0_RVT U2661 ( .A1(a2stg_shr_cnt_0[1]), .A2(n1925), .Y(n1932) );
  OA22X1_RVT U2662 ( .A1(n1947), .A2(n1926), .A3(n1954), .A4(n1932), .Y(n1933)
         );
  INVX1_RVT U2663 ( .A(n2176), .Y(n1960) );
  OA22X1_RVT U2664 ( .A1(n1933), .A2(n1960), .A3(n1986), .A4(n1927), .Y(n1930)
         );
  INVX1_RVT U2665 ( .A(a2stg_expadd_11), .Y(n1928) );
  NAND2X0_RVT U2666 ( .A1(a2stg_shr_frac2_max), .A2(n1928), .Y(n2528) );
  NAND2X0_RVT U2667 ( .A1(a3stg_frac2[62]), .A2(n2526), .Y(n1929) );
  NAND3X0_RVT U2668 ( .A1(n1930), .A2(n2528), .A3(n1929), .Y(n1931) );
  HADDX1_RVT U2669 ( .A0(a2stg_sub_step), .B0(n1931), .SO(n1730) );
  NAND2X0_RVT U2670 ( .A1(n2345), .A2(n1982), .Y(n1981) );
  INVX1_RVT U2671 ( .A(a2stg_frac2a[61]), .Y(n1991) );
  OA22X1_RVT U2672 ( .A1(n1954), .A2(n1981), .A3(n1991), .A4(n1948), .Y(n1937)
         );
  OA22X1_RVT U2673 ( .A1(n1937), .A2(n1957), .A3(n1947), .A4(n1932), .Y(n1938)
         );
  OA22X1_RVT U2674 ( .A1(n1938), .A2(n1960), .A3(n1933), .A4(n1986), .Y(n1935)
         );
  NAND2X0_RVT U2675 ( .A1(a3stg_frac2[61]), .A2(n2526), .Y(n1934) );
  NAND3X0_RVT U2676 ( .A1(n1935), .A2(n2528), .A3(n1934), .Y(n1936) );
  HADDX1_RVT U2677 ( .A0(a2stg_sub_step), .B0(n1936), .SO(n1729) );
  NAND2X0_RVT U2678 ( .A1(a3stg_frac2[60]), .A2(n2526), .Y(n1940) );
  INVX1_RVT U2679 ( .A(a2stg_frac2a[60]), .Y(n2000) );
  OA22X1_RVT U2680 ( .A1(n2000), .A2(n1948), .A3(n1947), .A4(n1981), .Y(n1942)
         );
  OA22X1_RVT U2681 ( .A1(n1942), .A2(n1957), .A3(n1937), .A4(n1958), .Y(n1943)
         );
  OA22X1_RVT U2682 ( .A1(n1938), .A2(n1986), .A3(n1943), .A4(n1960), .Y(n1939)
         );
  NAND3X0_RVT U2683 ( .A1(n1940), .A2(n2528), .A3(n1939), .Y(n1941) );
  HADDX1_RVT U2684 ( .A0(a2stg_sub_step), .B0(n1941), .SO(n1728) );
  NAND2X0_RVT U2685 ( .A1(a3stg_frac2[59]), .A2(n2526), .Y(n1945) );
  NAND2X0_RVT U2686 ( .A1(n2326), .A2(n1982), .Y(n1999) );
  INVX1_RVT U2687 ( .A(a2stg_frac2a[59]), .Y(n2008) );
  OA222X1_RVT U2688 ( .A1(n1954), .A2(n1999), .A3(n2008), .A4(n1948), .A5(
        n1991), .A6(n1981), .Y(n1949) );
  OA22X1_RVT U2689 ( .A1(n1949), .A2(n1957), .A3(n1942), .A4(n1958), .Y(n1950)
         );
  OA22X1_RVT U2690 ( .A1(n1950), .A2(n1960), .A3(n1943), .A4(n1986), .Y(n1944)
         );
  NAND3X0_RVT U2691 ( .A1(n1945), .A2(n2528), .A3(n1944), .Y(n1946) );
  HADDX1_RVT U2692 ( .A0(a2stg_sub_step), .B0(n1946), .SO(n1727) );
  NAND2X0_RVT U2693 ( .A1(a3stg_frac2[58]), .A2(n2526), .Y(n1952) );
  INVX1_RVT U2694 ( .A(a2stg_frac2a[58]), .Y(n2016) );
  OA222X1_RVT U2695 ( .A1(n2016), .A2(n1948), .A3(n2000), .A4(n1981), .A5(
        n1947), .A6(n1999), .Y(n1959) );
  OA22X1_RVT U2696 ( .A1(n1949), .A2(n1958), .A3(n1959), .A4(n1957), .Y(n1961)
         );
  OA22X1_RVT U2697 ( .A1(n1961), .A2(n1960), .A3(n1950), .A4(n1986), .Y(n1951)
         );
  NAND3X0_RVT U2698 ( .A1(n1952), .A2(n2528), .A3(n1951), .Y(n1953) );
  HADDX1_RVT U2699 ( .A0(a2stg_sub_step), .B0(n1953), .SO(n1726) );
  NAND2X0_RVT U2700 ( .A1(a3stg_frac2[57]), .A2(n2526), .Y(n1963) );
  INVX1_RVT U2701 ( .A(a2stg_frac2a[57]), .Y(n2025) );
  OA22X1_RVT U2702 ( .A1(n2467), .A2(n1991), .A3(n2448), .A4(n2025), .Y(n1956)
         );
  OA22X1_RVT U2703 ( .A1(n2465), .A2(n2008), .A3(n2456), .A4(n1954), .Y(n1955)
         );
  AO21X1_RVT U2704 ( .A1(n1956), .A2(n1955), .A3(n2035), .Y(n1965) );
  OA22X1_RVT U2705 ( .A1(n1959), .A2(n1958), .A3(n1957), .A4(n1965), .Y(n1970)
         );
  OA22X1_RVT U2706 ( .A1(n1961), .A2(n1986), .A3(n1970), .A4(n1960), .Y(n1962)
         );
  NAND3X0_RVT U2707 ( .A1(n1963), .A2(n2528), .A3(n1962), .Y(n1964) );
  HADDX1_RVT U2708 ( .A0(a2stg_sub_step), .B0(n1964), .SO(n1725) );
  AO22X1_RVT U2709 ( .A1(a2stg_frac2a[58]), .A2(n2345), .A3(a2stg_frac2a[62]), 
        .A4(n2476), .Y(n1967) );
  AO22X1_RVT U2710 ( .A1(a2stg_frac2a[60]), .A2(n2326), .A3(a2stg_frac2a[56]), 
        .A4(n2450), .Y(n1966) );
  OA21X1_RVT U2711 ( .A1(n1967), .A2(n1966), .A3(n1982), .Y(n1977) );
  AO22X1_RVT U2712 ( .A1(a2stg_shr_cnt_0[1]), .A2(n1968), .A3(
        a2stg_shr_cnt_0[0]), .A4(n1977), .Y(n1978) );
  AOI22X1_RVT U2713 ( .A1(n2176), .A2(n1978), .A3(a3stg_frac2[56]), .A4(n2526), 
        .Y(n1969) );
  AND2X1_RVT U2714 ( .A1(n2528), .A2(n1969), .Y(n1973) );
  INVX1_RVT U2715 ( .A(n1970), .Y(n1971) );
  NAND2X0_RVT U2716 ( .A1(n1971), .A2(a2stg_shr_frac2_shr_int), .Y(n1972) );
  AND2X1_RVT U2717 ( .A1(n1973), .A2(n1972), .Y(n1974) );
  HADDX1_RVT U2718 ( .A0(n1974), .B0(n2483), .SO(n1724) );
  NAND2X0_RVT U2719 ( .A1(n2476), .A2(n1982), .Y(n2017) );
  OA22X1_RVT U2720 ( .A1(n2008), .A2(n1999), .A3(n1991), .A4(n2017), .Y(n1976)
         );
  NAND2X0_RVT U2721 ( .A1(n2045), .A2(a2stg_shr_cnt_3[0]), .Y(n2112) );
  INVX1_RVT U2722 ( .A(n2112), .Y(n2054) );
  AOI22X1_RVT U2723 ( .A1(a2stg_frac2a[55]), .A2(n1982), .A3(a2stg_frac2a[63]), 
        .A4(n2054), .Y(n2026) );
  OA22X1_RVT U2724 ( .A1(n2026), .A2(n2448), .A3(n2025), .A4(n1981), .Y(n1975)
         );
  NAND2X0_RVT U2725 ( .A1(n1976), .A2(n1975), .Y(n1985) );
  AO22X1_RVT U2726 ( .A1(a2stg_shr_cnt_0[1]), .A2(n1977), .A3(
        a2stg_shr_cnt_0[0]), .A4(n1985), .Y(n1987) );
  NAND2X0_RVT U2727 ( .A1(a2stg_shr_frac2_shr_int), .A2(n1978), .Y(n1979) );
  NAND3X0_RVT U2728 ( .A1(n7), .A2(n2528), .A3(n1979), .Y(n1980) );
  HADDX1_RVT U2729 ( .A0(a2stg_sub_step), .B0(n1980), .SO(n1723) );
  INVX1_RVT U2730 ( .A(a2stg_frac2a[56]), .Y(n2036) );
  OA22X1_RVT U2731 ( .A1(n2000), .A2(n2017), .A3(n2036), .A4(n1981), .Y(n1984)
         );
  AOI22X1_RVT U2732 ( .A1(a2stg_frac2a[54]), .A2(n1982), .A3(a2stg_frac2a[62]), 
        .A4(n2054), .Y(n2034) );
  OA22X1_RVT U2733 ( .A1(n2034), .A2(n2448), .A3(n2016), .A4(n1999), .Y(n1983)
         );
  NAND2X0_RVT U2734 ( .A1(n1984), .A2(n1983), .Y(n1994) );
  AO22X1_RVT U2735 ( .A1(a2stg_shr_cnt_0[1]), .A2(n1985), .A3(
        a2stg_shr_cnt_0[0]), .A4(n1994), .Y(n1995) );
  AOI22X1_RVT U2736 ( .A1(n2176), .A2(n1995), .A3(a3stg_frac2[54]), .A4(n2526), 
        .Y(n1989) );
  NAND2X0_RVT U2737 ( .A1(a2stg_shr_frac2_shr_int), .A2(n1987), .Y(n1988) );
  NAND3X0_RVT U2738 ( .A1(n1989), .A2(n2528), .A3(n1988), .Y(n1990) );
  HADDX1_RVT U2739 ( .A0(a2stg_sub_step), .B0(n1990), .SO(n1722) );
  OA22X1_RVT U2740 ( .A1(n2025), .A2(n1999), .A3(n2008), .A4(n2017), .Y(n1993)
         );
  INVX1_RVT U2741 ( .A(a2stg_frac2a[53]), .Y(n2064) );
  OA22X1_RVT U2742 ( .A1(n2064), .A2(n2035), .A3(n1991), .A4(n2112), .Y(n2043)
         );
  OA22X1_RVT U2743 ( .A1(n2043), .A2(n2448), .A3(n2026), .A4(n2465), .Y(n1992)
         );
  NAND2X0_RVT U2744 ( .A1(n1993), .A2(n1992), .Y(n2003) );
  AO22X1_RVT U2745 ( .A1(a2stg_shr_cnt_0[1]), .A2(n1994), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2003), .Y(n2004) );
  AOI22X1_RVT U2746 ( .A1(n2176), .A2(n2004), .A3(a3stg_frac2[53]), .A4(n2526), 
        .Y(n1997) );
  NAND2X0_RVT U2747 ( .A1(a2stg_shr_frac2_shr_int), .A2(n1995), .Y(n1996) );
  NAND3X0_RVT U2748 ( .A1(n1997), .A2(n2528), .A3(n1996), .Y(n1998) );
  HADDX1_RVT U2749 ( .A0(a2stg_sub_step), .B0(n1998), .SO(n1721) );
  OA22X1_RVT U2750 ( .A1(n2016), .A2(n2017), .A3(n2036), .A4(n1999), .Y(n2002)
         );
  INVX1_RVT U2751 ( .A(a2stg_frac2a[52]), .Y(n2074) );
  OA22X1_RVT U2752 ( .A1(n2074), .A2(n2035), .A3(n2000), .A4(n2112), .Y(n2055)
         );
  OA22X1_RVT U2753 ( .A1(n2055), .A2(n2448), .A3(n2034), .A4(n2465), .Y(n2001)
         );
  NAND2X0_RVT U2754 ( .A1(n2002), .A2(n2001), .Y(n2011) );
  AO22X1_RVT U2755 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2003), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2011), .Y(n2012) );
  AOI22X1_RVT U2756 ( .A1(n2176), .A2(n2012), .A3(a3stg_frac2[52]), .A4(n2526), 
        .Y(n2006) );
  NAND2X0_RVT U2757 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2004), .Y(n2005) );
  NAND3X0_RVT U2758 ( .A1(n2006), .A2(n2528), .A3(n2005), .Y(n2007) );
  HADDX1_RVT U2759 ( .A0(a2stg_sub_step), .B0(n2007), .SO(n1720) );
  INVX1_RVT U2760 ( .A(a2stg_frac2a[51]), .Y(n2083) );
  OA22X1_RVT U2761 ( .A1(n2083), .A2(n2035), .A3(n2008), .A4(n2112), .Y(n2063)
         );
  OA22X1_RVT U2762 ( .A1(n2063), .A2(n2448), .A3(n2043), .A4(n2465), .Y(n2010)
         );
  OA22X1_RVT U2763 ( .A1(n2026), .A2(n2467), .A3(n2025), .A4(n2017), .Y(n2009)
         );
  NAND2X0_RVT U2764 ( .A1(n2010), .A2(n2009), .Y(n2020) );
  AO22X1_RVT U2765 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2011), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2020), .Y(n2021) );
  AOI22X1_RVT U2766 ( .A1(n2176), .A2(n2021), .A3(a3stg_frac2[51]), .A4(n2526), 
        .Y(n2014) );
  NAND2X0_RVT U2767 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2012), .Y(n2013) );
  NAND3X0_RVT U2768 ( .A1(n2014), .A2(n2528), .A3(n2013), .Y(n2015) );
  HADDX1_RVT U2769 ( .A0(a2stg_sub_step), .B0(n2015), .SO(n1719) );
  OA22X1_RVT U2770 ( .A1(n2055), .A2(n2465), .A3(n2034), .A4(n2467), .Y(n2019)
         );
  INVX1_RVT U2771 ( .A(a2stg_frac2a[50]), .Y(n2092) );
  OA22X1_RVT U2772 ( .A1(n2016), .A2(n2112), .A3(n2092), .A4(n2035), .Y(n2073)
         );
  OA22X1_RVT U2773 ( .A1(n2073), .A2(n2448), .A3(n2036), .A4(n2017), .Y(n2018)
         );
  NAND2X0_RVT U2774 ( .A1(n2019), .A2(n2018), .Y(n2029) );
  AO22X1_RVT U2775 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2020), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2029), .Y(n2030) );
  AOI22X1_RVT U2776 ( .A1(n2176), .A2(n2030), .A3(a3stg_frac2[50]), .A4(n2526), 
        .Y(n2023) );
  NAND2X0_RVT U2777 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2021), .Y(n2022) );
  NAND3X0_RVT U2778 ( .A1(n2023), .A2(n2528), .A3(n2022), .Y(n2024) );
  HADDX1_RVT U2779 ( .A0(a2stg_sub_step), .B0(n2024), .SO(n1718) );
  OA22X1_RVT U2780 ( .A1(n2025), .A2(n2112), .A3(n2103), .A4(n2035), .Y(n2085)
         );
  OA22X1_RVT U2781 ( .A1(n2085), .A2(n2448), .A3(n2063), .A4(n2465), .Y(n2028)
         );
  OA22X1_RVT U2782 ( .A1(n2043), .A2(n2467), .A3(n2026), .A4(n2456), .Y(n2027)
         );
  NAND2X0_RVT U2783 ( .A1(n2028), .A2(n2027), .Y(n2039) );
  AO22X1_RVT U2784 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2029), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2039), .Y(n2040) );
  AOI22X1_RVT U2785 ( .A1(n2176), .A2(n2040), .A3(a3stg_frac2[49]), .A4(n2526), 
        .Y(n2032) );
  NAND2X0_RVT U2786 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2030), .Y(n2031) );
  NAND3X0_RVT U2787 ( .A1(n2032), .A2(n2528), .A3(n2031), .Y(n2033) );
  HADDX1_RVT U2788 ( .A0(a2stg_sub_step), .B0(n2033), .SO(n1717) );
  OA22X1_RVT U2789 ( .A1(n2055), .A2(n2467), .A3(n2034), .A4(n2456), .Y(n2038)
         );
  OA22X1_RVT U2790 ( .A1(n2036), .A2(n2112), .A3(n2111), .A4(n2035), .Y(n2094)
         );
  OA22X1_RVT U2791 ( .A1(n2073), .A2(n2465), .A3(n2094), .A4(n2448), .Y(n2037)
         );
  NAND2X0_RVT U2792 ( .A1(n2038), .A2(n2037), .Y(n2048) );
  AO22X1_RVT U2793 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2039), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2048), .Y(n2049) );
  NAND2X0_RVT U2794 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2040), .Y(n2041) );
  NAND3X0_RVT U2795 ( .A1(n20), .A2(n2528), .A3(n2041), .Y(n2042) );
  HADDX1_RVT U2796 ( .A0(a2stg_sub_step), .B0(n2042), .SO(n1716) );
  OA22X1_RVT U2797 ( .A1(n2063), .A2(n2467), .A3(n2043), .A4(n2456), .Y(n2047)
         );
  AO22X1_RVT U2798 ( .A1(a2stg_frac2a[47]), .A2(n2045), .A3(a2stg_frac2a[63]), 
        .A4(n2044), .Y(n2122) );
  AOI22X1_RVT U2799 ( .A1(n2054), .A2(a2stg_frac2a[55]), .A3(n2449), .A4(n2122), .Y(n2102) );
  OA22X1_RVT U2800 ( .A1(n2102), .A2(n2448), .A3(n2085), .A4(n2465), .Y(n2046)
         );
  NAND2X0_RVT U2801 ( .A1(n2047), .A2(n2046), .Y(n2058) );
  AO22X1_RVT U2802 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2048), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2058), .Y(n2059) );
  AOI22X1_RVT U2803 ( .A1(n2176), .A2(n2059), .A3(a3stg_frac2[47]), .A4(n2526), 
        .Y(n2051) );
  NAND2X0_RVT U2804 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2049), .Y(n2050) );
  NAND3X0_RVT U2805 ( .A1(n2051), .A2(n2528), .A3(n2050), .Y(n2052) );
  HADDX1_RVT U2806 ( .A0(a2stg_sub_step), .B0(n2052), .SO(n1715) );
  AOI22X1_RVT U2807 ( .A1(n2054), .A2(a2stg_frac2a[54]), .A3(n2449), .A4(n2053), .Y(n2114) );
  OA22X1_RVT U2808 ( .A1(n2073), .A2(n2467), .A3(n2114), .A4(n2448), .Y(n2057)
         );
  OA22X1_RVT U2809 ( .A1(n2094), .A2(n2465), .A3(n2055), .A4(n2456), .Y(n2056)
         );
  NAND2X0_RVT U2810 ( .A1(n2057), .A2(n2056), .Y(n2068) );
  AO22X1_RVT U2811 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2058), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2068), .Y(n2069) );
  AOI22X1_RVT U2812 ( .A1(n2176), .A2(n2069), .A3(a3stg_frac2[46]), .A4(n2526), 
        .Y(n2061) );
  NAND2X0_RVT U2813 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2059), .Y(n2060) );
  NAND3X0_RVT U2814 ( .A1(n2061), .A2(n2528), .A3(n2060), .Y(n2062) );
  HADDX1_RVT U2815 ( .A0(a2stg_sub_step), .B0(n2062), .SO(n1714) );
  OA22X1_RVT U2816 ( .A1(n2085), .A2(n2467), .A3(n2063), .A4(n2456), .Y(n2067)
         );
  OA22X1_RVT U2817 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2065), .A3(n2112), .A4(
        n2064), .Y(n2123) );
  OA22X1_RVT U2818 ( .A1(n2102), .A2(n2465), .A3(n2123), .A4(n2448), .Y(n2066)
         );
  NAND2X0_RVT U2819 ( .A1(n2067), .A2(n2066), .Y(n2078) );
  AO22X1_RVT U2820 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2068), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2078), .Y(n2079) );
  AOI22X1_RVT U2821 ( .A1(n2176), .A2(n2079), .A3(a3stg_frac2[45]), .A4(n2526), 
        .Y(n2071) );
  NAND2X0_RVT U2822 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2069), .Y(n2070) );
  NAND3X0_RVT U2823 ( .A1(n2071), .A2(n2528), .A3(n2070), .Y(n2072) );
  HADDX1_RVT U2824 ( .A0(a2stg_sub_step), .B0(n2072), .SO(n1713) );
  OA22X1_RVT U2825 ( .A1(n2073), .A2(n2456), .A3(n2094), .A4(n2467), .Y(n2077)
         );
  OA22X1_RVT U2826 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2075), .A3(n2112), .A4(
        n2074), .Y(n2130) );
  OA22X1_RVT U2827 ( .A1(n2114), .A2(n2465), .A3(n2130), .A4(n2448), .Y(n2076)
         );
  NAND2X0_RVT U2828 ( .A1(n2077), .A2(n2076), .Y(n2088) );
  AO22X1_RVT U2829 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2078), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2088), .Y(n2089) );
  AOI22X1_RVT U2830 ( .A1(n2176), .A2(n2089), .A3(a3stg_frac2[44]), .A4(n2526), 
        .Y(n2081) );
  NAND2X0_RVT U2831 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2079), .Y(n2080) );
  NAND3X0_RVT U2832 ( .A1(n2081), .A2(n2528), .A3(n2080), .Y(n2082) );
  HADDX1_RVT U2833 ( .A0(a2stg_sub_step), .B0(n2082), .SO(n1712) );
  OA22X1_RVT U2834 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2084), .A3(n2112), .A4(
        n2083), .Y(n2137) );
  OA22X1_RVT U2835 ( .A1(n2123), .A2(n2465), .A3(n2137), .A4(n2448), .Y(n2087)
         );
  OA22X1_RVT U2836 ( .A1(n2102), .A2(n2467), .A3(n2085), .A4(n2456), .Y(n2086)
         );
  NAND2X0_RVT U2837 ( .A1(n2087), .A2(n2086), .Y(n2097) );
  AO22X1_RVT U2838 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2088), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2097), .Y(n2098) );
  NAND2X0_RVT U2839 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2089), .Y(n2090) );
  NAND3X0_RVT U2840 ( .A1(n21), .A2(n2528), .A3(n2090), .Y(n2091) );
  HADDX1_RVT U2841 ( .A0(a2stg_sub_step), .B0(n2091), .SO(n1711) );
  OA22X1_RVT U2842 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2093), .A3(n2112), .A4(
        n2092), .Y(n2144) );
  OA22X1_RVT U2843 ( .A1(n2130), .A2(n2465), .A3(n2144), .A4(n2448), .Y(n2096)
         );
  OA22X1_RVT U2844 ( .A1(n2094), .A2(n2456), .A3(n2114), .A4(n2467), .Y(n2095)
         );
  NAND2X0_RVT U2845 ( .A1(n2096), .A2(n2095), .Y(n2107) );
  AO22X1_RVT U2846 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2097), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2107), .Y(n2108) );
  AOI22X1_RVT U2847 ( .A1(n2176), .A2(n2108), .A3(a3stg_frac2[42]), .A4(n2526), 
        .Y(n2100) );
  NAND2X0_RVT U2848 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2098), .Y(n2099) );
  NAND3X0_RVT U2849 ( .A1(n2100), .A2(n2528), .A3(n2099), .Y(n2101) );
  HADDX1_RVT U2850 ( .A0(a2stg_sub_step), .B0(n2101), .SO(n1710) );
  OA22X1_RVT U2851 ( .A1(n2102), .A2(n2456), .A3(n2137), .A4(n2465), .Y(n2106)
         );
  OA22X1_RVT U2852 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2104), .A3(n2112), .A4(
        n2103), .Y(n2151) );
  OA22X1_RVT U2853 ( .A1(n2123), .A2(n2467), .A3(n2151), .A4(n2448), .Y(n2105)
         );
  NAND2X0_RVT U2854 ( .A1(n2106), .A2(n2105), .Y(n2117) );
  AO22X1_RVT U2855 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2107), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2117), .Y(n2118) );
  NAND2X0_RVT U2856 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2108), .Y(n2109) );
  NAND3X0_RVT U2857 ( .A1(n22), .A2(n2528), .A3(n2109), .Y(n2110) );
  HADDX1_RVT U2858 ( .A0(a2stg_sub_step), .B0(n2110), .SO(n1709) );
  OA22X1_RVT U2859 ( .A1(n2130), .A2(n2467), .A3(n2144), .A4(n2465), .Y(n2116)
         );
  OA22X1_RVT U2860 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2113), .A3(n2112), .A4(
        n2111), .Y(n2159) );
  OA22X1_RVT U2861 ( .A1(n2114), .A2(n2456), .A3(n2159), .A4(n2448), .Y(n2115)
         );
  NAND2X0_RVT U2862 ( .A1(n2116), .A2(n2115), .Y(n2126) );
  AO22X1_RVT U2863 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2117), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2126), .Y(n2127) );
  NAND2X0_RVT U2864 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2118), .Y(n2119) );
  NAND3X0_RVT U2865 ( .A1(n23), .A2(n2528), .A3(n2119), .Y(n2120) );
  HADDX1_RVT U2866 ( .A0(a2stg_sub_step), .B0(n2120), .SO(n1708) );
  AOI22X1_RVT U2867 ( .A1(a2stg_shr_cnt_3[1]), .A2(n2122), .A3(n2449), .A4(
        n2121), .Y(n2168) );
  OA22X1_RVT U2868 ( .A1(n2137), .A2(n2467), .A3(n2168), .A4(n2448), .Y(n2125)
         );
  OA22X1_RVT U2869 ( .A1(n2123), .A2(n2456), .A3(n2151), .A4(n2465), .Y(n2124)
         );
  NAND2X0_RVT U2870 ( .A1(n2125), .A2(n2124), .Y(n2133) );
  AO22X1_RVT U2871 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2126), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2133), .Y(n2134) );
  NAND2X0_RVT U2872 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2127), .Y(n2128) );
  NAND3X0_RVT U2873 ( .A1(n24), .A2(n2528), .A3(n2128), .Y(n2129) );
  HADDX1_RVT U2874 ( .A0(a2stg_sub_step), .B0(n2129), .SO(n1707) );
  OA22X1_RVT U2875 ( .A1(n2130), .A2(n2456), .A3(n2158), .A4(n2448), .Y(n2132)
         );
  OA22X1_RVT U2876 ( .A1(n2144), .A2(n2467), .A3(n2159), .A4(n2465), .Y(n2131)
         );
  NAND2X0_RVT U2877 ( .A1(n2132), .A2(n2131), .Y(n2140) );
  AO22X1_RVT U2878 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2133), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2140), .Y(n2141) );
  NAND2X0_RVT U2879 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2134), .Y(n2135) );
  NAND3X0_RVT U2880 ( .A1(n25), .A2(n2528), .A3(n2135), .Y(n2136) );
  HADDX1_RVT U2881 ( .A0(a2stg_sub_step), .B0(n2136), .SO(n1706) );
  OA22X1_RVT U2882 ( .A1(n2151), .A2(n2467), .A3(n2167), .A4(n2448), .Y(n2139)
         );
  OA22X1_RVT U2883 ( .A1(n2137), .A2(n2456), .A3(n2168), .A4(n2465), .Y(n2138)
         );
  NAND2X0_RVT U2884 ( .A1(n2139), .A2(n2138), .Y(n2147) );
  AO22X1_RVT U2885 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2140), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2147), .Y(n2148) );
  NAND2X0_RVT U2886 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2141), .Y(n2142) );
  NAND3X0_RVT U2887 ( .A1(n8), .A2(n2528), .A3(n2142), .Y(n2143) );
  HADDX1_RVT U2888 ( .A0(a2stg_sub_step), .B0(n2143), .SO(n1705) );
  OA22X1_RVT U2889 ( .A1(n2144), .A2(n2456), .A3(n2160), .A4(n2448), .Y(n2146)
         );
  OA22X1_RVT U2890 ( .A1(n2159), .A2(n2467), .A3(n2158), .A4(n2465), .Y(n2145)
         );
  NAND2X0_RVT U2891 ( .A1(n2146), .A2(n2145), .Y(n2154) );
  AO22X1_RVT U2892 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2147), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2154), .Y(n2155) );
  NAND2X0_RVT U2893 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2148), .Y(n2149) );
  NAND3X0_RVT U2894 ( .A1(n9), .A2(n2528), .A3(n2149), .Y(n2150) );
  HADDX1_RVT U2895 ( .A0(a2stg_sub_step), .B0(n2150), .SO(n1704) );
  OA22X1_RVT U2896 ( .A1(n2151), .A2(n2456), .A3(n2192), .A4(n2448), .Y(n2153)
         );
  OA22X1_RVT U2897 ( .A1(n2168), .A2(n2467), .A3(n2167), .A4(n2465), .Y(n2152)
         );
  NAND2X0_RVT U2898 ( .A1(n2153), .A2(n2152), .Y(n2163) );
  AO22X1_RVT U2899 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2154), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2163), .Y(n2164) );
  NAND2X0_RVT U2900 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2155), .Y(n2156) );
  NAND3X0_RVT U2901 ( .A1(n10), .A2(n2528), .A3(n2156), .Y(n2157) );
  HADDX1_RVT U2902 ( .A0(a2stg_sub_step), .B0(n2157), .SO(n1703) );
  OA22X1_RVT U2903 ( .A1(n2159), .A2(n2456), .A3(n2158), .A4(n2467), .Y(n2162)
         );
  OA22X1_RVT U2904 ( .A1(n2160), .A2(n2465), .A3(n2200), .A4(n2448), .Y(n2161)
         );
  NAND2X0_RVT U2905 ( .A1(n2162), .A2(n2161), .Y(n2171) );
  AO22X1_RVT U2906 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2163), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2171), .Y(n2172) );
  NAND2X0_RVT U2907 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2164), .Y(n2165) );
  NAND3X0_RVT U2908 ( .A1(n11), .A2(n2528), .A3(n2165), .Y(n2166) );
  HADDX1_RVT U2909 ( .A0(a2stg_sub_step), .B0(n2166), .SO(n1702) );
  OA22X1_RVT U2910 ( .A1(n2167), .A2(n2467), .A3(n2192), .A4(n2465), .Y(n2170)
         );
  OA22X1_RVT U2911 ( .A1(n2168), .A2(n2456), .A3(n2211), .A4(n2448), .Y(n2169)
         );
  NAND2X0_RVT U2912 ( .A1(n2170), .A2(n2169), .Y(n2175) );
  AO22X1_RVT U2913 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2171), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2175), .Y(n2177) );
  NAND2X0_RVT U2914 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2172), .Y(n2173) );
  NAND3X0_RVT U2915 ( .A1(n12), .A2(n2528), .A3(n2173), .Y(n2174) );
  HADDX1_RVT U2916 ( .A0(a2stg_sub_step), .B0(n2174), .SO(n1701) );
  AO22X1_RVT U2917 ( .A1(a2stg_shr_cnt_0[1]), .A2(n2175), .A3(
        a2stg_shr_cnt_0[0]), .A4(n2186), .Y(n2180) );
  NAND2X0_RVT U2918 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2177), .Y(n2178) );
  NAND3X0_RVT U2919 ( .A1(n13), .A2(n2528), .A3(n2178), .Y(n2179) );
  HADDX1_RVT U2920 ( .A0(a2stg_sub_step), .B0(n2179), .SO(n1700) );
  NAND3X0_RVT U2921 ( .A1(a2stg_expadd_11), .A2(a2stg_shr_frac2_shr_dbl), .A3(
        a2stg_shr_cnt_0[0]), .Y(n2387) );
  INVX1_RVT U2922 ( .A(n2387), .Y(n2525) );
  AOI22X1_RVT U2923 ( .A1(n2525), .A2(n2181), .A3(a2stg_shr_frac2_shr_int), 
        .A4(n2180), .Y(n2184) );
  NAND4X0_RVT U2924 ( .A1(a2stg_shr_frac2_shr_dbl), .A2(a2stg_expadd_11), .A3(
        a2stg_shr_cnt_0[1]), .A4(n2186), .Y(n2183) );
  NAND2X0_RVT U2925 ( .A1(a3stg_frac2[31]), .A2(n2526), .Y(n2182) );
  NAND4X0_RVT U2926 ( .A1(n2184), .A2(n2528), .A3(n2183), .A4(n2182), .Y(n2185) );
  HADDX1_RVT U2927 ( .A0(a2stg_sub_step), .B0(n2185), .SO(n1699) );
  AND3X1_RVT U2928 ( .A1(a2stg_expadd_11), .A2(a2stg_shr_frac2_shr_dbl), .A3(
        a2stg_shr_cnt_0[1]), .Y(n2523) );
  AO21X1_RVT U2929 ( .A1(a2stg_shr_cnt_0[0]), .A2(a2stg_shr_frac2_shr_int), 
        .A3(n2523), .Y(n2380) );
  INVX1_RVT U2930 ( .A(n2380), .Y(n2397) );
  OA22X1_RVT U2931 ( .A1(n2191), .A2(n2397), .A3(n2206), .A4(n2387), .Y(n2189)
         );
  NAND2X0_RVT U2932 ( .A1(a2stg_shr_cnt_0[1]), .A2(a2stg_shr_frac2_shr_int), 
        .Y(n2394) );
  INVX1_RVT U2933 ( .A(n2394), .Y(n2389) );
  NAND2X0_RVT U2934 ( .A1(n2389), .A2(n2186), .Y(n2188) );
  NAND2X0_RVT U2935 ( .A1(a3stg_frac2[30]), .A2(n2526), .Y(n2187) );
  NAND4X0_RVT U2936 ( .A1(n2189), .A2(n2528), .A3(n2188), .A4(n2187), .Y(n2190) );
  HADDX1_RVT U2937 ( .A0(a2stg_sub_step), .B0(n2190), .SO(n1698) );
  OA22X1_RVT U2938 ( .A1(n2206), .A2(n2397), .A3(n2191), .A4(n2394), .Y(n2197)
         );
  OA22X1_RVT U2939 ( .A1(n2192), .A2(n2456), .A3(n2211), .A4(n2467), .Y(n2194)
         );
  OA22X1_RVT U2940 ( .A1(n2227), .A2(n2465), .A3(n2244), .A4(n2448), .Y(n2193)
         );
  NAND2X0_RVT U2941 ( .A1(n2194), .A2(n2193), .Y(n2214) );
  NAND2X0_RVT U2942 ( .A1(n2525), .A2(n2214), .Y(n2196) );
  NAND2X0_RVT U2943 ( .A1(a3stg_frac2[29]), .A2(n2526), .Y(n2195) );
  NAND4X0_RVT U2944 ( .A1(n2197), .A2(n2528), .A3(n2196), .A4(n2195), .Y(n2198) );
  HADDX1_RVT U2945 ( .A0(a2stg_sub_step), .B0(n2198), .SO(n1697) );
  NAND2X0_RVT U2946 ( .A1(n2345), .A2(n2199), .Y(n2202) );
  OA22X1_RVT U2947 ( .A1(n2200), .A2(n2456), .A3(n2220), .A4(n2467), .Y(n2201)
         );
  AND2X1_RVT U2948 ( .A1(n2202), .A2(n2201), .Y(n2205) );
  NAND2X0_RVT U2949 ( .A1(n2203), .A2(n2450), .Y(n2204) );
  AND2X1_RVT U2950 ( .A1(n2205), .A2(n2204), .Y(n2219) );
  OA22X1_RVT U2951 ( .A1(n2206), .A2(n2394), .A3(n2219), .A4(n2387), .Y(n2209)
         );
  NAND2X0_RVT U2952 ( .A1(n2380), .A2(n2214), .Y(n2208) );
  NAND2X0_RVT U2953 ( .A1(a3stg_frac2[28]), .A2(n2526), .Y(n2207) );
  NAND4X0_RVT U2954 ( .A1(n2209), .A2(n2528), .A3(n2208), .A4(n2207), .Y(n2210) );
  HADDX1_RVT U2955 ( .A0(a2stg_sub_step), .B0(n2210), .SO(n1696) );
  OA22X1_RVT U2956 ( .A1(n2227), .A2(n2467), .A3(n2244), .A4(n2465), .Y(n2213)
         );
  OA22X1_RVT U2957 ( .A1(n2211), .A2(n2456), .A3(n2268), .A4(n2448), .Y(n2212)
         );
  AND2X1_RVT U2958 ( .A1(n2213), .A2(n2212), .Y(n2230) );
  OA22X1_RVT U2959 ( .A1(n2397), .A2(n2219), .A3(n2230), .A4(n2387), .Y(n2217)
         );
  NAND2X0_RVT U2960 ( .A1(n2389), .A2(n2214), .Y(n2216) );
  NAND2X0_RVT U2961 ( .A1(a3stg_frac2[27]), .A2(n2526), .Y(n2215) );
  NAND4X0_RVT U2962 ( .A1(n2217), .A2(n2528), .A3(n2216), .A4(n2215), .Y(n2218) );
  HADDX1_RVT U2963 ( .A0(a2stg_sub_step), .B0(n2218), .SO(n1695) );
  OA22X1_RVT U2964 ( .A1(n2397), .A2(n2230), .A3(n2219), .A4(n2394), .Y(n2225)
         );
  OA22X1_RVT U2965 ( .A1(n2256), .A2(n2465), .A3(n2278), .A4(n2448), .Y(n2222)
         );
  OA22X1_RVT U2966 ( .A1(n2220), .A2(n2456), .A3(n2235), .A4(n2467), .Y(n2221)
         );
  NAND2X0_RVT U2967 ( .A1(n2222), .A2(n2221), .Y(n2238) );
  NAND2X0_RVT U2968 ( .A1(n2525), .A2(n2238), .Y(n2224) );
  NAND2X0_RVT U2969 ( .A1(a3stg_frac2[26]), .A2(n2526), .Y(n2223) );
  NAND4X0_RVT U2970 ( .A1(n2225), .A2(n2528), .A3(n2224), .A4(n2223), .Y(n2226) );
  HADDX1_RVT U2971 ( .A0(a2stg_sub_step), .B0(n2226), .SO(n1694) );
  OA22X1_RVT U2972 ( .A1(n2227), .A2(n2456), .A3(n2244), .A4(n2467), .Y(n2229)
         );
  OA22X1_RVT U2973 ( .A1(n2268), .A2(n2465), .A3(n2287), .A4(n2448), .Y(n2228)
         );
  AND2X1_RVT U2974 ( .A1(n2229), .A2(n2228), .Y(n2243) );
  OA22X1_RVT U2975 ( .A1(n2230), .A2(n2394), .A3(n2243), .A4(n2387), .Y(n2233)
         );
  NAND2X0_RVT U2976 ( .A1(n2380), .A2(n2238), .Y(n2232) );
  NAND2X0_RVT U2977 ( .A1(a3stg_frac2[25]), .A2(n2526), .Y(n2231) );
  NAND4X0_RVT U2978 ( .A1(n2233), .A2(n2528), .A3(n2232), .A4(n2231), .Y(n2234) );
  HADDX1_RVT U2979 ( .A0(a2stg_sub_step), .B0(n2234), .SO(n1693) );
  OA22X1_RVT U2980 ( .A1(n2235), .A2(n2456), .A3(n2256), .A4(n2467), .Y(n2237)
         );
  OA22X1_RVT U2981 ( .A1(n2278), .A2(n2465), .A3(n2296), .A4(n2448), .Y(n2236)
         );
  AND2X1_RVT U2982 ( .A1(n2237), .A2(n2236), .Y(n2262) );
  OA22X1_RVT U2983 ( .A1(n2397), .A2(n2243), .A3(n2262), .A4(n2387), .Y(n2241)
         );
  NAND2X0_RVT U2984 ( .A1(n2389), .A2(n2238), .Y(n2240) );
  NAND2X0_RVT U2985 ( .A1(a3stg_frac2[24]), .A2(n2526), .Y(n2239) );
  NAND4X0_RVT U2986 ( .A1(n2241), .A2(n2528), .A3(n2240), .A4(n2239), .Y(n2242) );
  HADDX1_RVT U2987 ( .A0(a2stg_sub_step), .B0(n2242), .SO(n1692) );
  OA22X1_RVT U2988 ( .A1(n2397), .A2(n2262), .A3(n2243), .A4(n2394), .Y(n2251)
         );
  OA22X1_RVT U2989 ( .A1(n2244), .A2(n2456), .A3(n2287), .A4(n2465), .Y(n2248)
         );
  AOI22X1_RVT U2990 ( .A1(n2449), .A2(n2246), .A3(n2254), .A4(n2245), .Y(n2306) );
  OA22X1_RVT U2991 ( .A1(n2268), .A2(n2467), .A3(n2306), .A4(n2448), .Y(n2247)
         );
  NAND2X0_RVT U2992 ( .A1(n2248), .A2(n2247), .Y(n2271) );
  NAND2X0_RVT U2993 ( .A1(n2525), .A2(n2271), .Y(n2250) );
  NAND2X0_RVT U2994 ( .A1(a3stg_frac2[23]), .A2(n2526), .Y(n2249) );
  NAND4X0_RVT U2995 ( .A1(n2251), .A2(n2528), .A3(n2250), .A4(n2249), .Y(n2252) );
  HADDX1_RVT U2996 ( .A0(a2stg_sub_step), .B0(n2252), .SO(n1691) );
  AO22X1_RVT U2997 ( .A1(n2449), .A2(n2255), .A3(n2254), .A4(n2253), .Y(n2279)
         );
  NAND2X0_RVT U2998 ( .A1(n2450), .A2(n2279), .Y(n2258) );
  OA22X1_RVT U2999 ( .A1(n2256), .A2(n2456), .A3(n2296), .A4(n2465), .Y(n2257)
         );
  AND2X1_RVT U3000 ( .A1(n2258), .A2(n2257), .Y(n2261) );
  NAND2X0_RVT U3001 ( .A1(n2259), .A2(n2326), .Y(n2260) );
  AND2X1_RVT U3002 ( .A1(n2261), .A2(n2260), .Y(n2276) );
  OA22X1_RVT U3003 ( .A1(n2262), .A2(n2394), .A3(n2276), .A4(n2387), .Y(n2265)
         );
  NAND2X0_RVT U3004 ( .A1(n2380), .A2(n2271), .Y(n2264) );
  NAND2X0_RVT U3005 ( .A1(a3stg_frac2[22]), .A2(n2526), .Y(n2263) );
  NAND4X0_RVT U3006 ( .A1(n2265), .A2(n2528), .A3(n2264), .A4(n2263), .Y(n2266) );
  HADDX1_RVT U3007 ( .A0(a2stg_sub_step), .B0(n2266), .SO(n1690) );
  OA22X1_RVT U3008 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2349), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2267), .Y(n2323) );
  OA22X1_RVT U3009 ( .A1(n2306), .A2(n2465), .A3(n2323), .A4(n2448), .Y(n2270)
         );
  OA22X1_RVT U3010 ( .A1(n2268), .A2(n2456), .A3(n2287), .A4(n2467), .Y(n2269)
         );
  AND2X1_RVT U3011 ( .A1(n2270), .A2(n2269), .Y(n2290) );
  OA22X1_RVT U3012 ( .A1(n2397), .A2(n2276), .A3(n2290), .A4(n2387), .Y(n2274)
         );
  NAND2X0_RVT U3013 ( .A1(n2389), .A2(n2271), .Y(n2273) );
  NAND2X0_RVT U3014 ( .A1(a3stg_frac2[21]), .A2(n2526), .Y(n2272) );
  NAND4X0_RVT U3015 ( .A1(n2274), .A2(n2528), .A3(n2273), .A4(n2272), .Y(n2275) );
  HADDX1_RVT U3016 ( .A0(a2stg_sub_step), .B0(n2275), .SO(n1689) );
  OA22X1_RVT U3017 ( .A1(n2397), .A2(n2290), .A3(n2276), .A4(n2394), .Y(n2284)
         );
  OA22X1_RVT U3018 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2357), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2277), .Y(n2337) );
  OA22X1_RVT U3019 ( .A1(n2278), .A2(n2456), .A3(n2337), .A4(n2448), .Y(n2281)
         );
  INVX1_RVT U3020 ( .A(n2279), .Y(n2314) );
  OA22X1_RVT U3021 ( .A1(n2296), .A2(n2467), .A3(n2314), .A4(n2465), .Y(n2280)
         );
  NAND2X0_RVT U3022 ( .A1(n2281), .A2(n2280), .Y(n2299) );
  NAND2X0_RVT U3023 ( .A1(n2525), .A2(n2299), .Y(n2283) );
  NAND2X0_RVT U3024 ( .A1(a3stg_frac2[20]), .A2(n2526), .Y(n2282) );
  NAND4X0_RVT U3025 ( .A1(n2284), .A2(n2528), .A3(n2283), .A4(n2282), .Y(n2285) );
  HADDX1_RVT U3026 ( .A0(a2stg_sub_step), .B0(n2285), .SO(n1688) );
  OA22X1_RVT U3027 ( .A1(n2306), .A2(n2467), .A3(n2323), .A4(n2465), .Y(n2289)
         );
  OA22X1_RVT U3028 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2367), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2286), .Y(n2346) );
  OA22X1_RVT U3029 ( .A1(n2287), .A2(n2456), .A3(n2346), .A4(n2448), .Y(n2288)
         );
  AND2X1_RVT U3030 ( .A1(n2289), .A2(n2288), .Y(n2304) );
  OA22X1_RVT U3031 ( .A1(n2290), .A2(n2394), .A3(n2304), .A4(n2387), .Y(n2293)
         );
  NAND2X0_RVT U3032 ( .A1(n2380), .A2(n2299), .Y(n2292) );
  NAND2X0_RVT U3033 ( .A1(a3stg_frac2[19]), .A2(n2526), .Y(n2291) );
  NAND4X0_RVT U3034 ( .A1(n2293), .A2(n2528), .A3(n2292), .A4(n2291), .Y(n2294) );
  HADDX1_RVT U3035 ( .A0(a2stg_sub_step), .B0(n2294), .SO(n1687) );
  OA22X1_RVT U3036 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2375), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2295), .Y(n2358) );
  OA22X1_RVT U3037 ( .A1(n2337), .A2(n2465), .A3(n2358), .A4(n2448), .Y(n2298)
         );
  OA22X1_RVT U3038 ( .A1(n2296), .A2(n2456), .A3(n2314), .A4(n2467), .Y(n2297)
         );
  AND2X1_RVT U3039 ( .A1(n2298), .A2(n2297), .Y(n2317) );
  OA22X1_RVT U3040 ( .A1(n2397), .A2(n2304), .A3(n2317), .A4(n2387), .Y(n2302)
         );
  NAND2X0_RVT U3041 ( .A1(n2389), .A2(n2299), .Y(n2301) );
  NAND2X0_RVT U3042 ( .A1(a3stg_frac2[18]), .A2(n2526), .Y(n2300) );
  NAND4X0_RVT U3043 ( .A1(n2302), .A2(n2528), .A3(n2301), .A4(n2300), .Y(n2303) );
  HADDX1_RVT U3044 ( .A0(a2stg_sub_step), .B0(n2303), .SO(n1686) );
  OA22X1_RVT U3045 ( .A1(n2397), .A2(n2317), .A3(n2304), .A4(n2394), .Y(n2311)
         );
  OA22X1_RVT U3046 ( .A1(n2323), .A2(n2467), .A3(n2346), .A4(n2465), .Y(n2308)
         );
  OA22X1_RVT U3047 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2487), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2305), .Y(n2368) );
  OA22X1_RVT U3048 ( .A1(n2306), .A2(n2456), .A3(n2368), .A4(n2448), .Y(n2307)
         );
  NAND2X0_RVT U3049 ( .A1(n2308), .A2(n2307), .Y(n2330) );
  NAND2X0_RVT U3050 ( .A1(n2525), .A2(n2330), .Y(n2310) );
  NAND2X0_RVT U3051 ( .A1(a3stg_frac2[17]), .A2(n2526), .Y(n2309) );
  NAND4X0_RVT U3052 ( .A1(n2311), .A2(n2528), .A3(n2310), .A4(n2309), .Y(n2312) );
  HADDX1_RVT U3053 ( .A0(a2stg_sub_step), .B0(n2312), .SO(n1685) );
  OA22X1_RVT U3054 ( .A1(n2337), .A2(n2467), .A3(n2358), .A4(n2465), .Y(n2316)
         );
  OA22X1_RVT U3055 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2398), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2313), .Y(n2376) );
  OA22X1_RVT U3056 ( .A1(n2314), .A2(n2456), .A3(n2376), .A4(n2448), .Y(n2315)
         );
  AND2X1_RVT U3057 ( .A1(n2316), .A2(n2315), .Y(n2335) );
  OA22X1_RVT U3058 ( .A1(n2317), .A2(n2394), .A3(n2335), .A4(n2387), .Y(n2320)
         );
  NAND2X0_RVT U3059 ( .A1(n2380), .A2(n2330), .Y(n2319) );
  NAND2X0_RVT U3060 ( .A1(a3stg_frac2[16]), .A2(n2526), .Y(n2318) );
  NAND4X0_RVT U3061 ( .A1(n2320), .A2(n2528), .A3(n2319), .A4(n2318), .Y(n2321) );
  HADDX1_RVT U3062 ( .A0(a2stg_sub_step), .B0(n2321), .SO(n1684) );
  OA22X1_RVT U3063 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2410), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2322), .Y(n2502) );
  INVX1_RVT U3064 ( .A(n2502), .Y(n2344) );
  NAND2X0_RVT U3065 ( .A1(n2450), .A2(n2344), .Y(n2325) );
  OA22X1_RVT U3066 ( .A1(n2323), .A2(n2456), .A3(n2368), .A4(n2465), .Y(n2324)
         );
  AND2X1_RVT U3067 ( .A1(n2325), .A2(n2324), .Y(n2329) );
  NAND2X0_RVT U3068 ( .A1(n2327), .A2(n2326), .Y(n2328) );
  AND2X1_RVT U3069 ( .A1(n2329), .A2(n2328), .Y(n2352) );
  OA22X1_RVT U3070 ( .A1(n2397), .A2(n2335), .A3(n2352), .A4(n2387), .Y(n2333)
         );
  NAND2X0_RVT U3071 ( .A1(n2389), .A2(n2330), .Y(n2332) );
  NAND2X0_RVT U3072 ( .A1(a3stg_frac2[15]), .A2(n2526), .Y(n2331) );
  NAND4X0_RVT U3073 ( .A1(n2333), .A2(n2528), .A3(n2332), .A4(n2331), .Y(n2334) );
  HADDX1_RVT U3074 ( .A0(a2stg_sub_step), .B0(n2334), .SO(n1683) );
  OA22X1_RVT U3075 ( .A1(n2397), .A2(n2352), .A3(n2335), .A4(n2394), .Y(n2342)
         );
  OA22X1_RVT U3076 ( .A1(n2358), .A2(n2467), .A3(n2376), .A4(n2465), .Y(n2339)
         );
  OA22X1_RVT U3077 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2405), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2336), .Y(n2501) );
  OA22X1_RVT U3078 ( .A1(n2501), .A2(n2448), .A3(n2337), .A4(n2456), .Y(n2338)
         );
  NAND2X0_RVT U3079 ( .A1(n2339), .A2(n2338), .Y(n2361) );
  NAND2X0_RVT U3080 ( .A1(n2525), .A2(n2361), .Y(n2341) );
  NAND2X0_RVT U3081 ( .A1(a3stg_frac2[14]), .A2(n2526), .Y(n2340) );
  NAND4X0_RVT U3082 ( .A1(n2342), .A2(n2528), .A3(n2341), .A4(n2340), .Y(n2343) );
  HADDX1_RVT U3083 ( .A0(a2stg_sub_step), .B0(n2343), .SO(n1682) );
  NAND2X0_RVT U3084 ( .A1(n2345), .A2(n2344), .Y(n2348) );
  OA22X1_RVT U3085 ( .A1(n2346), .A2(n2456), .A3(n2368), .A4(n2467), .Y(n2347)
         );
  AND2X1_RVT U3086 ( .A1(n2348), .A2(n2347), .Y(n2351) );
  OA22X1_RVT U3087 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2416), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2349), .Y(n2409) );
  INVX1_RVT U3088 ( .A(n2409), .Y(n2505) );
  NAND2X0_RVT U3089 ( .A1(n2505), .A2(n2450), .Y(n2350) );
  AND2X1_RVT U3090 ( .A1(n2351), .A2(n2350), .Y(n2366) );
  OA22X1_RVT U3091 ( .A1(n2352), .A2(n2394), .A3(n2366), .A4(n2387), .Y(n2355)
         );
  NAND2X0_RVT U3092 ( .A1(n2380), .A2(n2361), .Y(n2354) );
  NAND2X0_RVT U3093 ( .A1(a3stg_frac2[13]), .A2(n2526), .Y(n2353) );
  NAND4X0_RVT U3094 ( .A1(n2355), .A2(n2528), .A3(n2354), .A4(n2353), .Y(n2356) );
  HADDX1_RVT U3095 ( .A0(a2stg_sub_step), .B0(n2356), .SO(n1681) );
  OA22X1_RVT U3096 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2424), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2357), .Y(n2510) );
  OA22X1_RVT U3097 ( .A1(n2510), .A2(n2448), .A3(n2501), .A4(n2465), .Y(n2360)
         );
  OA22X1_RVT U3098 ( .A1(n2358), .A2(n2456), .A3(n2376), .A4(n2467), .Y(n2359)
         );
  AND2X1_RVT U3099 ( .A1(n2360), .A2(n2359), .Y(n2379) );
  OA22X1_RVT U3100 ( .A1(n2397), .A2(n2366), .A3(n2379), .A4(n2387), .Y(n2364)
         );
  NAND2X0_RVT U3101 ( .A1(n2389), .A2(n2361), .Y(n2363) );
  NAND2X0_RVT U3102 ( .A1(a3stg_frac2[12]), .A2(n2526), .Y(n2362) );
  NAND4X0_RVT U3103 ( .A1(n2364), .A2(n2528), .A3(n2363), .A4(n2362), .Y(n2365) );
  HADDX1_RVT U3104 ( .A0(a2stg_sub_step), .B0(n2365), .SO(n1680) );
  OA22X1_RVT U3105 ( .A1(n2397), .A2(n2379), .A3(n2366), .A4(n2394), .Y(n2373)
         );
  OA22X1_RVT U3106 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2432), .A3(
        a2stg_shr_cnt_3[2]), .A4(n2367), .Y(n2418) );
  OA22X1_RVT U3107 ( .A1(n2418), .A2(n2448), .A3(n2368), .A4(n2456), .Y(n2370)
         );
  OA22X1_RVT U3108 ( .A1(n2409), .A2(n2465), .A3(n2502), .A4(n2467), .Y(n2369)
         );
  NAND2X0_RVT U3109 ( .A1(n2370), .A2(n2369), .Y(n2388) );
  NAND2X0_RVT U3110 ( .A1(n2525), .A2(n2388), .Y(n2372) );
  NAND2X0_RVT U3111 ( .A1(a3stg_frac2[11]), .A2(n2526), .Y(n2371) );
  NAND4X0_RVT U3112 ( .A1(n2373), .A2(n2528), .A3(n2372), .A4(n2371), .Y(n2374) );
  HADDX1_RVT U3113 ( .A0(a2stg_sub_step), .B0(n2374), .SO(n1679) );
  OA22X1_RVT U3114 ( .A1(n2510), .A2(n2465), .A3(n2501), .A4(n2467), .Y(n2378)
         );
  OA22X1_RVT U3115 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2441), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2375), .Y(n2426) );
  OA22X1_RVT U3116 ( .A1(n2426), .A2(n2448), .A3(n2376), .A4(n2456), .Y(n2377)
         );
  AND2X1_RVT U3117 ( .A1(n2378), .A2(n2377), .Y(n2395) );
  OA22X1_RVT U3118 ( .A1(n2379), .A2(n2394), .A3(n2395), .A4(n2387), .Y(n2383)
         );
  NAND2X0_RVT U3119 ( .A1(n2380), .A2(n2388), .Y(n2382) );
  NAND2X0_RVT U3120 ( .A1(a3stg_frac2[10]), .A2(n2526), .Y(n2381) );
  NAND4X0_RVT U3121 ( .A1(n2383), .A2(n2528), .A3(n2382), .A4(n2381), .Y(n2384) );
  HADDX1_RVT U3122 ( .A0(a2stg_sub_step), .B0(n2384), .SO(n1678) );
  OA22X1_RVT U3123 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2452), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2487), .Y(n2434) );
  OA22X1_RVT U3124 ( .A1(n2434), .A2(n2448), .A3(n2502), .A4(n2456), .Y(n2386)
         );
  OA22X1_RVT U3125 ( .A1(n2418), .A2(n2465), .A3(n2409), .A4(n2467), .Y(n2385)
         );
  AND2X1_RVT U3126 ( .A1(n2386), .A2(n2385), .Y(n2396) );
  OA22X1_RVT U3127 ( .A1(n2397), .A2(n2395), .A3(n2396), .A4(n2387), .Y(n2392)
         );
  NAND2X0_RVT U3128 ( .A1(n2389), .A2(n2388), .Y(n2391) );
  NAND2X0_RVT U3129 ( .A1(a3stg_frac2[9]), .A2(n2526), .Y(n2390) );
  NAND4X0_RVT U3130 ( .A1(n2392), .A2(n2528), .A3(n2391), .A4(n2390), .Y(n2393) );
  HADDX1_RVT U3131 ( .A0(a2stg_sub_step), .B0(n2393), .SO(n1677) );
  OA22X1_RVT U3132 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .Y(n2403)
         );
  OA22X1_RVT U3133 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2472), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2398), .Y(n2440) );
  OA22X1_RVT U3134 ( .A1(n2501), .A2(n2456), .A3(n2440), .A4(n2448), .Y(n2400)
         );
  OA22X1_RVT U3135 ( .A1(n2510), .A2(n2467), .A3(n2426), .A4(n2465), .Y(n2399)
         );
  NAND2X0_RVT U3136 ( .A1(n2400), .A2(n2399), .Y(n2522) );
  NAND2X0_RVT U3137 ( .A1(n2525), .A2(n2522), .Y(n2402) );
  NAND2X0_RVT U3138 ( .A1(a3stg_frac2[8]), .A2(n2526), .Y(n2401) );
  NAND4X0_RVT U3139 ( .A1(n2403), .A2(n2528), .A3(n2402), .A4(n2401), .Y(n2404) );
  HADDX1_RVT U3140 ( .A0(a2stg_sub_step), .B0(n2404), .SO(n1676) );
  OA22X1_RVT U3141 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2406), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2405), .Y(n2475) );
  OA22X1_RVT U3142 ( .A1(n2426), .A2(n2467), .A3(n2475), .A4(n2448), .Y(n2408)
         );
  OA22X1_RVT U3143 ( .A1(n2510), .A2(n2456), .A3(n2440), .A4(n2465), .Y(n2407)
         );
  NAND2X0_RVT U3144 ( .A1(n2408), .A2(n2407), .Y(n2421) );
  OA22X1_RVT U3145 ( .A1(n2418), .A2(n2467), .A3(n2409), .A4(n2456), .Y(n2413)
         );
  OA22X1_RVT U3146 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2411), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2410), .Y(n2455) );
  OA22X1_RVT U3147 ( .A1(n2434), .A2(n2465), .A3(n2455), .A4(n2448), .Y(n2412)
         );
  NAND2X0_RVT U3148 ( .A1(n2413), .A2(n2412), .Y(n2524) );
  NAND2X0_RVT U3149 ( .A1(n2523), .A2(n2524), .Y(n2414) );
  NAND3X0_RVT U3150 ( .A1(n14), .A2(n2528), .A3(n2414), .Y(n2415) );
  HADDX1_RVT U3151 ( .A0(a2stg_sub_step), .B0(n2415), .SO(n1675) );
  OA22X1_RVT U3152 ( .A1(n2434), .A2(n2467), .A3(n2455), .A4(n2465), .Y(n2420)
         );
  OA22X1_RVT U3153 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2417), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2416), .Y(n2454) );
  OA22X1_RVT U3154 ( .A1(n2418), .A2(n2456), .A3(n2454), .A4(n2448), .Y(n2419)
         );
  NAND2X0_RVT U3155 ( .A1(n2420), .A2(n2419), .Y(n2429) );
  NAND2X0_RVT U3156 ( .A1(n2523), .A2(n2421), .Y(n2422) );
  NAND3X0_RVT U3157 ( .A1(n15), .A2(n2528), .A3(n2422), .Y(n2423) );
  HADDX1_RVT U3158 ( .A0(a2stg_sub_step), .B0(n2423), .SO(n1674) );
  OA22X1_RVT U3159 ( .A1(n2440), .A2(n2467), .A3(n2475), .A4(n2465), .Y(n2428)
         );
  OA22X1_RVT U3160 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2425), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2424), .Y(n2468) );
  OA22X1_RVT U3161 ( .A1(n2426), .A2(n2456), .A3(n2468), .A4(n2448), .Y(n2427)
         );
  NAND2X0_RVT U3162 ( .A1(n2428), .A2(n2427), .Y(n2437) );
  NAND2X0_RVT U3163 ( .A1(n2523), .A2(n2429), .Y(n2430) );
  NAND3X0_RVT U3164 ( .A1(n16), .A2(n2528), .A3(n2430), .Y(n2431) );
  HADDX1_RVT U3165 ( .A0(a2stg_sub_step), .B0(n2431), .SO(n1673) );
  OA22X1_RVT U3166 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2433), .A3(
        a2stg_shr_cnt_3[3]), .A4(n2432), .Y(n2453) );
  OA22X1_RVT U3167 ( .A1(n2454), .A2(n2465), .A3(n2453), .A4(n2448), .Y(n2436)
         );
  OA22X1_RVT U3168 ( .A1(n2434), .A2(n2456), .A3(n2455), .A4(n2467), .Y(n2435)
         );
  NAND2X0_RVT U3169 ( .A1(n2436), .A2(n2435), .Y(n2445) );
  NAND2X0_RVT U3170 ( .A1(n2523), .A2(n2437), .Y(n2438) );
  NAND3X0_RVT U3171 ( .A1(n17), .A2(n2528), .A3(n2438), .Y(n2439) );
  HADDX1_RVT U3172 ( .A0(a2stg_sub_step), .B0(n2439), .SO(n1672) );
  OA22X1_RVT U3173 ( .A1(n2440), .A2(n2456), .A3(n2475), .A4(n2467), .Y(n2444)
         );
  OA22X1_RVT U3174 ( .A1(a2stg_shr_cnt_3[4]), .A2(n2442), .A3(n2441), .A4(
        a2stg_shr_cnt_3[3]), .Y(n2466) );
  OA22X1_RVT U3175 ( .A1(n2468), .A2(n2465), .A3(n2466), .A4(n2448), .Y(n2443)
         );
  NAND2X0_RVT U3176 ( .A1(n2444), .A2(n2443), .Y(n2460) );
  NAND2X0_RVT U3177 ( .A1(n2523), .A2(n2445), .Y(n2446) );
  NAND3X0_RVT U3178 ( .A1(n18), .A2(n2528), .A3(n2446), .Y(n2447) );
  HADDX1_RVT U3179 ( .A0(a2stg_sub_step), .B0(n2447), .SO(n1671) );
  OR2X1_RVT U3180 ( .A1(n2448), .A2(a2stg_shr_cnt_3[3]), .Y(n2471) );
  NAND2X0_RVT U3181 ( .A1(n2450), .A2(n2449), .Y(n2469) );
  OA22X1_RVT U3182 ( .A1(n2452), .A2(n2471), .A3(n2451), .A4(n2469), .Y(n2459)
         );
  OA22X1_RVT U3183 ( .A1(n2454), .A2(n2467), .A3(n2453), .A4(n2465), .Y(n2458)
         );
  OR2X1_RVT U3184 ( .A1(n2456), .A2(n2455), .Y(n2457) );
  NAND3X0_RVT U3185 ( .A1(n2459), .A2(n2458), .A3(n2457), .Y(n2463) );
  NAND2X0_RVT U3186 ( .A1(n2523), .A2(n2460), .Y(n2461) );
  NAND3X0_RVT U3187 ( .A1(n19), .A2(n2528), .A3(n2461), .Y(n2462) );
  HADDX1_RVT U3188 ( .A0(a2stg_sub_step), .B0(n2462), .SO(n1670) );
  AOI22X1_RVT U3189 ( .A1(n2523), .A2(n2463), .A3(a3stg_frac2[0]), .A4(n2526), 
        .Y(n2464) );
  AND2X1_RVT U3190 ( .A1(n2528), .A2(n2464), .Y(n2482) );
  OA22X1_RVT U3191 ( .A1(n2468), .A2(n2467), .A3(n2466), .A4(n2465), .Y(n2474)
         );
  OA22X1_RVT U3192 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .Y(n2473)
         );
  AND2X1_RVT U3193 ( .A1(n2474), .A2(n2473), .Y(n2479) );
  NAND2X0_RVT U3194 ( .A1(n2477), .A2(n2476), .Y(n2478) );
  NAND2X0_RVT U3195 ( .A1(n2479), .A2(n2478), .Y(n2480) );
  NAND2X0_RVT U3196 ( .A1(n2480), .A2(n2525), .Y(n2481) );
  AND2X1_RVT U3197 ( .A1(n2482), .A2(n2481), .Y(n2484) );
  HADDX1_RVT U3198 ( .A0(n2484), .B0(n2483), .SO(n1669) );
  AO22X1_RVT U3199 ( .A1(a2stg_shr_cnt[3]), .A2(n2487), .A3(n2486), .A4(n2485), 
        .Y(n2508) );
  AOI22X1_RVT U3200 ( .A1(a2stg_shr_cnt[3]), .A2(n2489), .A3(n2504), .A4(n2488), .Y(n2514) );
  NAND2X0_RVT U3201 ( .A1(a2stg_shr_cnt[3]), .A2(n2491), .Y(n2492) );
  AND2X1_RVT U3202 ( .A1(n2493), .A2(n2492), .Y(n2497) );
  NAND2X0_RVT U3203 ( .A1(a2stg_shr_cnt[3]), .A2(n2494), .Y(n2495) );
  NAND3X0_RVT U3204 ( .A1(n2496), .A2(n2497), .A3(n2495), .Y(n2500) );
  AND2X1_RVT U3205 ( .A1(n2500), .A2(a2stg_shr_cnt[1]), .Y(n2499) );
  NAND2X0_RVT U3206 ( .A1(n2503), .A2(n2497), .Y(n2498) );
  NAND2X0_RVT U3207 ( .A1(n2499), .A2(n2498), .Y(n2513) );
  OAI21X1_RVT U3208 ( .A1(n2503), .A2(n2502), .A3(n2501), .Y(n2506) );
  AOI22X1_RVT U3209 ( .A1(a2stg_shr_cnt[1]), .A2(n2506), .A3(n2505), .A4(n2504), .Y(n2507) );
  NAND4X0_RVT U3210 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .Y(n2511) );
  NAND2X0_RVT U3211 ( .A1(a2stg_shr_cnt[2]), .A2(n2511), .Y(n2512) );
  NAND3X0_RVT U3212 ( .A1(n2514), .A2(n2513), .A3(n2512), .Y(n2532) );
  NOR4X1_RVT U3213 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .Y(n2519)
         );
  NAND3X0_RVT U3214 ( .A1(n2521), .A2(n2520), .A3(n2519), .Y(n2531) );
  AOI22X1_RVT U3215 ( .A1(n2525), .A2(n2524), .A3(n2523), .A4(n2522), .Y(n2529) );
  NAND2X0_RVT U3216 ( .A1(a3stg_frac2[7]), .A2(n2526), .Y(n2527) );
  NAND3X0_RVT U3217 ( .A1(n2529), .A2(n2528), .A3(n2527), .Y(n2530) );
  AO221X1_RVT U3218 ( .A1(a2stg_shr_frac2_shr_int), .A2(n2532), .A3(
        a2stg_shr_frac2_shr_int), .A4(n2531), .A5(n2530), .Y(n2533) );
  HADDX1_RVT U3219 ( .A0(a2stg_sub_step), .B0(n2533), .SO(n1668) );
endmodule


module fpu_add ( inq_op, inq_rnd_mode, inq_id, inq_fcc, inq_in1, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, fadd_clken_l, arst_l, 
        grst_l, rclk, add_pipe_active, a1stg_step, a6stg_fadd_in, 
        add_id_out_in, a6stg_fcmpop, add_exc_out, a6stg_dbl_dst, a6stg_sng_dst, 
        a6stg_long_dst, a6stg_int_dst, add_sign_out, add_exp_out, add_frac_out, 
        add_cc_out, add_fcc_out, se_add_exp, se_add_frac, si, so, 
        add_dest_rdy_BAR );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [1:0] inq_fcc;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] add_id_out_in;
  output [4:0] add_exc_out;
  output [10:0] add_exp_out;
  output [63:0] add_frac_out;
  output [1:0] add_cc_out;
  output [1:0] add_fcc_out;
  input inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0,
         inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0,
         inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, fadd_clken_l, arst_l,
         grst_l, rclk, se_add_exp, se_add_frac, si, add_dest_rdy_BAR;
  output add_pipe_active, a1stg_step, a6stg_fadd_in, a6stg_fcmpop,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         add_sign_out, so;
  wire   add_dest_rdy, a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac,
         a1stg_in2_eq_in1_exp, a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0,
         a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a2stg_frac2_63, add_of_out_cout,
         a4stg_frac_neq_0, a4stg_shl_data_neq_0, a4stg_frac_dbl_nx,
         a4stg_frac_sng_nx, a3stg_denorm, a4stg_denorm_inv, a4stg_round,
         a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac_11,
         a4stg_rnd_frac_10, a4stg_frac_38_0_nx, a4stg_frac_9_0_nx,
         a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1, a1stg_denorm_sng_in2,
         a1stg_denorm_dbl_in2, a1stg_norm_sng_in1, a1stg_norm_dbl_in1,
         a1stg_norm_sng_in2, a1stg_norm_dbl_in2, a1stg_stepa, a1stg_sngop,
         a1stg_intlngop, a1stg_fsdtoix, a1stg_fstod, a1stg_fstoi, a1stg_fstox,
         a1stg_fdtoi, a1stg_fdtox, a1stg_faddsubs, a1stg_faddsubd, a1stg_fdtos,
         a2stg_faddsubop, a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod,
         a2stg_fxtos, a2stg_fxtod, a3stg_faddsubop, a4stg_dblop, a6stg_step,
         a3stg_sub_in, a4stg_in_of, a2stg_frac1_in_frac1, a2stg_frac1_in_frac2,
         a1stg_2nan_in_inv, a1stg_faddsubop_inv, a2stg_frac1_in_qnan,
         a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, a2stg_frac2_in_frac1,
         a2stg_frac2_in_qnan, a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add,
         a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0,
         a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1,
         add_exp_out_expadd, a4stg_to_0_inv, a3stg_inc_exp_inv,
         a3stg_same_exp_inv, a3stg_dec_exp_inv, a4stg_rndadd_cout,
         a1stg_expadd3_11, net211161, net211162, net211163, net211164;
  wire   [11:0] a1stg_expadd1_11_0;
  wire   [12:0] a2stg_expadd;
  wire   [11:0] a2stg_exp;
  wire   [11:0] a4stg_exp_11_0;
  wire   [5:0] a1stg_expadd2_5_0;
  wire   [10:0] a1stg_expadd4_inv;
  wire   [10:0] a3stg_exp_10_0;
  wire   [5:0] a3stg_lead0;
  wire   [1:0] a3stg_faddsubopa;
  wire   [5:0] a2stg_shr_cnt_in;
  wire   [9:0] a4stg_shl_cnt_in;
  wire   [5:0] a4stg_shl_cnt;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign add_dest_rdy = add_dest_rdy_BAR;

  fpu_add_ctl fpu_add_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_63(inq_in1[63]), .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(inq_in1_exp_neq_ffs), 
        .inq_in2_51(inq_in2[51]), .inq_in2_54(inq_in2[54]), .inq_in2_63(
        inq_in2[63]), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0), .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(
        inq_op), .inq_rnd_mode(inq_rnd_mode), .inq_id(inq_id), .inq_fcc(
        inq_fcc), .inq_add(inq_add), .a1stg_in2_neq_in1_frac(
        a1stg_in2_neq_in1_frac), .a1stg_in2_gt_in1_frac(a1stg_in2_gt_in1_frac), 
        .a1stg_in2_eq_in1_exp(a1stg_in2_eq_in1_exp), .a1stg_expadd1(
        a1stg_expadd1_11_0), .a2stg_expadd(a2stg_expadd[11:0]), 
        .a2stg_frac2hi_neq_0(a2stg_frac2hi_neq_0), .a2stg_frac2lo_neq_0(
        a2stg_frac2lo_neq_0), .a2stg_exp(a2stg_exp), .a3stg_fsdtoix_nx(
        a3stg_fsdtoix_nx), .a3stg_fsdtoi_nx(a3stg_fsdtoi_nx), .a2stg_frac2_63(
        a2stg_frac2_63), .a4stg_exp(a4stg_exp_11_0), .add_of_out_cout(
        add_of_out_cout), .a4stg_frac_neq_0(a4stg_frac_neq_0), 
        .a4stg_shl_data_neq_0(a4stg_shl_data_neq_0), .a4stg_frac_dbl_nx(
        a4stg_frac_dbl_nx), .a4stg_frac_sng_nx(a4stg_frac_sng_nx), 
        .a1stg_expadd2(a1stg_expadd2_5_0), .a1stg_expadd4_inv(
        a1stg_expadd4_inv), .a3stg_denorm(a3stg_denorm), .a3stg_denorm_inv(
        net211163), .a4stg_denorm_inv(a4stg_denorm_inv), .a3stg_exp(
        a3stg_exp_10_0), .a3stg_lead0(a3stg_lead0), .a4stg_rnd_frac_40(
        a4stg_rnd_frac_40), .a4stg_rnd_frac_39(a4stg_rnd_frac_39), 
        .a4stg_rnd_frac_11(a4stg_rnd_frac_11), .a4stg_rnd_frac_10(
        a4stg_rnd_frac_10), .a4stg_frac_38_0_nx(a4stg_frac_38_0_nx), 
        .a4stg_frac_9_0_nx(a4stg_frac_9_0_nx), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), .add_pipe_active(add_pipe_active), .a1stg_denorm_sng_in1(
        a1stg_denorm_sng_in1), .a1stg_denorm_dbl_in1(a1stg_denorm_dbl_in1), 
        .a1stg_denorm_sng_in2(a1stg_denorm_sng_in2), .a1stg_denorm_dbl_in2(
        a1stg_denorm_dbl_in2), .a1stg_norm_sng_in1(a1stg_norm_sng_in1), 
        .a1stg_norm_dbl_in1(a1stg_norm_dbl_in1), .a1stg_norm_sng_in2(
        a1stg_norm_sng_in2), .a1stg_norm_dbl_in2(a1stg_norm_dbl_in2), 
        .a1stg_step(a1stg_step), .a1stg_stepa(a1stg_stepa), .a1stg_sngop(
        a1stg_sngop), .a1stg_intlngop(a1stg_intlngop), .a1stg_fsdtoix(
        a1stg_fsdtoix), .a1stg_fstod(a1stg_fstod), .a1stg_fstoi(a1stg_fstoi), 
        .a1stg_fstox(a1stg_fstox), .a1stg_fdtoi(a1stg_fdtoi), .a1stg_fdtox(
        a1stg_fdtox), .a1stg_faddsubs(a1stg_faddsubs), .a1stg_faddsubd(
        a1stg_faddsubd), .a1stg_fdtos(a1stg_fdtos), .a2stg_faddsubop(
        a2stg_faddsubop), .a2stg_fsdtoix_fdtos(a2stg_fsdtoix_fdtos), 
        .a2stg_fitos(a2stg_fitos), .a2stg_fitod(a2stg_fitod), .a2stg_fxtos(
        a2stg_fxtos), .a2stg_fxtod(a2stg_fxtod), .a3stg_faddsubop(
        a3stg_faddsubop), .a3stg_faddsubopa(a3stg_faddsubopa), .a4stg_dblop(
        a4stg_dblop), .a6stg_fadd_in(a6stg_fadd_in), .add_id_out_in(
        add_id_out_in), .add_fcc_out(add_fcc_out), .a6stg_dbl_dst(
        a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), .a6stg_long_dst(
        a6stg_long_dst), .a6stg_int_dst(a6stg_int_dst), .a6stg_fcmpop(
        a6stg_fcmpop), .a6stg_step(a6stg_step), .a3stg_sub_in(a3stg_sub_in), 
        .add_sign_out(add_sign_out), .add_cc_out(add_cc_out), .a4stg_in_of(
        a4stg_in_of), .add_exc_out({add_exc_out[4:2], SYNOPSYS_UNCONNECTED__0, 
        add_exc_out[0]}), .a2stg_frac1_in_frac1(a2stg_frac1_in_frac1), 
        .a2stg_frac1_in_frac2(a2stg_frac1_in_frac2), .a1stg_2nan_in_inv(
        a1stg_2nan_in_inv), .a1stg_faddsubop_inv(a1stg_faddsubop_inv), 
        .a2stg_frac1_in_qnan(a2stg_frac1_in_qnan), .a2stg_frac1_in_nv(
        a2stg_frac1_in_nv), .a2stg_frac1_in_nv_dbl(a2stg_frac1_in_nv_dbl), 
        .a2stg_frac2_in_frac1(a2stg_frac2_in_frac1), .a2stg_frac2_in_qnan(
        a2stg_frac2_in_qnan), .a2stg_shr_cnt_in(a2stg_shr_cnt_in), 
        .a2stg_shr_cnt_5_inv_in(a2stg_shr_cnt_5_inv_in), 
        .a2stg_shr_frac2_shr_int(a2stg_shr_frac2_shr_int), 
        .a2stg_shr_frac2_shr_dbl(a2stg_shr_frac2_shr_dbl), 
        .a2stg_shr_frac2_shr_sng(a2stg_shr_frac2_shr_sng), 
        .a2stg_shr_frac2_max(a2stg_shr_frac2_max), .a2stg_sub_step(
        a2stg_sub_step), .a2stg_fracadd_frac2_inv_in(
        a2stg_fracadd_frac2_inv_in), .a2stg_fracadd_frac2_inv_shr1_in(
        a2stg_fracadd_frac2_inv_shr1_in), .a2stg_fracadd_frac2(
        a2stg_fracadd_frac2), .a2stg_fracadd_cin_in(a2stg_fracadd_cin_in), 
        .a3stg_exp_7ff(a3stg_exp_7ff), .a3stg_exp_ff(a3stg_exp_ff), 
        .a3stg_exp_add(a3stg_exp_add), .a2stg_expdec_neq_0(a2stg_expdec_neq_0), 
        .a3stg_exp10_0_eq0(a3stg_exp10_0_eq0), .a3stg_exp10_1_eq0(
        a3stg_exp10_1_eq0), .a3stg_fdtos_inv(a3stg_fdtos_inv), 
        .a4stg_fixtos_fxtod_inv(a4stg_fixtos_fxtod_inv), 
        .a4stg_rnd_frac_add_inv(a4stg_rnd_frac_add_inv), .a4stg_shl_cnt_in(
        a4stg_shl_cnt_in), .a4stg_rnd_sng(a4stg_rnd_sng), .a4stg_rnd_dbl(
        a4stg_rnd_dbl), .add_frac_out_rndadd(add_frac_out_rndadd), 
        .add_frac_out_rnd_frac(add_frac_out_rnd_frac), .add_frac_out_shl(
        add_frac_out_shl), .a4stg_to_0(a4stg_to_0), .add_exp_out_expinc(
        add_exp_out_expinc), .add_exp_out_exp(add_exp_out_exp), 
        .add_exp_out_exp1(add_exp_out_exp1), .add_exp_out_expadd(
        add_exp_out_expadd), .a4stg_to_0_inv(a4stg_to_0_inv), .se(se_add_exp), 
        .si(net211164), .add_dest_rdy_BAR(add_dest_rdy), .a4stg_round_BAR(
        a4stg_round) );
  fpu_add_exp_dp fpu_add_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .inq_op(inq_op[1:0]), .inq_op_7(inq_op[7]), 
        .a1stg_step(a1stg_stepa), .a1stg_faddsubd(a1stg_faddsubd), 
        .a1stg_faddsubs(a1stg_faddsubs), .a1stg_fsdtoix(a1stg_fsdtoix), 
        .a6stg_step(a6stg_step), .a1stg_fstod(a1stg_fstod), .a1stg_fdtos(
        a1stg_fdtos), .a1stg_fstoi(a1stg_fstoi), .a1stg_fstox(a1stg_fstox), 
        .a1stg_fdtoi(a1stg_fdtoi), .a1stg_fdtox(a1stg_fdtox), 
        .a2stg_fsdtoix_fdtos(a2stg_fsdtoix_fdtos), .a2stg_faddsubop(
        a2stg_faddsubop), .a2stg_fitos(a2stg_fitos), .a2stg_fitod(a2stg_fitod), 
        .a2stg_fxtos(a2stg_fxtos), .a2stg_fxtod(a2stg_fxtod), .a3stg_exp_7ff(
        a3stg_exp_7ff), .a3stg_exp_ff(a3stg_exp_ff), .a3stg_exp_add(
        a3stg_exp_add), .a3stg_inc_exp_inv(a3stg_inc_exp_inv), 
        .a3stg_same_exp_inv(a3stg_same_exp_inv), .a3stg_dec_exp_inv(
        a3stg_dec_exp_inv), .a3stg_faddsubop(a3stg_faddsubop), 
        .a3stg_fdtos_inv(a3stg_fdtos_inv), .a4stg_fixtos_fxtod_inv(
        a4stg_fixtos_fxtod_inv), .a4stg_shl_cnt(a4stg_shl_cnt), 
        .a4stg_denorm_inv(a4stg_denorm_inv), .a4stg_rndadd_cout(
        a4stg_rndadd_cout), .add_exp_out_expinc(add_exp_out_expinc), 
        .add_exp_out_exp(add_exp_out_exp), .add_exp_out_exp1(add_exp_out_exp1), 
        .a4stg_in_of(a4stg_in_of), .add_exp_out_expadd(add_exp_out_expadd), 
        .a4stg_dblop(a4stg_dblop), .a4stg_to_0_inv(a4stg_to_0_inv), 
        .fadd_clken_l(fadd_clken_l), .rclk(rclk), .a1stg_expadd3_11(
        a1stg_expadd3_11), .a1stg_expadd1_11_0(a1stg_expadd1_11_0), 
        .a1stg_expadd4_inv(a1stg_expadd4_inv), .a1stg_expadd2_5_0(
        a1stg_expadd2_5_0), .a2stg_exp(a2stg_exp), .a2stg_expadd(a2stg_expadd), 
        .a3stg_exp_10_0(a3stg_exp_10_0), .a4stg_exp_11_0(a4stg_exp_11_0), 
        .add_exp_out(add_exp_out), .se(se_add_exp), .si(net211162) );
  fpu_add_frac_dp fpu_add_frac_dp ( .inq_in1(inq_in1[62:0]), .inq_in2(inq_in2), 
        .a1stg_step(a1stg_stepa), .a1stg_sngop(a1stg_sngop), 
        .a1stg_expadd3_11(a1stg_expadd3_11), .a1stg_norm_dbl_in1(
        a1stg_norm_dbl_in1), .a1stg_denorm_dbl_in1(a1stg_denorm_dbl_in1), 
        .a1stg_norm_sng_in1(a1stg_norm_sng_in1), .a1stg_denorm_sng_in1(
        a1stg_denorm_sng_in1), .a1stg_norm_dbl_in2(a1stg_norm_dbl_in2), 
        .a1stg_denorm_dbl_in2(a1stg_denorm_dbl_in2), .a1stg_norm_sng_in2(
        a1stg_norm_sng_in2), .a1stg_denorm_sng_in2(a1stg_denorm_sng_in2), 
        .a1stg_intlngop(a1stg_intlngop), .a2stg_frac1_in_frac1(
        a2stg_frac1_in_frac1), .a2stg_frac1_in_frac2(a2stg_frac1_in_frac2), 
        .a1stg_2nan_in_inv(a1stg_2nan_in_inv), .a1stg_faddsubop_inv(
        a1stg_faddsubop_inv), .a2stg_frac1_in_qnan(a2stg_frac1_in_qnan), 
        .a2stg_frac1_in_nv(a2stg_frac1_in_nv), .a2stg_frac1_in_nv_dbl(
        a2stg_frac1_in_nv_dbl), .a6stg_step(a6stg_step), 
        .a2stg_frac2_in_frac1(a2stg_frac2_in_frac1), .a2stg_frac2_in_qnan(
        a2stg_frac2_in_qnan), .a2stg_shr_cnt_in(a2stg_shr_cnt_in), 
        .a2stg_shr_cnt_5_inv_in(a2stg_shr_cnt_5_inv_in), 
        .a2stg_shr_frac2_shr_int(a2stg_shr_frac2_shr_int), 
        .a2stg_shr_frac2_shr_dbl(a2stg_shr_frac2_shr_dbl), 
        .a2stg_shr_frac2_shr_sng(a2stg_shr_frac2_shr_sng), 
        .a2stg_shr_frac2_max(a2stg_shr_frac2_max), .a2stg_expadd_11(
        a2stg_expadd[12]), .a2stg_sub_step(a2stg_sub_step), 
        .a2stg_fracadd_frac2_inv_in(a2stg_fracadd_frac2_inv_in), 
        .a2stg_fracadd_frac2_inv_shr1_in(a2stg_fracadd_frac2_inv_shr1_in), 
        .a2stg_fracadd_frac2(a2stg_fracadd_frac2), .a2stg_fracadd_cin_in(
        a2stg_fracadd_cin_in), .a2stg_exp(a2stg_exp[5:0]), 
        .a2stg_expdec_neq_0(a2stg_expdec_neq_0), .a3stg_faddsubopa(
        a3stg_faddsubopa), .a3stg_sub_in(a3stg_sub_in), .a3stg_exp10_0_eq0(
        a3stg_exp10_0_eq0), .a3stg_exp10_1_eq0(a3stg_exp10_1_eq0), 
        .a3stg_exp_0(a3stg_exp_10_0[0]), .a4stg_rnd_frac_add_inv(
        a4stg_rnd_frac_add_inv), .a3stg_fdtos_inv(a3stg_fdtos_inv), 
        .a4stg_fixtos_fxtod_inv(a4stg_fixtos_fxtod_inv), .a4stg_rnd_sng(
        a4stg_rnd_sng), .a4stg_rnd_dbl(a4stg_rnd_dbl), .a4stg_shl_cnt_in(
        a4stg_shl_cnt_in), .add_frac_out_rndadd(add_frac_out_rndadd), 
        .add_frac_out_rnd_frac(add_frac_out_rnd_frac), .a4stg_in_of(
        a4stg_in_of), .add_frac_out_shl(add_frac_out_shl), .a4stg_to_0(
        a4stg_to_0), .fadd_clken_l(fadd_clken_l), .rclk(rclk), 
        .a1stg_in2_neq_in1_frac(a1stg_in2_neq_in1_frac), 
        .a1stg_in2_gt_in1_frac(a1stg_in2_gt_in1_frac), .a1stg_in2_eq_in1_exp(
        a1stg_in2_eq_in1_exp), .a2stg_frac2_63(a2stg_frac2_63), 
        .a2stg_frac2hi_neq_0(a2stg_frac2hi_neq_0), .a2stg_frac2lo_neq_0(
        a2stg_frac2lo_neq_0), .a3stg_fsdtoix_nx(a3stg_fsdtoix_nx), 
        .a3stg_fsdtoi_nx(a3stg_fsdtoi_nx), .a3stg_denorm(a3stg_denorm), 
        .a3stg_lead0(a3stg_lead0), .a4stg_shl_cnt(a4stg_shl_cnt), 
        .a4stg_denorm_inv(a4stg_denorm_inv), .a3stg_inc_exp_inv(
        a3stg_inc_exp_inv), .a3stg_same_exp_inv(a3stg_same_exp_inv), 
        .a3stg_dec_exp_inv(a3stg_dec_exp_inv), .a4stg_rnd_frac_40(
        a4stg_rnd_frac_40), .a4stg_rnd_frac_39(a4stg_rnd_frac_39), 
        .a4stg_rnd_frac_11(a4stg_rnd_frac_11), .a4stg_rnd_frac_10(
        a4stg_rnd_frac_10), .a4stg_rndadd_cout(a4stg_rndadd_cout), 
        .a4stg_frac_9_0_nx(a4stg_frac_9_0_nx), .a4stg_frac_dbl_nx(
        a4stg_frac_dbl_nx), .a4stg_frac_38_0_nx(a4stg_frac_38_0_nx), 
        .a4stg_frac_sng_nx(a4stg_frac_sng_nx), .a4stg_frac_neq_0(
        a4stg_frac_neq_0), .a4stg_shl_data_neq_0(a4stg_shl_data_neq_0), 
        .add_of_out_cout(add_of_out_cout), .add_frac_out(add_frac_out), .se(
        se_add_frac), .si(net211161), .a4stg_round_BAR(a4stg_round) );
endmodule


module dffrl_async_SIZE1_3 ( din, clk, rst_l, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  wire   N4, n1;

  DFFARX1_RVT \q_reg[0]  ( .D(N4), .CLK(clk), .RSTB(rst_l), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
endmodule


module dffe_SIZE1_87 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_86 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_85 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_84 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_83 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_82 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_81 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_80 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_79 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_78 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_77 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_76 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_75 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_74 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_73 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_72 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_71 ( din, en, clk, se, si, so, \q[0]  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0] ;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(\q[0] ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_70 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_69 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n2, n3, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n2) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n3), .A4(din[0]), .A5(n2), .Y(n5)
         );
endmodule


module dffe_SIZE1_68 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_67 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_66 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_65 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_64 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_63 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dff_SIZE8_3 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;

  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
endmodule


module dff_SIZE1_30 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dffe_SIZE1_62 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE4_2 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N4, net24462, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_2 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24462), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24462), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24462), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24462), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24462), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE1_61 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE4_1 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N4, net24462, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE4_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24462), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24462), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24462), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24462), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24462), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE1_60 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE2_9 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_10 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_10 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE5 ( din, rst, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input rst, en, clk, se;
  wire   N11, N12, N13, N14, N15, net24444, n4, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE5 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24444), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N15), .CLK(net24444), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N14), .CLK(net24444), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N13), .CLK(net24444), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N12), .CLK(net24444), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N11), .CLK(net24444), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N11) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N12) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N13) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N14) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N15) );
  NAND2X0_RVT U11 ( .A1(n3), .A2(n2), .Y(n4) );
endmodule


module dffe_SIZE2_8 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_9 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_9 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_5 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_5 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffe_SIZE2_7 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_8 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_8 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_4 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_4 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffe_SIZE2_6 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_7 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_7 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_3 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_3 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffe_SIZE2_5 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_6 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_6 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_2 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_2 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffe_SIZE2_4 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_5 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_5 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE4_1 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N10, N11, N12, N13, net24426, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE4_1 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24426), .TE(1'b0) );
  DFFX1_RVT \q_reg[3]  ( .D(N13), .CLK(net24426), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N12), .CLK(net24426), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N11), .CLK(net24426), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N10), .CLK(net24426), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N11) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N12) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N13) );
  NAND2X0_RVT U10 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffe_SIZE2_3 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_4 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_4 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffre_SIZE1_9 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_3 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_3 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE10_1 ( din, en, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, net24408, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE10_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24408), .TE(1'b0) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24408), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24408), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24408), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24408), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24408), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24408), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24408), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24408), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24408), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24408), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  OR2X1_RVT U14 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffre_SIZE1_8 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffe_SIZE1_59 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_58 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_57 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_56 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_55 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_54 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_53 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_52 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_51 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_50 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_49 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_48 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_47 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_46 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_45 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_44 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_43 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_42 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_41 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_40 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_39 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_38 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_37 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_36 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_35 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_34 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_33 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE6_0 ( din, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, net24390, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE6_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24390), .TE(1'b0) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24390), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24390), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24390), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24390), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24390), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24390), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  OR2X1_RVT U10 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE6_1 ( din, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, net24390, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE6_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24390), .TE(1'b0) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24390), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24390), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24390), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24390), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24390), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24390), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  OR2X1_RVT U10 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE7_0 ( din, en, clk, q, se, si, so );
  input [6:0] din;
  output [6:0] q;
  input [6:0] si;
  output [6:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, net24372, n3, n1;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE7_0 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24372), .TE(1'b0) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24372), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24372), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24372), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24372), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24372), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24372), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24372), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  OR2X1_RVT U11 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE7_1 ( din, en, clk, q, se, si, so );
  input [6:0] din;
  output [6:0] q;
  input [6:0] si;
  output [6:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, net24372, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE7_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24372), .TE(1'b0) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24372), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24372), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24372), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24372), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24372), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24372), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24372), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  OR2X1_RVT U11 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE1_32 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_31 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module fpu_mul_ctl ( inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, inq_op, inq_mul, inq_rnd_mode, inq_id, inq_in1_63, 
        inq_in2_63, mul_dest_rdy, m5stg_exp, m5stg_fracadd_cout, 
        m5stg_frac_neq_0, m5stg_frac_dbl_nx, m5stg_frac_sng_nx, m1stg_ld0_1, 
        m1stg_ld0_2, m3stg_exp, m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv, 
        m3stg_ld0_inv, m4stg_exp, m4stg_frac_105, m5stg_frac, arst_l, grst_l, 
        rclk, mul_pipe_active, m1stg_snan_sng_in1, m1stg_snan_dbl_in1, 
        m1stg_snan_sng_in2, m1stg_snan_dbl_in2, m1stg_step, m1stg_sngop, 
        m1stg_dblop, m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld, m2stg_fmuls, 
        m2stg_fmuld, m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda, 
        m6stg_fmul_in, m6stg_id_in, m6stg_fmul_dbl_dst, m6stg_fmuls, 
        m6stg_step, mul_sign_out, m5stg_in_of, mul_exc_out, 
        m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm, m2stg_frac1_sng_norm, 
        m2stg_frac1_sng_dnrm, m2stg_frac1_inf, m2stg_frac2_dbl_norm, 
        m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, m2stg_frac2_sng_dnrm, 
        m2stg_frac2_inf, m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, 
        m2stg_exp_expadd, m2stg_exp_0bff, m2stg_exp_017f, m2stg_exp_04ff, 
        m2stg_exp_zero, m3bstg_ld0_inv, m4stg_sh_cnt_in, m4stg_inc_exp_54, 
        m4stg_inc_exp_55, m4stg_inc_exp_105, m4stg_left_shift_step, 
        m4stg_right_shift_step, m5stg_to_0, m5stg_to_0_inv, 
        mul_frac_out_fracadd, mul_frac_out_frac, mul_exp_out_exp_plus1, 
        mul_exp_out_exp, mula_rst_l, se, si, so, mul_dest_rdya_BAR );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [12:0] m5stg_exp;
  input [5:0] m1stg_ld0_1;
  input [5:0] m1stg_ld0_2;
  input [12:0] m3stg_exp;
  input [5:0] m3stg_ld0_inv;
  input [12:0] m4stg_exp;
  input [32:0] m5stg_frac;
  output [9:0] m6stg_id_in;
  output [4:0] mul_exc_out;
  output [6:0] m3bstg_ld0_inv;
  output [5:0] m4stg_sh_cnt_in;
  input inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_mul,
         inq_in1_63, inq_in2_63, mul_dest_rdy, m5stg_fracadd_cout,
         m5stg_frac_neq_0, m5stg_frac_dbl_nx, m5stg_frac_sng_nx,
         m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv, m4stg_frac_105, arst_l,
         grst_l, rclk, se, si, mul_dest_rdya_BAR;
  output mul_pipe_active, m1stg_snan_sng_in1, m1stg_snan_dbl_in1,
         m1stg_snan_sng_in2, m1stg_snan_dbl_in2, m1stg_step, m1stg_sngop,
         m1stg_dblop, m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld, m2stg_fmuls,
         m2stg_fmuld, m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda,
         m6stg_fmul_in, m6stg_fmul_dbl_dst, m6stg_fmuls, m6stg_step,
         mul_sign_out, m5stg_in_of, m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm,
         m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, m2stg_frac1_inf,
         m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm,
         m2stg_frac2_sng_dnrm, m2stg_frac2_inf, m1stg_inf_zero_in,
         m1stg_inf_zero_in_dbl, m2stg_exp_expadd, m2stg_exp_0bff,
         m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero, m4stg_inc_exp_54,
         m4stg_inc_exp_55, m4stg_inc_exp_105, m4stg_left_shift_step,
         m4stg_right_shift_step, m5stg_to_0, m5stg_to_0_inv,
         mul_frac_out_fracadd, mul_frac_out_frac, mul_exp_out_exp_plus1,
         mul_exp_out_exp, mula_rst_l, so;
  wire   mul_dest_rdya, mul_exc_out_0, mul_frac_out_fracadd, mul_frac_out_frac,
         mul_frac_in1_51, mul_frac_in1_54, mul_frac_in1_53_0_neq_0,
         mul_frac_in1_50_0_neq_0, mul_frac_in1_53_32_neq_0,
         mul_exp_in1_exp_eq_0, mul_exp_in1_exp_neq_ffs, mul_frac_in2_51,
         mul_frac_in2_54, mul_frac_in2_53_0_neq_0, mul_frac_in2_50_0_neq_0,
         mul_frac_in2_53_32_neq_0, mul_exp_in2_exp_eq_0,
         mul_exp_in2_exp_neq_ffs, m1stg_snan_in1, m1stg_snan_in2,
         m1stg_qnan_in1, m1stg_qnan_in2, m2stg_snan_in1, m2stg_snan_in2,
         m2stg_qnan_in1, m2stg_qnan_in2, m1stg_nan_in2, m2stg_nan_in2,
         m1stg_inf_in1, m1stg_inf_in2, m1stg_inf_in, m2stg_inf_in1,
         m2stg_inf_in2, m2stg_inf_in, m1stg_zero_in1, m1stg_zero_in2,
         m1stg_zero_in, m2stg_zero_in1, m2stg_zero_in2, m2stg_zero_in,
         m1stg_mul, m1stg_mul_in, \m1stg_opdec[3] , \m6stg_opdec[4] ,
         mul_pipe_active_in, m1stg_sign1, m1stg_sign2, m2stg_sign1,
         m2stg_sign2, m2stg_of_mask, m2stg_sign, m3astg_sign, m2stg_nv,
         m3astg_nv, m3astg_of_mask, m3bstg_sign, m3bstg_nv, m3bstg_of_mask,
         m3stg_sign, m3stg_nv, m3stg_of_mask, m4stg_sign, m4stg_nv,
         m4stg_of_mask, m5stg_sign, m5stg_nv, m5stg_of_mask,
         mul_of_out_tmp1_in, mul_of_out_tmp1, mul_of_out_tmp2, mul_of_out_cout,
         mul_uf_out_in, mul_nx_out_in, mul_nx_out, m4stg_expadd_eq_0,
         m4stg_right_shift_in, m4stg_right_shift, \m3stg_exp_inv_plus2[1] ,
         n153, n154, n155, n157, n160, n161, n162, n163, n164, n165, n166,
         n168, \intadd_4/CI , \intadd_4/SUM[4] , \intadd_4/SUM[3] ,
         \intadd_4/SUM[2] , \intadd_4/SUM[1] , \intadd_4/SUM[0] ,
         \intadd_4/n5 , \intadd_4/n4 , \intadd_4/n3 , \intadd_4/n2 ,
         \intadd_4/n1 , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n156,
         n158, n159, n167, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n200;
  wire   [3:0] m1stg_sngopa;
  wire   [3:0] m1stg_dblopa;
  wire   [7:0] m1stg_op;
  wire   [7:0] m1stg_op_in;
  wire   [1:0] m1stg_rnd_mode;
  wire   [4:0] m1stg_id;
  wire   [4:3] m2stg_opdec;
  wire   [1:0] m2stg_rnd_mode;
  wire   [4:0] m2stg_id;
  wire   [4:1] m3astg_opdec;
  wire   [1:0] m3astg_rnd_mode;
  wire   [4:0] m3astg_id;
  wire   [4:1] m3bstg_opdec;
  wire   [1:0] m3bstg_rnd_mode;
  wire   [4:0] m3bstg_id;
  wire   [4:1] m3stg_opdec;
  wire   [1:0] m3stg_rnd_mode;
  wire   [4:0] m3stg_id;
  wire   [4:1] m4stg_opdec;
  wire   [1:0] m4stg_rnd_mode;
  wire   [4:0] m4stg_id;
  wire   [4:3] m5stg_opdec;
  wire   [1:0] m5stg_rnd_mode;
  wire   [4:0] m5stg_id;
  wire   [9:0] m6stg_id;
  wire   [5:0] m2stg_ld0_1_in;
  wire   [5:0] m2stg_ld0_1;
  wire   [5:0] m2stg_ld0_2_in;
  wire   [5:0] m2stg_ld0_2;
  wire   [6:0] m3astg_ld0_inv;
  assign mul_dest_rdya = mul_dest_rdya_BAR;
  assign mul_exc_out[0] = mul_exc_out_0;
  assign mul_exp_out_exp_plus1 = mul_frac_out_fracadd;
  assign mul_exp_out_exp = mul_frac_out_frac;
  assign \m3stg_exp_inv_plus2[1]  = m3stg_exp[1];
  assign so = 1'b0;
  assign mul_exc_out[1] = 1'b0;

  dffrl_async_SIZE1_3 dffrl_mul_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(mula_rst_l), .se(se), .si(1'b0) );
  dffe_SIZE1_87 i_mul_frac_in1_51 ( .din(inq_in1_51), .en(n200), .clk(rclk), 
        .q(mul_frac_in1_51), .se(se), .si(1'b0) );
  dffe_SIZE1_86 i_mul_frac_in1_54 ( .din(inq_in1_54), .en(n200), .clk(rclk), 
        .q(mul_frac_in1_54), .se(se), .si(1'b0) );
  dffe_SIZE1_85 i_mul_frac_in1_53_0_neq_0 ( .din(inq_in1_53_0_neq_0), .en(n200), .clk(rclk), .q(mul_frac_in1_53_0_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_84 i_mul_frac_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(n200), .clk(rclk), .q(mul_frac_in1_50_0_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_83 i_mul_frac_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        n200), .clk(rclk), .q(mul_frac_in1_53_32_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_82 i_mul_exp_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(n200), 
        .clk(rclk), .q(mul_exp_in1_exp_eq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_81 i_mul_exp_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        n200), .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (
        mul_exp_in1_exp_neq_ffs) );
  dffe_SIZE1_80 i_mul_frac_in2_51 ( .din(inq_in2_51), .en(n200), .clk(rclk), 
        .q(mul_frac_in2_51), .se(se), .si(1'b0) );
  dffe_SIZE1_79 i_mul_frac_in2_54 ( .din(inq_in2_54), .en(n200), .clk(rclk), 
        .q(mul_frac_in2_54), .se(se), .si(1'b0) );
  dffe_SIZE1_78 i_mul_frac_in2_53_0_neq_0 ( .din(inq_in2_53_0_neq_0), .en(n200), .clk(rclk), .q(mul_frac_in2_53_0_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_77 i_mul_frac_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(n200), .clk(rclk), .q(mul_frac_in2_50_0_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_76 i_mul_frac_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        n200), .clk(rclk), .q(mul_frac_in2_53_32_neq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_75 i_mul_exp_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(n200), 
        .clk(rclk), .q(mul_exp_in2_exp_eq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_74 i_mul_exp_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        n200), .clk(rclk), .q(mul_exp_in2_exp_neq_ffs), .se(se), .si(1'b0) );
  dffe_SIZE1_73 i_m2stg_snan_in1 ( .din(m1stg_snan_in1), .en(n200), .clk(rclk), 
        .se(se), .si(1'b0), .\q[0]_BAR (m2stg_snan_in1) );
  dffe_SIZE1_72 i_m2stg_snan_in2 ( .din(m1stg_snan_in2), .en(n200), .clk(rclk), 
        .q(m2stg_snan_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_71 i_m2stg_qnan_in1 ( .din(m1stg_qnan_in1), .en(n200), .clk(rclk), 
        .se(se), .si(1'b0), .\q[0] (m2stg_qnan_in1) );
  dffe_SIZE1_70 i_m2stg_qnan_in2 ( .din(m1stg_qnan_in2), .en(n200), .clk(rclk), 
        .q(m2stg_qnan_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_69 i_m2stg_nan_in2 ( .din(m1stg_nan_in2), .en(n200), .clk(rclk), 
        .se(se), .si(1'b0), .\q[0]_BAR (m2stg_nan_in2) );
  dffe_SIZE1_68 i_m2stg_inf_in1 ( .din(m1stg_inf_in1), .en(n200), .clk(rclk), 
        .q(m2stg_inf_in1), .se(se), .si(1'b0) );
  dffe_SIZE1_67 i_m2stg_inf_in2 ( .din(m1stg_inf_in2), .en(n200), .clk(rclk), 
        .q(m2stg_inf_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_66 i_m2stg_inf_in ( .din(m1stg_inf_in), .en(n200), .clk(rclk), 
        .q(m2stg_inf_in), .se(se), .si(1'b0) );
  dffe_SIZE1_65 i_m2stg_zero_in1 ( .din(m1stg_zero_in1), .en(n200), .clk(rclk), 
        .q(m2stg_zero_in1), .se(se), .si(1'b0) );
  dffe_SIZE1_64 i_m2stg_zero_in2 ( .din(m1stg_zero_in2), .en(n200), .clk(rclk), 
        .q(m2stg_zero_in2), .se(se), .si(1'b0) );
  dffe_SIZE1_63 i_m2stg_zero_in ( .din(m1stg_zero_in), .en(n200), .clk(rclk), 
        .q(m2stg_zero_in), .se(se), .si(1'b0) );
  dff_SIZE8_3 i_m1stg_op ( .din(m1stg_op_in), .clk(rclk), .q(m1stg_op), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE1_30 i_m1stg_mul ( .din(m1stg_mul_in), .clk(rclk), .q(m1stg_mul), 
        .se(se), .si(1'b0) );
  dffe_SIZE1_62 i_m1stg_sngop ( .din(inq_op[0]), .en(n200), .clk(rclk), .q(
        m1stg_sngop), .se(se), .si(1'b0) );
  dffe_SIZE4_2 i_m1stg_sngopa ( .din({1'b0, 1'b0, 1'b0, inq_op[0]}), .en(n200), 
        .clk(rclk), .q(m1stg_sngopa), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0})
         );
  dffe_SIZE1_61 i_m1stg_dblop ( .din(inq_op[1]), .en(n200), .clk(rclk), .q(
        m1stg_dblop), .se(se), .si(1'b0) );
  dffe_SIZE4_1 i_m1stg_dblopa ( .din({1'b0, 1'b0, 1'b0, inq_op[1]}), .en(n200), 
        .clk(rclk), .q(m1stg_dblopa), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0})
         );
  dffe_SIZE1_60 i_m1stg_dblop_inv ( .din(n168), .en(n200), .clk(rclk), .q(
        m1stg_dblop_inv), .se(se), .si(1'b0) );
  dffe_SIZE2_9 i_m1stg_rnd_mode ( .din(inq_rnd_mode), .en(n200), .clk(rclk), 
        .q(m1stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_10 i_m1stg_id ( .din(inq_id), .en(n200), .clk(rclk), .q(m1stg_id), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE5 i_m2stg_opdec ( .din({m1stg_fmul, \m1stg_opdec[3] , n155, n157, 
        m1stg_fsmuld}), .rst(n153), .en(n200), .clk(rclk), .q({m2stg_opdec, 
        m2stg_fmuls, m2stg_fmuld, m2stg_fsmuld}), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_8 i_m2stg_rnd_mode ( .din(m1stg_rnd_mode), .en(n200), .clk(rclk), 
        .q(m2stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_9 i_m2stg_id ( .din(m1stg_id), .en(n200), .clk(rclk), .q(m2stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_5 i_m3astg_opdec ( .din({m2stg_opdec, m2stg_fmuls, m2stg_fmuld}), 
        .rst(n153), .en(n200), .clk(rclk), .q(m3astg_opdec), .se(se), .si({
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_7 i_m3astg_rnd_mode ( .din(m2stg_rnd_mode), .en(n200), .clk(rclk), 
        .q(m3astg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_8 i_m3astg_id ( .din(m2stg_id), .en(n200), .clk(rclk), .q(
        m3astg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_4 i_m3bstg_opdec ( .din(m3astg_opdec), .rst(n153), .en(n200), 
        .clk(rclk), .q(m3bstg_opdec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0})
         );
  dffe_SIZE2_6 i_m3bstg_rnd_mode ( .din(m3astg_rnd_mode), .en(n200), .clk(rclk), .q(m3bstg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_7 i_m3bstg_id ( .din(m3astg_id), .en(n200), .clk(rclk), .q(
        m3bstg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_3 i_m3stg_opdec ( .din(m3bstg_opdec), .rst(n153), .en(n200), 
        .clk(rclk), .q(m3stg_opdec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_5 i_m3stg_rnd_mode ( .din(m3bstg_rnd_mode), .en(n200), .clk(rclk), 
        .q(m3stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_6 i_m3stg_id ( .din(m3bstg_id), .en(n200), .clk(rclk), .q(
        m3stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_2 i_m4stg_opdec ( .din(m3stg_opdec), .rst(n153), .en(n200), 
        .clk(rclk), .q(m4stg_opdec), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_4 i_m4stg_rnd_mode ( .din(m3stg_rnd_mode), .en(n200), .clk(rclk), 
        .q(m4stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_5 i_m4stg_id ( .din(m3stg_id), .en(n200), .clk(rclk), .q(m4stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE4_1 i_m5stg_opdec ( .din(m4stg_opdec), .rst(n153), .en(n200), 
        .clk(rclk), .q({m5stg_opdec, m5stg_fmuls, m5stg_fmuld}), .se(se), .si(
        {1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE2_3 i_m5stg_rnd_mode ( .din(m4stg_rnd_mode), .en(n200), .clk(rclk), 
        .q(m5stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_4 i_m5stg_id ( .din(m4stg_id), .en(n200), .clk(rclk), .q(m5stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_9 i_m5stg_fmulda ( .din(m4stg_opdec[1]), .rst(n153), .en(n200), 
        .clk(rclk), .q(m5stg_fmulda), .se(se), .si(1'b0) );
  dffre_SIZE3_3 i_m6stg_opdec ( .din({m5stg_opdec, m5stg_fmuls}), .rst(n153), 
        .en(n200), .clk(rclk), .q({\m6stg_opdec[4] , m6stg_fmul_dbl_dst, 
        m6stg_fmuls}), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dffe_SIZE10_1 i_m6stg_id ( .din(m6stg_id_in), .en(n200), .clk(rclk), .q(
        m6stg_id), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_8 i_mul_pipe_active ( .din(mul_pipe_active_in), .rst(n153), .en(
        1'b1), .clk(rclk), .q(mul_pipe_active), .se(se), .si(1'b0) );
  dffe_SIZE1_59 i_m1stg_sign1 ( .din(inq_in1_63), .en(n200), .clk(rclk), .q(
        m1stg_sign1), .se(se), .si(1'b0) );
  dffe_SIZE1_58 i_m1stg_sign2 ( .din(inq_in2_63), .en(n200), .clk(rclk), .q(
        m1stg_sign2), .se(se), .si(1'b0) );
  dffe_SIZE1_57 i_m2stg_sign1 ( .din(m1stg_sign1), .en(n200), .clk(rclk), .q(
        m2stg_sign1), .se(se), .si(1'b0) );
  dffe_SIZE1_56 i_m2stg_sign2 ( .din(m1stg_sign2), .en(n200), .clk(rclk), .q(
        m2stg_sign2), .se(se), .si(1'b0) );
  dffe_SIZE1_55 i_m2stg_of_mask ( .din(n154), .en(n200), .clk(rclk), .q(
        m2stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_54 i_m3astg_sign ( .din(m2stg_sign), .en(n200), .clk(rclk), .q(
        m3astg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_53 i_m3astg_nv ( .din(m2stg_nv), .en(n200), .clk(rclk), .q(
        m3astg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_52 i_m3astg_of_mask ( .din(m2stg_of_mask), .en(n200), .clk(rclk), 
        .q(m3astg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_51 i_m3bstg_sign ( .din(m3astg_sign), .en(n200), .clk(rclk), .q(
        m3bstg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_50 i_m3bstg_nv ( .din(m3astg_nv), .en(n200), .clk(rclk), .q(
        m3bstg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_49 i_m3bstg_of_mask ( .din(m3astg_of_mask), .en(n200), .clk(rclk), 
        .q(m3bstg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_48 i_m3stg_sign ( .din(m3bstg_sign), .en(n200), .clk(rclk), .q(
        m3stg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_47 i_m3stg_nv ( .din(m3bstg_nv), .en(n200), .clk(rclk), .q(
        m3stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_46 i_m3stg_of_mask ( .din(m3bstg_of_mask), .en(n200), .clk(rclk), 
        .q(m3stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_45 i_m4stg_sign ( .din(m3stg_sign), .en(n200), .clk(rclk), .q(
        m4stg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_44 i_m4stg_nv ( .din(m3stg_nv), .en(n200), .clk(rclk), .q(
        m4stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_43 i_m4stg_of_mask ( .din(m3stg_of_mask), .en(n200), .clk(rclk), 
        .q(m4stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_42 i_m5stg_sign ( .din(m4stg_sign), .en(n200), .clk(rclk), .q(
        m5stg_sign), .se(se), .si(1'b0) );
  dffe_SIZE1_41 i_m5stg_nv ( .din(m4stg_nv), .en(n200), .clk(rclk), .q(
        m5stg_nv), .se(se), .si(1'b0) );
  dffe_SIZE1_40 i_m5stg_of_mask ( .din(m4stg_of_mask), .en(n200), .clk(rclk), 
        .q(m5stg_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_39 i_mul_sign_out ( .din(m5stg_sign), .en(n200), .clk(rclk), .q(
        mul_sign_out), .se(se), .si(1'b0) );
  dffe_SIZE1_38 i_mul_nv_out ( .din(m5stg_nv), .en(n200), .clk(rclk), .q(
        mul_exc_out[4]), .se(se), .si(1'b0) );
  dffe_SIZE1_37 i_mul_of_out_tmp1 ( .din(mul_of_out_tmp1_in), .en(n200), .clk(
        rclk), .q(mul_of_out_tmp1), .se(se), .si(1'b0) );
  dffe_SIZE1_36 i_mul_of_out_tmp2 ( .din(m5stg_in_of), .en(n200), .clk(rclk), 
        .q(mul_of_out_tmp2), .se(se), .si(1'b0) );
  dffe_SIZE1_35 i_mul_of_out_cout ( .din(m5stg_fracadd_cout), .en(n200), .clk(
        rclk), .q(mul_of_out_cout), .se(se), .si(1'b0) );
  dffe_SIZE1_34 i_mul_uf_out ( .din(mul_uf_out_in), .en(n200), .clk(rclk), .q(
        mul_exc_out[2]), .se(se), .si(1'b0) );
  dffe_SIZE1_33 i_mul_nx_out ( .din(mul_nx_out_in), .en(n200), .clk(rclk), .q(
        mul_nx_out), .se(se), .si(1'b0) );
  dffe_SIZE6_0 i_m2stg_ld0_1 ( .din(m2stg_ld0_1_in), .en(n200), .clk(rclk), 
        .q(m2stg_ld0_1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE6_1 i_m2stg_ld0_2 ( .din(m2stg_ld0_2_in), .en(n200), .clk(rclk), 
        .q(m2stg_ld0_2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE7_0 i_m3astg_ld0_inv ( .din({n160, n161, n162, n163, n164, n165, 
        n166}), .en(n200), .clk(rclk), .q(m3astg_ld0_inv), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE7_1 i_m3bstg_ld0_inv ( .din(m3astg_ld0_inv), .en(n200), .clk(rclk), 
        .q(m3bstg_ld0_inv), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE1_32 i_m4stg_expadd_eq_0 ( .din(m3stg_expadd_eq_0), .en(n200), 
        .clk(rclk), .q(m4stg_expadd_eq_0), .se(se), .si(1'b0) );
  dffe_SIZE1_31 i_m4stg_right_shift ( .din(m4stg_right_shift_in), .en(n200), 
        .clk(rclk), .q(m4stg_right_shift), .se(se), .si(1'b0) );
  FADDX1_RVT \intadd_4/U6  ( .A(m2stg_ld0_2[1]), .B(m2stg_ld0_1[1]), .CI(
        \intadd_4/CI ), .CO(\intadd_4/n5 ), .S(\intadd_4/SUM[0] ) );
  FADDX1_RVT \intadd_4/U5  ( .A(m2stg_ld0_2[2]), .B(m2stg_ld0_1[2]), .CI(
        \intadd_4/n5 ), .CO(\intadd_4/n4 ), .S(\intadd_4/SUM[1] ) );
  FADDX1_RVT \intadd_4/U4  ( .A(m2stg_ld0_2[3]), .B(m2stg_ld0_1[3]), .CI(
        \intadd_4/n4 ), .CO(\intadd_4/n3 ), .S(\intadd_4/SUM[2] ) );
  FADDX1_RVT \intadd_4/U3  ( .A(m2stg_ld0_2[4]), .B(m2stg_ld0_1[4]), .CI(
        \intadd_4/n3 ), .CO(\intadd_4/n2 ), .S(\intadd_4/SUM[3] ) );
  FADDX1_RVT \intadd_4/U2  ( .A(m2stg_ld0_2[5]), .B(m2stg_ld0_1[5]), .CI(
        \intadd_4/n2 ), .CO(\intadd_4/n1 ), .S(\intadd_4/SUM[4] ) );
  OR3X1_RVT U3 ( .A1(\m3stg_exp_inv_plus2[1] ), .A2(n185), .A3(m3stg_exp[0]), 
        .Y(n186) );
  INVX0_RVT U4 ( .A(inq_op[1]), .Y(n168) );
  INVX0_RVT U5 ( .A(m5stg_in_of), .Y(n34) );
  INVX0_RVT U6 ( .A(n16), .Y(n17) );
  INVX0_RVT U7 ( .A(n180), .Y(n177) );
  INVX0_RVT U8 ( .A(n126), .Y(n88) );
  INVX0_RVT U9 ( .A(n21), .Y(n11) );
  INVX0_RVT U10 ( .A(m5stg_frac[32]), .Y(n18) );
  INVX0_RVT U11 ( .A(m3stg_exp[0]), .Y(n182) );
  OR3X1_RVT U12 ( .A1(m5stg_frac[3]), .A2(m5stg_frac[0]), .A3(m5stg_frac[1]), 
        .Y(n21) );
  INVX0_RVT U13 ( .A(m1stg_snan_in1), .Y(n86) );
  INVX0_RVT U14 ( .A(n69), .Y(n60) );
  INVX0_RVT U15 ( .A(n70), .Y(n44) );
  INVX0_RVT U16 ( .A(n122), .Y(n51) );
  INVX0_RVT U17 ( .A(n76), .Y(m1stg_snan_sng_in2) );
  INVX0_RVT U18 ( .A(n77), .Y(m1stg_snan_dbl_in2) );
  INVX0_RVT U19 ( .A(n121), .Y(n39) );
  INVX0_RVT U20 ( .A(m1stg_dblopa[0]), .Y(n128) );
  INVX0_RVT U21 ( .A(m1stg_sngopa[0]), .Y(n127) );
  INVX0_RVT U22 ( .A(m5stg_fmuls), .Y(n29) );
  INVX0_RVT U23 ( .A(m1stg_dblopa[2]), .Y(n82) );
  INVX0_RVT U24 ( .A(m1stg_sngopa[2]), .Y(n80) );
  INVX0_RVT U25 ( .A(m1stg_op[1]), .Y(n57) );
  INVX0_RVT U26 ( .A(mul_exp_in1_exp_neq_ffs), .Y(n35) );
  INVX0_RVT U27 ( .A(m2stg_snan_in2), .Y(n113) );
  INVX0_RVT U28 ( .A(m1stg_op[0]), .Y(n56) );
  INVX0_RVT U29 ( .A(mul_frac_in2_51), .Y(n37) );
  INVX0_RVT U30 ( .A(mul_frac_in1_54), .Y(n48) );
  INVX0_RVT U31 ( .A(mul_frac_in1_51), .Y(n36) );
  INVX0_RVT U32 ( .A(mul_frac_in2_54), .Y(n49) );
  INVX0_RVT U33 ( .A(m5stg_rnd_mode[1]), .Y(n24) );
  OAI22X1_RVT U34 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .Y(n1) );
  NAND2X0_RVT U35 ( .A1(mul_dest_rdya), .A2(\m6stg_opdec[4] ), .Y(m6stg_step)
         );
  INVX1_RVT U36 ( .A(m6stg_step), .Y(n103) );
  INVX1_RVT U37 ( .A(n103), .Y(n200) );
  NAND2X0_RVT U38 ( .A1(m5stg_sign), .A2(m5stg_rnd_mode[1]), .Y(n3) );
  HADDX1_RVT U39 ( .A0(m5stg_rnd_mode[0]), .B0(n3), .SO(m5stg_to_0_inv) );
  NOR4X1_RVT U40 ( .A1(m5stg_frac[2]), .A2(m5stg_frac[30]), .A3(m5stg_frac[28]), .A4(m5stg_frac[21]), .Y(n7) );
  NOR4X1_RVT U41 ( .A1(m5stg_frac[11]), .A2(m5stg_frac[8]), .A3(m5stg_frac[10]), .A4(m5stg_frac[9]), .Y(n6) );
  NOR4X1_RVT U42 ( .A1(m5stg_frac[24]), .A2(m5stg_frac[25]), .A3(
        m5stg_frac[26]), .A4(m5stg_frac[27]), .Y(n5) );
  NOR4X1_RVT U43 ( .A1(m5stg_frac[29]), .A2(m5stg_frac[20]), .A3(
        m5stg_frac[22]), .A4(m5stg_frac[23]), .Y(n4) );
  NAND4X0_RVT U44 ( .A1(n7), .A2(n6), .A3(n5), .A4(n4), .Y(n13) );
  NOR4X1_RVT U45 ( .A1(m5stg_frac[14]), .A2(m5stg_frac[15]), .A3(
        m5stg_frac[12]), .A4(m5stg_frac[13]), .Y(n10) );
  NOR4X1_RVT U46 ( .A1(m5stg_frac[4]), .A2(m5stg_frac[5]), .A3(m5stg_frac[6]), 
        .A4(m5stg_frac[7]), .Y(n9) );
  NOR4X1_RVT U47 ( .A1(m5stg_frac[17]), .A2(m5stg_frac[18]), .A3(
        m5stg_frac[16]), .A4(m5stg_frac[19]), .Y(n8) );
  NAND4X0_RVT U48 ( .A1(n11), .A2(n10), .A3(n9), .A4(n8), .Y(n12) );
  OR2X1_RVT U49 ( .A1(n13), .A2(n12), .Y(n16) );
  AO222X1_RVT U50 ( .A1(m5stg_fmuld), .A2(m5stg_frac[1]), .A3(m5stg_fmuld), 
        .A4(m5stg_frac[0]), .A5(m5stg_fmuld), .A6(m5stg_frac[2]), .Y(n14) );
  AO221X1_RVT U51 ( .A1(m5stg_fmuls), .A2(m5stg_frac[31]), .A3(m5stg_fmuls), 
        .A4(n16), .A5(n14), .Y(n15) );
  AND2X1_RVT U52 ( .A1(m5stg_to_0_inv), .A2(n15), .Y(n26) );
  AND2X1_RVT U53 ( .A1(m5stg_frac[31]), .A2(m5stg_fmuls), .Y(n20) );
  NAND2X0_RVT U54 ( .A1(n18), .A2(n17), .Y(n19) );
  AND2X1_RVT U55 ( .A1(n20), .A2(n19), .Y(n22) );
  OAI222X1_RVT U56 ( .A1(n22), .A2(m5stg_fmuld), .A3(n22), .A4(m5stg_frac[2]), 
        .A5(n22), .A6(n21), .Y(n23) );
  NAND2X0_RVT U57 ( .A1(n24), .A2(n23), .Y(n25) );
  AND2X1_RVT U58 ( .A1(n26), .A2(n25), .Y(n191) );
  AND4X1_RVT U59 ( .A1(m5stg_exp[7]), .A2(m5stg_exp[3]), .A3(m5stg_exp[6]), 
        .A4(m5stg_exp[4]), .Y(n27) );
  AND4X1_RVT U60 ( .A1(m5stg_exp[5]), .A2(m5stg_exp[1]), .A3(m5stg_exp[2]), 
        .A4(n27), .Y(n31) );
  NAND4X0_RVT U61 ( .A1(m5stg_exp[9]), .A2(m5stg_exp[10]), .A3(m5stg_fmuld), 
        .A4(m5stg_exp[8]), .Y(n28) );
  NAND2X0_RVT U62 ( .A1(n29), .A2(n28), .Y(n30) );
  AND2X1_RVT U63 ( .A1(n31), .A2(n30), .Y(n116) );
  AO22X1_RVT U64 ( .A1(m5stg_fmuld), .A2(m5stg_exp[11]), .A3(n116), .A4(
        m5stg_exp[0]), .Y(n33) );
  OR4X1_RVT U65 ( .A1(m5stg_exp[9]), .A2(m5stg_exp[10]), .A3(m5stg_exp[8]), 
        .A4(m5stg_exp[11]), .Y(n118) );
  INVX1_RVT U66 ( .A(m5stg_exp[12]), .Y(n115) );
  AND2X1_RVT U67 ( .A1(m5stg_of_mask), .A2(n115), .Y(n32) );
  OA221X1_RVT U68 ( .A1(n33), .A2(m5stg_fmuls), .A3(n33), .A4(n118), .A5(n32), 
        .Y(m5stg_in_of) );
  AND2X1_RVT U69 ( .A1(n191), .A2(n34), .Y(mul_frac_out_fracadd) );
  NAND2X0_RVT U70 ( .A1(mul_exp_in2_exp_neq_ffs), .A2(n35), .Y(n47) );
  NAND2X0_RVT U71 ( .A1(m1stg_dblopa[3]), .A2(n47), .Y(n70) );
  AND3X1_RVT U72 ( .A1(m1stg_dblopa[0]), .A2(mul_exp_in1_exp_eq_0), .A3(n70), 
        .Y(m2stg_frac1_dbl_dnrm) );
  INVX1_RVT U73 ( .A(mul_exp_in1_exp_eq_0), .Y(n66) );
  AND2X1_RVT U74 ( .A1(n66), .A2(m1stg_dblopa[0]), .Y(n42) );
  NAND3X0_RVT U75 ( .A1(mul_exp_in1_exp_neq_ffs), .A2(mul_frac_in1_51), .A3(
        m1stg_dblopa[1]), .Y(n121) );
  OA21X1_RVT U76 ( .A1(mul_frac_in2_51), .A2(mul_frac_in2_50_0_neq_0), .A3(
        m1stg_dblopa[2]), .Y(n75) );
  INVX1_RVT U77 ( .A(mul_exp_in2_exp_neq_ffs), .Y(n73) );
  NAND2X0_RVT U78 ( .A1(n75), .A2(n73), .Y(n38) );
  AND4X1_RVT U79 ( .A1(mul_frac_in1_50_0_neq_0), .A2(mul_exp_in1_exp_neq_ffs), 
        .A3(m1stg_dblopa[1]), .A4(n36), .Y(m1stg_snan_dbl_in1) );
  NAND4X0_RVT U80 ( .A1(mul_frac_in2_50_0_neq_0), .A2(m1stg_dblopa[1]), .A3(
        n73), .A4(n37), .Y(n77) );
  AOI22X1_RVT U81 ( .A1(n39), .A2(n38), .A3(m1stg_snan_dbl_in1), .A4(n77), .Y(
        n40) );
  NAND2X0_RVT U82 ( .A1(n44), .A2(n40), .Y(n41) );
  AND2X1_RVT U83 ( .A1(n42), .A2(n41), .Y(m2stg_frac1_dbl_norm) );
  INVX1_RVT U84 ( .A(mul_exp_in2_exp_eq_0), .Y(n68) );
  AND2X1_RVT U85 ( .A1(n68), .A2(m1stg_dblopa[0]), .Y(n46) );
  NAND3X0_RVT U86 ( .A1(mul_frac_in2_51), .A2(m1stg_dblopa[1]), .A3(n73), .Y(
        n78) );
  OA21X1_RVT U87 ( .A1(m1stg_snan_dbl_in1), .A2(n78), .A3(n77), .Y(n43) );
  NAND2X0_RVT U88 ( .A1(n44), .A2(n43), .Y(n45) );
  AND2X1_RVT U89 ( .A1(n46), .A2(n45), .Y(m2stg_frac2_dbl_norm) );
  AND3X1_RVT U90 ( .A1(m1stg_dblopa[0]), .A2(mul_exp_in2_exp_eq_0), .A3(n70), 
        .Y(m2stg_frac2_dbl_dnrm) );
  AND2X1_RVT U91 ( .A1(n66), .A2(m1stg_sngopa[0]), .Y(n54) );
  NAND2X0_RVT U92 ( .A1(m1stg_sngopa[3]), .A2(n47), .Y(n69) );
  NAND3X0_RVT U93 ( .A1(mul_exp_in1_exp_neq_ffs), .A2(mul_frac_in1_54), .A3(
        m1stg_sngopa[1]), .Y(n122) );
  OA21X1_RVT U94 ( .A1(mul_frac_in2_54), .A2(mul_frac_in2_53_32_neq_0), .A3(
        m1stg_sngopa[2]), .Y(n74) );
  NAND2X0_RVT U95 ( .A1(n74), .A2(n73), .Y(n50) );
  AND4X1_RVT U96 ( .A1(mul_exp_in1_exp_neq_ffs), .A2(mul_frac_in1_53_32_neq_0), 
        .A3(m1stg_sngopa[1]), .A4(n48), .Y(m1stg_snan_sng_in1) );
  NAND4X0_RVT U97 ( .A1(mul_frac_in2_53_32_neq_0), .A2(m1stg_sngopa[1]), .A3(
        n73), .A4(n49), .Y(n76) );
  AOI22X1_RVT U98 ( .A1(n51), .A2(n50), .A3(m1stg_snan_sng_in1), .A4(n76), .Y(
        n52) );
  NAND2X0_RVT U99 ( .A1(n60), .A2(n52), .Y(n53) );
  AND2X1_RVT U100 ( .A1(n54), .A2(n53), .Y(m2stg_frac1_sng_norm) );
  AND3X1_RVT U101 ( .A1(m1stg_sngopa[0]), .A2(mul_exp_in1_exp_eq_0), .A3(n69), 
        .Y(m2stg_frac1_sng_dnrm) );
  AND3X1_RVT U102 ( .A1(m1stg_sngopa[0]), .A2(mul_exp_in2_exp_eq_0), .A3(n69), 
        .Y(m2stg_frac2_sng_dnrm) );
  NAND2X0_RVT U103 ( .A1(m1stg_op[6]), .A2(m1stg_op[3]), .Y(n55) );
  NOR4X1_RVT U104 ( .A1(m1stg_op[4]), .A2(m1stg_op[7]), .A3(m1stg_op[2]), .A4(
        n55), .Y(n58) );
  INVX1_RVT U105 ( .A(m1stg_op[5]), .Y(n134) );
  AND4X1_RVT U106 ( .A1(m1stg_op[1]), .A2(n58), .A3(n56), .A4(n134), .Y(n157)
         );
  AND3X1_RVT U107 ( .A1(n58), .A2(m1stg_op[0]), .A3(n57), .Y(n135) );
  OR2X1_RVT U108 ( .A1(n135), .A2(n157), .Y(m1stg_fmul) );
  NOR2X0_RVT U109 ( .A1(n103), .A2(m1stg_mul), .Y(m1stg_step) );
  AND2X1_RVT U110 ( .A1(n68), .A2(m1stg_sngopa[0]), .Y(n62) );
  NAND3X0_RVT U111 ( .A1(mul_frac_in2_54), .A2(m1stg_sngopa[1]), .A3(n73), .Y(
        n79) );
  OA21X1_RVT U112 ( .A1(m1stg_snan_sng_in1), .A2(n79), .A3(n76), .Y(n59) );
  NAND2X0_RVT U113 ( .A1(n60), .A2(n59), .Y(n61) );
  AND2X1_RVT U114 ( .A1(n62), .A2(n61), .Y(m2stg_frac2_sng_norm) );
  NOR2X0_RVT U115 ( .A1(mul_frac_in2_51), .A2(mul_frac_in2_50_0_neq_0), .Y(n64) );
  NOR2X0_RVT U116 ( .A1(mul_frac_in2_54), .A2(mul_frac_in2_53_32_neq_0), .Y(
        n63) );
  AO22X1_RVT U117 ( .A1(n64), .A2(m1stg_dblopa[2]), .A3(n63), .A4(
        m1stg_sngopa[2]), .Y(n65) );
  AND2X1_RVT U118 ( .A1(n73), .A2(n65), .Y(m1stg_inf_in2) );
  NOR3X0_RVT U119 ( .A1(mul_frac_in1_54), .A2(mul_frac_in1_53_0_neq_0), .A3(
        n66), .Y(m1stg_zero_in1) );
  NOR2X0_RVT U120 ( .A1(mul_frac_in1_50_0_neq_0), .A2(mul_frac_in1_51), .Y(n83) );
  NOR2X0_RVT U121 ( .A1(mul_frac_in1_54), .A2(mul_frac_in1_53_32_neq_0), .Y(
        n81) );
  AO22X1_RVT U122 ( .A1(m1stg_dblopa[2]), .A2(n83), .A3(m1stg_sngopa[2]), .A4(
        n81), .Y(n67) );
  AND2X1_RVT U123 ( .A1(mul_exp_in1_exp_neq_ffs), .A2(n67), .Y(m1stg_inf_in1)
         );
  NOR3X0_RVT U124 ( .A1(mul_frac_in2_54), .A2(mul_frac_in2_53_0_neq_0), .A3(
        n68), .Y(m1stg_zero_in2) );
  AO22X1_RVT U125 ( .A1(m1stg_inf_in2), .A2(m1stg_zero_in1), .A3(m1stg_inf_in1), .A4(m1stg_zero_in2), .Y(m1stg_inf_zero_in) );
  INVX1_RVT U126 ( .A(mula_rst_l), .Y(n153) );
  OR2X1_RVT U127 ( .A1(m1stg_zero_in1), .A2(m1stg_zero_in2), .Y(m1stg_zero_in)
         );
  NAND2X0_RVT U128 ( .A1(n70), .A2(n69), .Y(n136) );
  NOR2X0_RVT U129 ( .A1(n136), .A2(m1stg_zero_in), .Y(m2stg_exp_expadd) );
  INVX1_RVT U130 ( .A(n136), .Y(n154) );
  INVX1_RVT U131 ( .A(m4stg_right_shift), .Y(m4stg_inc_exp_55) );
  AND2X1_RVT U132 ( .A1(n200), .A2(m4stg_inc_exp_55), .Y(m4stg_left_shift_step) );
  AND2X1_RVT U133 ( .A1(m4stg_right_shift), .A2(n200), .Y(
        m4stg_right_shift_step) );
  INVX1_RVT U134 ( .A(\intadd_4/SUM[0] ), .Y(n165) );
  INVX1_RVT U135 ( .A(\intadd_4/SUM[1] ), .Y(n164) );
  INVX1_RVT U136 ( .A(\intadd_4/SUM[2] ), .Y(n163) );
  INVX1_RVT U137 ( .A(\intadd_4/SUM[3] ), .Y(n162) );
  INVX1_RVT U138 ( .A(\intadd_4/n1 ), .Y(n160) );
  INVX1_RVT U139 ( .A(\intadd_4/SUM[4] ), .Y(n161) );
  NAND2X0_RVT U140 ( .A1(m2stg_ld0_2[0]), .A2(m2stg_ld0_1[0]), .Y(n192) );
  INVX1_RVT U141 ( .A(n192), .Y(\intadd_4/CI ) );
  OR2X1_RVT U142 ( .A1(m1stg_snan_dbl_in1), .A2(m1stg_snan_sng_in1), .Y(
        m1stg_snan_in1) );
  INVX1_RVT U143 ( .A(m3stg_expadd_lte_0_inv), .Y(n188) );
  INVX1_RVT U144 ( .A(m3stg_exp[3]), .Y(n167) );
  INVX1_RVT U145 ( .A(m3stg_exp[4]), .Y(n146) );
  INVX1_RVT U146 ( .A(m3stg_exp[2]), .Y(n173) );
  INVX1_RVT U147 ( .A(\m3stg_exp_inv_plus2[1] ), .Y(n183) );
  NAND4X0_RVT U148 ( .A1(n167), .A2(n146), .A3(n173), .A4(n183), .Y(n140) );
  INVX1_RVT U149 ( .A(n140), .Y(n145) );
  NOR4X1_RVT U150 ( .A1(m3stg_exp[0]), .A2(m3stg_exp[10]), .A3(m3stg_exp[6]), 
        .A4(m3stg_exp[7]), .Y(n72) );
  NOR4X1_RVT U151 ( .A1(m3stg_exp[5]), .A2(m3stg_exp[11]), .A3(m3stg_exp[9]), 
        .A4(m3stg_exp[8]), .Y(n71) );
  OA222X1_RVT U152 ( .A1(m3stg_exp[12]), .A2(n145), .A3(m3stg_exp[12]), .A4(
        n72), .A5(m3stg_exp[12]), .A6(n71), .Y(n151) );
  NAND2X0_RVT U153 ( .A1(n188), .A2(n151), .Y(n181) );
  INVX1_RVT U154 ( .A(n181), .Y(m4stg_right_shift_in) );
  INVX1_RVT U155 ( .A(m5stg_to_0_inv), .Y(m5stg_to_0) );
  OA21X1_RVT U156 ( .A1(n75), .A2(n74), .A3(n73), .Y(m1stg_nan_in2) );
  NAND2X0_RVT U157 ( .A1(n77), .A2(n76), .Y(m1stg_snan_in2) );
  NAND2X0_RVT U164 ( .A1(n79), .A2(n78), .Y(m1stg_qnan_in2) );
  OR2X1_RVT U165 ( .A1(m1stg_inf_in2), .A2(m1stg_inf_in1), .Y(m1stg_inf_in) );
  INVX1_RVT U166 ( .A(m1stg_snan_in2), .Y(n124) );
  INVX1_RVT U167 ( .A(m1stg_nan_in2), .Y(n123) );
  AND2X1_RVT U168 ( .A1(m1stg_inf_in), .A2(n123), .Y(n85) );
  NAND2X0_RVT U169 ( .A1(n1), .A2(mul_exp_in1_exp_neq_ffs), .Y(n84) );
  AND2X1_RVT U170 ( .A1(n85), .A2(n84), .Y(n126) );
  NAND2X0_RVT U171 ( .A1(n86), .A2(m1stg_qnan_in2), .Y(n87) );
  NAND3X0_RVT U172 ( .A1(n124), .A2(n88), .A3(n87), .Y(m2stg_frac1_inf) );
  OR3X2_RVT U173 ( .A1(m4stg_right_shift), .A2(m4stg_exp[2]), .A3(
        m4stg_exp[11]), .Y(n92) );
  NOR4X1_RVT U174 ( .A1(m4stg_exp[1]), .A2(m4stg_exp[0]), .A3(m4stg_exp[5]), 
        .A4(m4stg_exp[3]), .Y(n90) );
  NOR4X1_RVT U175 ( .A1(m4stg_exp[4]), .A2(m4stg_exp[6]), .A3(m4stg_exp[8]), 
        .A4(m4stg_exp[10]), .Y(n89) );
  NAND2X0_RVT U176 ( .A1(n90), .A2(n89), .Y(n91) );
  NOR4X1_RVT U177 ( .A1(m4stg_exp[9]), .A2(m4stg_exp[7]), .A3(n92), .A4(n91), 
        .Y(m4stg_inc_exp_54) );
  AND2X1_RVT U180 ( .A1(mula_rst_l), .A2(n103), .Y(n94) );
  AND3X1_RVT U181 ( .A1(mula_rst_l), .A2(m1stg_step), .A3(inq_mul), .Y(n93) );
  AO22X1_RVT U182 ( .A1(m1stg_op[7]), .A2(n94), .A3(n93), .A4(inq_op[7]), .Y(
        m1stg_op_in[7]) );
  AO22X1_RVT U183 ( .A1(m1stg_op[6]), .A2(n94), .A3(n93), .A4(inq_op[6]), .Y(
        m1stg_op_in[6]) );
  AO22X1_RVT U184 ( .A1(m1stg_op[5]), .A2(n94), .A3(n93), .A4(inq_op[5]), .Y(
        m1stg_op_in[5]) );
  AO22X1_RVT U185 ( .A1(m1stg_op[4]), .A2(n94), .A3(n93), .A4(inq_op[4]), .Y(
        m1stg_op_in[4]) );
  AO22X1_RVT U186 ( .A1(m1stg_op[3]), .A2(n94), .A3(n93), .A4(inq_op[3]), .Y(
        m1stg_op_in[3]) );
  AO22X1_RVT U187 ( .A1(m1stg_op[2]), .A2(n94), .A3(n93), .A4(inq_op[2]), .Y(
        m1stg_op_in[2]) );
  AO22X1_RVT U188 ( .A1(m1stg_op[1]), .A2(n94), .A3(n93), .A4(inq_op[1]), .Y(
        m1stg_op_in[1]) );
  AO22X1_RVT U189 ( .A1(m1stg_op[0]), .A2(n94), .A3(n93), .A4(inq_op[0]), .Y(
        m1stg_op_in[0]) );
  AO21X1_RVT U190 ( .A1(m1stg_mul), .A2(n94), .A3(n93), .Y(m1stg_mul_in) );
  OA21X1_RVT U191 ( .A1(m5stg_opdec[4]), .A2(n103), .A3(mula_rst_l), .Y(
        m6stg_fmul_in) );
  AND2X1_RVT U192 ( .A1(m5stg_id[3]), .A2(n200), .Y(n99) );
  AND2X1_RVT U193 ( .A1(m5stg_id[2]), .A2(m5stg_id[4]), .Y(n95) );
  AO22X1_RVT U194 ( .A1(n103), .A2(m6stg_id[9]), .A3(n99), .A4(n95), .Y(
        m6stg_id_in[9]) );
  INVX1_RVT U195 ( .A(m5stg_id[2]), .Y(n98) );
  AND2X1_RVT U196 ( .A1(m5stg_id[4]), .A2(n98), .Y(n96) );
  AO22X1_RVT U197 ( .A1(n103), .A2(m6stg_id[8]), .A3(n99), .A4(n96), .Y(
        m6stg_id_in[8]) );
  NOR2X0_RVT U198 ( .A1(n103), .A2(m5stg_id[3]), .Y(n102) );
  AO22X1_RVT U199 ( .A1(n103), .A2(m6stg_id[7]), .A3(n95), .A4(n102), .Y(
        m6stg_id_in[7]) );
  AO22X1_RVT U200 ( .A1(n103), .A2(m6stg_id[6]), .A3(n96), .A4(n102), .Y(
        m6stg_id_in[6]) );
  INVX1_RVT U201 ( .A(m5stg_id[4]), .Y(n97) );
  AND2X1_RVT U202 ( .A1(m5stg_id[2]), .A2(n97), .Y(n100) );
  AO22X1_RVT U203 ( .A1(n103), .A2(m6stg_id[5]), .A3(n99), .A4(n100), .Y(
        m6stg_id_in[5]) );
  AND2X1_RVT U204 ( .A1(n98), .A2(n97), .Y(n101) );
  AO22X1_RVT U205 ( .A1(n103), .A2(m6stg_id[4]), .A3(n99), .A4(n101), .Y(
        m6stg_id_in[4]) );
  AO22X1_RVT U206 ( .A1(n103), .A2(m6stg_id[3]), .A3(n102), .A4(n100), .Y(
        m6stg_id_in[3]) );
  AO22X1_RVT U207 ( .A1(n103), .A2(m6stg_id[2]), .A3(n102), .A4(n101), .Y(
        m6stg_id_in[2]) );
  AO22X1_RVT U208 ( .A1(n103), .A2(m6stg_id[1]), .A3(n200), .A4(m5stg_id[1]), 
        .Y(m6stg_id_in[1]) );
  AO22X1_RVT U209 ( .A1(n103), .A2(m6stg_id[0]), .A3(n200), .A4(m5stg_id[0]), 
        .Y(m6stg_id_in[0]) );
  NOR4X1_RVT U210 ( .A1(m3bstg_opdec[4]), .A2(m3stg_opdec[4]), .A3(
        m4stg_opdec[4]), .A4(m2stg_opdec[4]), .Y(n105) );
  NOR4X1_RVT U211 ( .A1(m3astg_opdec[4]), .A2(\m6stg_opdec[4] ), .A3(
        m5stg_opdec[4]), .A4(m1stg_fmul), .Y(n104) );
  NAND2X0_RVT U212 ( .A1(n105), .A2(n104), .Y(mul_pipe_active_in) );
  OR2X1_RVT U213 ( .A1(m2stg_snan_in2), .A2(m2stg_snan_in1), .Y(n106) );
  AND2X1_RVT U214 ( .A1(n106), .A2(m2stg_sign2), .Y(n108) );
  NAND2X0_RVT U215 ( .A1(m2stg_qnan_in1), .A2(m2stg_nan_in2), .Y(n107) );
  AND2X1_RVT U216 ( .A1(n108), .A2(n107), .Y(n112) );
  NAND2X0_RVT U217 ( .A1(m2stg_snan_in1), .A2(m2stg_qnan_in2), .Y(n109) );
  AND3X1_RVT U218 ( .A1(n113), .A2(m2stg_sign1), .A3(n109), .Y(n111) );
  AOI22X1_RVT U219 ( .A1(m2stg_zero_in), .A2(m2stg_inf_in), .A3(n112), .A4(
        n111), .Y(n110) );
  OA21X1_RVT U220 ( .A1(n112), .A2(n111), .A3(n110), .Y(m2stg_sign) );
  AOI22X1_RVT U221 ( .A1(m2stg_zero_in2), .A2(m2stg_inf_in1), .A3(
        m2stg_inf_in2), .A4(m2stg_zero_in1), .Y(n114) );
  NAND3X0_RVT U222 ( .A1(m2stg_snan_in1), .A2(n114), .A3(n113), .Y(m2stg_nv)
         );
  AND4X1_RVT U223 ( .A1(m5stg_of_mask), .A2(n191), .A3(n116), .A4(n115), .Y(
        mul_of_out_tmp1_in) );
  NOR4X1_RVT U224 ( .A1(m5stg_exp[1]), .A2(m5stg_exp[2]), .A3(m5stg_exp[7]), 
        .A4(m5stg_exp[3]), .Y(n120) );
  OR2X1_RVT U225 ( .A1(m5stg_exp[6]), .A2(m5stg_exp[4]), .Y(n117) );
  NOR4X1_RVT U226 ( .A1(m5stg_exp[5]), .A2(m5stg_exp[0]), .A3(n118), .A4(n117), 
        .Y(n119) );
  OA221X1_RVT U227 ( .A1(m5stg_exp[12]), .A2(n120), .A3(m5stg_exp[12]), .A4(
        n119), .A5(m5stg_frac_neq_0), .Y(mul_uf_out_in) );
  AO22X1_RVT U228 ( .A1(m5stg_fmuls), .A2(m5stg_frac_sng_nx), .A3(m5stg_fmuld), 
        .A4(m5stg_frac_dbl_nx), .Y(mul_nx_out_in) );
  AO21X1_RVT U229 ( .A1(mul_of_out_cout), .A2(mul_of_out_tmp1), .A3(
        mul_of_out_tmp2), .Y(mul_exc_out[3]) );
  OR2X1_RVT U230 ( .A1(mul_nx_out), .A2(mul_exc_out[3]), .Y(mul_exc_out_0) );
  NAND2X0_RVT U231 ( .A1(n122), .A2(n121), .Y(m1stg_qnan_in1) );
  AO22X1_RVT U232 ( .A1(n124), .A2(m1stg_snan_in1), .A3(n123), .A4(
        m1stg_qnan_in1), .Y(n125) );
  OR2X1_RVT U233 ( .A1(n126), .A2(n125), .Y(m2stg_frac2_inf) );
  AND2X1_RVT U234 ( .A1(n135), .A2(m1stg_op[5]), .Y(m1stg_fsmuld) );
  OR2X1_RVT U235 ( .A1(m1stg_fsmuld), .A2(n157), .Y(\m1stg_opdec[3] ) );
  AND2X1_RVT U236 ( .A1(\m1stg_opdec[3] ), .A2(m1stg_inf_zero_in), .Y(
        m1stg_inf_zero_in_dbl) );
  AND2X1_RVT U237 ( .A1(n154), .A2(mul_exp_in1_exp_eq_0), .Y(n129) );
  NAND2X0_RVT U238 ( .A1(n128), .A2(n127), .Y(n131) );
  AND2X1_RVT U239 ( .A1(n129), .A2(n131), .Y(n130) );
  AND2X1_RVT U240 ( .A1(n130), .A2(m1stg_ld0_1[5]), .Y(m2stg_ld0_1_in[5]) );
  AND2X1_RVT U241 ( .A1(n130), .A2(m1stg_ld0_1[4]), .Y(m2stg_ld0_1_in[4]) );
  AND2X1_RVT U242 ( .A1(n130), .A2(m1stg_ld0_1[3]), .Y(m2stg_ld0_1_in[3]) );
  AND2X1_RVT U243 ( .A1(n130), .A2(m1stg_ld0_1[2]), .Y(m2stg_ld0_1_in[2]) );
  AND2X1_RVT U244 ( .A1(n130), .A2(m1stg_ld0_1[1]), .Y(m2stg_ld0_1_in[1]) );
  AND2X1_RVT U245 ( .A1(n130), .A2(m1stg_ld0_1[0]), .Y(m2stg_ld0_1_in[0]) );
  AND2X1_RVT U246 ( .A1(n154), .A2(mul_exp_in2_exp_eq_0), .Y(n132) );
  AND2X1_RVT U247 ( .A1(n132), .A2(n131), .Y(n133) );
  AND2X1_RVT U248 ( .A1(n133), .A2(m1stg_ld0_2[5]), .Y(m2stg_ld0_2_in[5]) );
  AND2X1_RVT U249 ( .A1(n133), .A2(m1stg_ld0_2[4]), .Y(m2stg_ld0_2_in[4]) );
  AND2X1_RVT U250 ( .A1(n133), .A2(m1stg_ld0_2[3]), .Y(m2stg_ld0_2_in[3]) );
  AND2X1_RVT U251 ( .A1(n133), .A2(m1stg_ld0_2[2]), .Y(m2stg_ld0_2_in[2]) );
  AND2X1_RVT U252 ( .A1(n133), .A2(m1stg_ld0_2[1]), .Y(m2stg_ld0_2_in[1]) );
  AND2X1_RVT U253 ( .A1(n133), .A2(m1stg_ld0_2[0]), .Y(m2stg_ld0_2_in[0]) );
  AND2X1_RVT U254 ( .A1(n157), .A2(n136), .Y(m2stg_exp_0bff) );
  AND2X1_RVT U255 ( .A1(n135), .A2(n134), .Y(n155) );
  AND2X1_RVT U256 ( .A1(n155), .A2(n136), .Y(m2stg_exp_017f) );
  AND2X1_RVT U257 ( .A1(m1stg_fsmuld), .A2(n136), .Y(m2stg_exp_04ff) );
  AND2X1_RVT U258 ( .A1(n154), .A2(m1stg_zero_in), .Y(m2stg_exp_zero) );
  INVX1_RVT U259 ( .A(n151), .Y(n156) );
  NAND2X0_RVT U260 ( .A1(n156), .A2(n188), .Y(n185) );
  NAND2X0_RVT U261 ( .A1(n173), .A2(n183), .Y(n176) );
  NOR2X0_RVT U262 ( .A1(n176), .A2(m3stg_exp[0]), .Y(n152) );
  NAND2X0_RVT U263 ( .A1(n152), .A2(n167), .Y(n158) );
  INVX1_RVT U264 ( .A(n158), .Y(n147) );
  NAND2X0_RVT U265 ( .A1(n146), .A2(n147), .Y(n148) );
  HADDX1_RVT U266 ( .A0(m3stg_exp[5]), .B0(n148), .SO(n137) );
  OA22X1_RVT U267 ( .A1(m3stg_ld0_inv[5]), .A2(n188), .A3(n185), .A4(n137), 
        .Y(n143) );
  AND4X1_RVT U268 ( .A1(m3stg_exp[9]), .A2(m3stg_exp[8]), .A3(m3stg_exp[10]), 
        .A4(m3stg_exp[6]), .Y(n139) );
  INVX1_RVT U269 ( .A(m3stg_exp[5]), .Y(n141) );
  NAND3X0_RVT U270 ( .A1(n167), .A2(n146), .A3(n141), .Y(n138) );
  NAND4X0_RVT U271 ( .A1(m3stg_exp[7]), .A2(m3stg_exp[11]), .A3(n139), .A4(
        n138), .Y(n180) );
  NAND3X0_RVT U272 ( .A1(m3stg_exp[12]), .A2(n188), .A3(n180), .Y(n189) );
  AO221X1_RVT U273 ( .A1(n145), .A2(n141), .A3(n140), .A4(m3stg_exp[5]), .A5(
        n181), .Y(n142) );
  NAND3X0_RVT U274 ( .A1(n143), .A2(n189), .A3(n142), .Y(m4stg_sh_cnt_in[5])
         );
  AO221X1_RVT U275 ( .A1(m3stg_exp[4]), .A2(m3stg_exp[3]), .A3(m3stg_exp[4]), 
        .A4(n176), .A5(n181), .Y(n144) );
  OA22X1_RVT U276 ( .A1(n145), .A2(n144), .A3(m3stg_ld0_inv[4]), .A4(n188), 
        .Y(n150) );
  AO221X1_RVT U277 ( .A1(n148), .A2(n147), .A3(n148), .A4(n146), .A5(n185), 
        .Y(n149) );
  NAND3X0_RVT U278 ( .A1(n150), .A2(n189), .A3(n149), .Y(m4stg_sh_cnt_in[4])
         );
  AO221X1_RVT U279 ( .A1(n156), .A2(n152), .A3(n151), .A4(n176), .A5(
        m3stg_expadd_lte_0_inv), .Y(n159) );
  OA22X1_RVT U280 ( .A1(n159), .A2(n167), .A3(n185), .A4(n158), .Y(n172) );
  NAND3X0_RVT U281 ( .A1(m4stg_right_shift_in), .A2(n167), .A3(n176), .Y(n171)
         );
  OR2X1_RVT U282 ( .A1(m3stg_ld0_inv[3]), .A2(n188), .Y(n170) );
  NAND4X0_RVT U283 ( .A1(n172), .A2(n171), .A3(n189), .A4(n170), .Y(
        m4stg_sh_cnt_in[3]) );
  OA222X1_RVT U284 ( .A1(n173), .A2(n183), .A3(n173), .A4(n182), .A5(
        m3stg_exp[0]), .A6(n176), .Y(n174) );
  OA22X1_RVT U285 ( .A1(n174), .A2(n185), .A3(m3stg_ld0_inv[2]), .A4(n188), 
        .Y(n179) );
  NAND2X0_RVT U286 ( .A1(m3stg_exp[2]), .A2(\m3stg_exp_inv_plus2[1] ), .Y(n175) );
  NAND4X0_RVT U287 ( .A1(m4stg_right_shift_in), .A2(n177), .A3(n176), .A4(n175), .Y(n178) );
  NAND2X0_RVT U288 ( .A1(n179), .A2(n178), .Y(m4stg_sh_cnt_in[2]) );
  OA22X1_RVT U289 ( .A1(n182), .A2(n185), .A3(n181), .A4(n180), .Y(n184) );
  OA22X1_RVT U290 ( .A1(n184), .A2(n183), .A3(m3stg_ld0_inv[1]), .A4(n188), 
        .Y(n187) );
  NAND2X0_RVT U291 ( .A1(n187), .A2(n186), .Y(m4stg_sh_cnt_in[1]) );
  AO22X1_RVT U292 ( .A1(m3stg_expadd_lte_0_inv), .A2(m3stg_ld0_inv[0]), .A3(
        n188), .A4(m3stg_exp[0]), .Y(n190) );
  NAND2X0_RVT U293 ( .A1(n190), .A2(n189), .Y(m4stg_sh_cnt_in[0]) );
  AND3X1_RVT U294 ( .A1(m4stg_right_shift), .A2(m4stg_frac_105), .A3(
        m4stg_expadd_eq_0), .Y(m4stg_inc_exp_105) );
  NOR2X0_RVT U295 ( .A1(n191), .A2(m5stg_in_of), .Y(mul_frac_out_frac) );
  OAI21X1_RVT U296 ( .A1(m2stg_ld0_2[0]), .A2(m2stg_ld0_1[0]), .A3(n192), .Y(
        n166) );
endmodule


module clken_buf_9 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_5 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_5 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_4 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_4 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_8 ( din, en, clk, se, si, so, \q[12] , \q[11]_BAR , \q[9] , 
        \q[8] , \q[7] , \q[6] , \q[5] , \q[4] , \q[3] , \q[2] , \q[1] , \q[0] , 
        \q[10]_BAR  );
  input [12:0] din;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  output \q[12] , \q[11]_BAR , \q[9] , \q[8] , \q[7] , \q[6] , \q[5] , \q[4] ,
         \q[3] , \q[2] , \q[1] , \q[0] , \q[10]_BAR ;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n4, n5;
  wire   [12:0] q;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_8 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .QN(\q[11]_BAR ) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .QN(\q[10]_BAR ) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n4) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n4), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n4), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n4), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n4), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n4), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n4), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n4), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n4), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n4), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n4), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n4), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n4), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n4), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_7 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_7 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_6 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_6 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_5 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2, n4;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_5 clk_gate_q_reg ( .CLK(clk), .EN(n4), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  INVX1_RVT U14 ( .A(se), .Y(n2) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n2), .Y(N15) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  OR2X1_RVT U18 ( .A1(se), .A2(en), .Y(n4) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_4 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_4 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_3 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, net24246, n1,
         n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_3 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N15) );
  OR2X1_RVT U16 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dff_SIZE13_3 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, n1;

  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
endmodule


module dff_SIZE13_2 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, n1;

  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
endmodule


module dff_SIZE13_1 ( din, clk, se, si, so, \q[12]_BAR , \q[11]_BAR , 
        \q[10]_BAR , \q[9]_BAR , \q[8]_BAR , \q[7]_BAR , \q[6]_BAR , 
        \q[5]_BAR , \q[4]_BAR , \q[3]_BAR , \q[2]_BAR , \q[1]_BAR , \q[0]_BAR 
 );
  input [12:0] din;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  output \q[12]_BAR , \q[11]_BAR , \q[10]_BAR , \q[9]_BAR , \q[8]_BAR ,
         \q[7]_BAR , \q[6]_BAR , \q[5]_BAR , \q[4]_BAR , \q[3]_BAR ,
         \q[2]_BAR , \q[1]_BAR , \q[0]_BAR ;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, n1;

  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .QN(\q[12]_BAR ) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .QN(\q[11]_BAR ) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .QN(\q[10]_BAR ) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .QN(\q[9]_BAR ) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .QN(\q[8]_BAR ) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .QN(\q[7]_BAR ) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .QN(\q[6]_BAR ) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .QN(\q[5]_BAR ) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .QN(\q[4]_BAR ) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .QN(\q[3]_BAR ) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .QN(\q[2]_BAR ) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .QN(\q[1]_BAR ) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .QN(\q[0]_BAR ) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
endmodule


module dff_SIZE5_1 ( din, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, n1;

  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_3 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_3 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module fpu_mul_exp_dp ( inq_in1, inq_in2, m6stg_step, m1stg_dblop, m1stg_sngop, 
        m2stg_exp_expadd, m2stg_exp_0bff, m2stg_exp_017f, m2stg_exp_04ff, 
        m2stg_exp_zero, m1stg_fsmuld, m2stg_fmuld, m2stg_fmuls, m2stg_fsmuld, 
        m3stg_ld0_inv, m5stg_fracadd_cout, mul_exp_out_exp_plus1, 
        mul_exp_out_exp, m5stg_in_of, m5stg_fmuld, m5stg_to_0_inv, 
        m4stg_shl_54, m4stg_shl_55, m4stg_inc_exp_54, m4stg_inc_exp_55, 
        m4stg_inc_exp_105, fmul_clken_l, rclk, m3stg_exp, m3stg_expadd_eq_0, 
        m3stg_expadd_lte_0_inv, m4stg_exp, m5stg_exp, mul_exp_out, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [6:0] m3stg_ld0_inv;
  output [12:0] m3stg_exp;
  output [12:0] m4stg_exp;
  output [12:0] m5stg_exp;
  output [10:0] mul_exp_out;
  input m6stg_step, m1stg_dblop, m1stg_sngop, m2stg_exp_expadd, m2stg_exp_0bff,
         m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero, m1stg_fsmuld,
         m2stg_fmuld, m2stg_fmuls, m2stg_fsmuld, m5stg_fracadd_cout,
         mul_exp_out_exp_plus1, mul_exp_out_exp, m5stg_in_of, m5stg_fmuld,
         m5stg_to_0_inv, m4stg_shl_54, m4stg_shl_55, m4stg_inc_exp_54,
         m4stg_inc_exp_55, m4stg_inc_exp_105, fmul_clken_l, rclk, se, si;
  output m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv, so;
  wire   clk, m5stg_shl_55, m5stg_shl_54, m5stg_inc_exp_54, m5stg_inc_exp_55,
         m5stg_inc_exp_105, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, \intadd_7/B[0] , \intadd_7/CI , \intadd_7/SUM[1] ,
         \intadd_7/SUM[0] , \intadd_7/n3 , \intadd_7/n2 , \intadd_5/A[9] ,
         \intadd_5/A[8] , \intadd_5/A[7] , \intadd_5/A[6] , \intadd_5/A[5] ,
         \intadd_5/A[4] , \intadd_5/A[3] , \intadd_5/A[2] , \intadd_5/A[1] ,
         \intadd_5/A[0] , \intadd_5/B[9] , \intadd_5/B[8] , \intadd_5/B[7] ,
         \intadd_5/B[6] , \intadd_5/B[5] , \intadd_5/B[4] , \intadd_5/B[3] ,
         \intadd_5/B[2] , \intadd_5/B[1] , \intadd_5/B[0] , \intadd_5/CI ,
         \intadd_5/SUM[9] , \intadd_5/SUM[8] , \intadd_5/SUM[7] ,
         \intadd_5/SUM[6] , \intadd_5/SUM[5] , \intadd_5/SUM[4] ,
         \intadd_5/SUM[3] , \intadd_5/SUM[2] , \intadd_5/SUM[1] ,
         \intadd_5/SUM[0] , \intadd_5/n10 , \intadd_5/n9 , \intadd_5/n8 ,
         \intadd_5/n7 , \intadd_5/n6 , \intadd_5/n5 , \intadd_5/n4 ,
         \intadd_5/n3 , \intadd_5/n2 , \intadd_5/n1 , \intadd_6/CI ,
         \intadd_6/SUM[5] , \intadd_6/SUM[4] , \intadd_6/SUM[3] ,
         \intadd_6/SUM[2] , \intadd_6/SUM[1] , \intadd_6/SUM[0] ,
         \intadd_6/n6 , \intadd_6/n5 , \intadd_6/n4 , \intadd_6/n3 ,
         \intadd_6/n2 , \intadd_6/n1 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156;
  wire   [10:0] m1stg_exp_in1;
  wire   [10:0] m1stg_exp_in2;
  wire   [12:0] m2stg_exp_in;
  wire   [12:0] m2stg_exp;
  wire   [12:0] m2stg_expadd;
  wire   [12:0] m3astg_exp;
  wire   [12:0] m3bstg_exp;
  wire   [12:0] m3stg_expa;
  wire   [12:0] m4stg_exp_in;
  wire   [12:0] m5stg_exp_pre1_in;
  wire   [12:0] m5stg_exp_pre1;
  wire   [12:0] m5stg_exp_pre2_in;
  wire   [12:0] m5stg_exp_pre2;
  wire   [12:0] m5stg_exp_pre3;
  wire   [10:0] mul_exp_out_in;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign so = 1'b0;

  clken_buf_9 ckbuf_mul_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fmul_clken_l), 
        .tmb_l(n156) );
  dffe_SIZE11_5 i_m1stg_exp_in1 ( .din(inq_in1), .en(m6stg_step), .clk(clk), 
        .q(m1stg_exp_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_4 i_m1stg_exp_in2 ( .din(inq_in2), .en(m6stg_step), .clk(clk), 
        .q(m1stg_exp_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_8 i_m2stg_exp ( .din(m2stg_exp_in), .en(m6stg_step), .clk(clk), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .\q[12] (m2stg_exp[12]), .\q[11]_BAR (
        m2stg_exp[11]), .\q[9] (m2stg_exp[9]), .\q[8] (m2stg_exp[8]), .\q[7] (
        m2stg_exp[7]), .\q[6] (m2stg_expadd[6]), .\q[5] (m2stg_expadd[5]), 
        .\q[4] (m2stg_expadd[4]), .\q[3] (m2stg_expadd[3]), .\q[2] (
        m2stg_expadd[2]), .\q[1] (m2stg_expadd[1]), .\q[0] (m2stg_expadd[0]), 
        .\q[10]_BAR (m2stg_exp[10]) );
  dffe_SIZE13_7 i_m3astg_exp ( .din(m2stg_expadd), .en(m6stg_step), .clk(clk), 
        .q(m3astg_exp), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_6 i_m3bstg_exp ( .din(m3astg_exp), .en(m6stg_step), .clk(clk), 
        .q(m3bstg_exp), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_5 i_m3stg_exp ( .din(m3bstg_exp), .en(m6stg_step), .clk(clk), 
        .q(m3stg_exp), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_4 i_m3stg_expa ( .din(m3bstg_exp), .en(m6stg_step), .clk(clk), 
        .q(m3stg_expa), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_3 i_m4stg_exp ( .din({1'b0, m4stg_exp_in[11:0]}), .en(m6stg_step), .clk(clk), .q({SYNOPSYS_UNCONNECTED__0, m4stg_exp[11:0]}), .se(se), .si({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dff_SIZE13_3 i_m5stg_exp_pre1 ( .din(m5stg_exp_pre1_in), .clk(clk), .q(
        m5stg_exp_pre1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE13_2 i_m5stg_exp_pre2 ( .din({1'b0, m5stg_exp_pre2_in[11:0]}), .clk(
        clk), .q({SYNOPSYS_UNCONNECTED__1, m5stg_exp_pre2[11:0]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  dff_SIZE13_1 i_m5stg_exp_pre3 ( .din({n69, n68, n67, n66, n65, n64, n63, n62, 
        n61, n60, n59, n58, n57}), .clk(clk), .se(se), .si({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .\q[12]_BAR (m5stg_exp_pre3[12]), .\q[11]_BAR (m5stg_exp_pre3[11]), 
        .\q[10]_BAR (m5stg_exp_pre3[10]), .\q[9]_BAR (m5stg_exp_pre3[9]), 
        .\q[8]_BAR (m5stg_exp_pre3[8]), .\q[7]_BAR (m5stg_exp_pre3[7]), 
        .\q[6]_BAR (m5stg_exp_pre3[6]), .\q[5]_BAR (m5stg_exp_pre3[5]), 
        .\q[4]_BAR (m5stg_exp_pre3[4]), .\q[3]_BAR (m5stg_exp_pre3[3]), 
        .\q[2]_BAR (m5stg_exp_pre3[2]), .\q[1]_BAR (m5stg_exp_pre3[1]), 
        .\q[0]_BAR (m5stg_exp_pre3[0]) );
  dff_SIZE5_1 i_m5stg_inc_exp ( .din({m4stg_shl_55, m4stg_shl_54, 
        m4stg_inc_exp_54, m4stg_inc_exp_55, m4stg_inc_exp_105}), .clk(clk), 
        .q({m5stg_shl_55, m5stg_shl_54, m5stg_inc_exp_54, m5stg_inc_exp_55, 
        m5stg_inc_exp_105}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_3 i_mul_exp_out ( .din(mul_exp_out_in), .en(m6stg_step), .clk(
        clk), .q(mul_exp_out), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  FADDX1_RVT \intadd_7/U4  ( .A(\intadd_7/B[0] ), .B(m2stg_exp[10]), .CI(
        \intadd_7/CI ), .CO(\intadd_7/n3 ), .S(\intadd_7/SUM[0] ) );
  FADDX1_RVT \intadd_7/U3  ( .A(\intadd_7/CI ), .B(m2stg_exp[11]), .CI(
        \intadd_7/n3 ), .CO(\intadd_7/n2 ), .S(\intadd_7/SUM[1] ) );
  FADDX1_RVT \intadd_5/U11  ( .A(\intadd_5/B[0] ), .B(\intadd_5/A[0] ), .CI(
        \intadd_5/CI ), .CO(\intadd_5/n10 ), .S(\intadd_5/SUM[0] ) );
  FADDX1_RVT \intadd_5/U10  ( .A(\intadd_5/B[1] ), .B(\intadd_5/A[1] ), .CI(
        \intadd_5/n10 ), .CO(\intadd_5/n9 ), .S(\intadd_5/SUM[1] ) );
  FADDX1_RVT \intadd_5/U9  ( .A(\intadd_5/B[2] ), .B(\intadd_5/A[2] ), .CI(
        \intadd_5/n9 ), .CO(\intadd_5/n8 ), .S(\intadd_5/SUM[2] ) );
  FADDX1_RVT \intadd_5/U8  ( .A(\intadd_5/B[3] ), .B(\intadd_5/A[3] ), .CI(
        \intadd_5/n8 ), .CO(\intadd_5/n7 ), .S(\intadd_5/SUM[3] ) );
  FADDX1_RVT \intadd_5/U7  ( .A(\intadd_5/B[4] ), .B(\intadd_5/A[4] ), .CI(
        \intadd_5/n7 ), .CO(\intadd_5/n6 ), .S(\intadd_5/SUM[4] ) );
  FADDX1_RVT \intadd_5/U6  ( .A(\intadd_5/B[5] ), .B(\intadd_5/A[5] ), .CI(
        \intadd_5/n6 ), .CO(\intadd_5/n5 ), .S(\intadd_5/SUM[5] ) );
  FADDX1_RVT \intadd_5/U5  ( .A(\intadd_5/B[6] ), .B(\intadd_5/A[6] ), .CI(
        \intadd_5/n5 ), .CO(\intadd_5/n4 ), .S(\intadd_5/SUM[6] ) );
  FADDX1_RVT \intadd_5/U4  ( .A(\intadd_5/B[7] ), .B(\intadd_5/A[7] ), .CI(
        \intadd_5/n4 ), .CO(\intadd_5/n3 ), .S(\intadd_5/SUM[7] ) );
  FADDX1_RVT \intadd_5/U3  ( .A(\intadd_5/B[8] ), .B(\intadd_5/A[8] ), .CI(
        \intadd_5/n3 ), .CO(\intadd_5/n2 ), .S(\intadd_5/SUM[8] ) );
  FADDX1_RVT \intadd_5/U2  ( .A(\intadd_5/B[9] ), .B(\intadd_5/A[9] ), .CI(
        \intadd_5/n2 ), .CO(\intadd_5/n1 ), .S(\intadd_5/SUM[9] ) );
  FADDX1_RVT \intadd_6/U7  ( .A(m3stg_expa[1]), .B(m3stg_ld0_inv[1]), .CI(
        \intadd_6/CI ), .CO(\intadd_6/n6 ), .S(\intadd_6/SUM[0] ) );
  FADDX1_RVT \intadd_6/U6  ( .A(m3stg_expa[2]), .B(m3stg_ld0_inv[2]), .CI(
        \intadd_6/n6 ), .CO(\intadd_6/n5 ), .S(\intadd_6/SUM[1] ) );
  FADDX1_RVT \intadd_6/U5  ( .A(m3stg_expa[3]), .B(m3stg_ld0_inv[3]), .CI(
        \intadd_6/n5 ), .CO(\intadd_6/n4 ), .S(\intadd_6/SUM[2] ) );
  FADDX1_RVT \intadd_6/U4  ( .A(m3stg_expa[4]), .B(m3stg_ld0_inv[4]), .CI(
        \intadd_6/n4 ), .CO(\intadd_6/n3 ), .S(\intadd_6/SUM[3] ) );
  FADDX1_RVT \intadd_6/U3  ( .A(m3stg_expa[5]), .B(m3stg_ld0_inv[5]), .CI(
        \intadd_6/n3 ), .CO(\intadd_6/n2 ), .S(\intadd_6/SUM[4] ) );
  FADDX1_RVT \intadd_6/U2  ( .A(m3stg_expa[6]), .B(m3stg_ld0_inv[6]), .CI(
        \intadd_6/n2 ), .CO(\intadd_6/n1 ), .S(\intadd_6/SUM[5] ) );
  OR3X1_RVT U3 ( .A1(m5stg_exp[10]), .A2(n104), .A3(n103), .Y(n100) );
  INVX0_RVT U4 ( .A(n142), .Y(n143) );
  INVX0_RVT U5 ( .A(n50), .Y(n51) );
  INVX0_RVT U6 ( .A(n52), .Y(n53) );
  INVX0_RVT U7 ( .A(n78), .Y(n38) );
  INVX0_RVT U8 ( .A(n54), .Y(n55) );
  INVX0_RVT U9 ( .A(n56), .Y(n70) );
  INVX0_RVT U10 ( .A(m5stg_in_of), .Y(n140) );
  OR3X1_RVT U11 ( .A1(m3stg_expa[8]), .A2(m3stg_expa[7]), .A3(\intadd_6/n1 ), 
        .Y(n56) );
  INVX0_RVT U12 ( .A(n82), .Y(n33) );
  INVX0_RVT U13 ( .A(m5stg_exp[0]), .Y(n145) );
  INVX0_RVT U14 ( .A(m5stg_exp[1]), .Y(n139) );
  INVX0_RVT U15 ( .A(m5stg_exp[2]), .Y(n134) );
  INVX0_RVT U16 ( .A(n86), .Y(n28) );
  INVX0_RVT U17 ( .A(m5stg_exp[6]), .Y(n117) );
  INVX0_RVT U18 ( .A(m5stg_exp[7]), .Y(n115) );
  INVX0_RVT U19 ( .A(m5stg_exp[4]), .Y(n125) );
  INVX0_RVT U20 ( .A(m5stg_exp[5]), .Y(n124) );
  INVX0_RVT U21 ( .A(m5stg_exp[3]), .Y(n132) );
  INVX0_RVT U22 ( .A(m5stg_exp[8]), .Y(n106) );
  INVX0_RVT U23 ( .A(m5stg_exp[9]), .Y(n103) );
  INVX0_RVT U24 ( .A(m5stg_exp[10]), .Y(n99) );
  INVX0_RVT U25 ( .A(n84), .Y(m5stg_exp_pre2_in[8]) );
  INVX0_RVT U26 ( .A(n88), .Y(m5stg_exp_pre2_in[6]) );
  INVX0_RVT U27 ( .A(n91), .Y(m5stg_exp_pre2_in[4]) );
  INVX0_RVT U28 ( .A(n80), .Y(m5stg_exp_pre2_in[10]) );
  INVX0_RVT U29 ( .A(m2stg_exp_04ff), .Y(n18) );
  INVX0_RVT U30 ( .A(m2stg_exp_017f), .Y(n15) );
  INVX0_RVT U31 ( .A(m4stg_exp[3]), .Y(n24) );
  INVX0_RVT U32 ( .A(m4stg_exp[5]), .Y(n29) );
  INVX0_RVT U33 ( .A(m4stg_exp[7]), .Y(n34) );
  INVX0_RVT U34 ( .A(m4stg_exp[9]), .Y(n39) );
  INVX0_RVT U35 ( .A(m4stg_exp[1]), .Y(n96) );
  INVX0_RVT U36 ( .A(m4stg_exp[2]), .Y(n93) );
  INVX0_RVT U37 ( .A(m4stg_exp[11]), .Y(n76) );
  NOR2X0_RVT U38 ( .A1(m2stg_fmuls), .A2(m2stg_fmuld), .Y(\intadd_7/CI ) );
  XOR2X1_RVT U39 ( .A1(\intadd_7/CI ), .A2(m2stg_exp[12]), .Y(n1) );
  XOR2X1_RVT U40 ( .A1(\intadd_7/n2 ), .A2(n1), .Y(m2stg_expadd[12]) );
  AOI22X1_RVT U41 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[1]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[4]), .Y(\intadd_5/CI ) );
  AOI22X1_RVT U42 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[1]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[4]), .Y(\intadd_5/B[0] ) );
  AOI22X1_RVT U43 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[2]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[5]), .Y(\intadd_5/A[1] ) );
  AOI22X1_RVT U44 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[2]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[5]), .Y(\intadd_5/B[1] ) );
  AOI22X1_RVT U45 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[3]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[6]), .Y(\intadd_5/A[2] ) );
  AOI22X1_RVT U46 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[3]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[6]), .Y(\intadd_5/B[2] ) );
  AOI22X1_RVT U47 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[4]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[7]), .Y(\intadd_5/A[3] ) );
  AOI22X1_RVT U48 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[4]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[7]), .Y(\intadd_5/B[3] ) );
  AOI22X1_RVT U49 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[5]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[8]), .Y(\intadd_5/A[4] ) );
  AOI22X1_RVT U50 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[5]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[8]), .Y(\intadd_5/B[4] ) );
  AOI22X1_RVT U51 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[6]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[9]), .Y(\intadd_5/A[5] ) );
  AOI22X1_RVT U52 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[6]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[9]), .Y(\intadd_5/B[5] ) );
  AOI22X1_RVT U53 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[7]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[10]), .Y(\intadd_5/A[6] ) );
  AOI22X1_RVT U54 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[7]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[10]), .Y(\intadd_5/B[6] ) );
  INVX1_RVT U55 ( .A(se), .Y(n156) );
  NAND2X0_RVT U56 ( .A1(m6stg_step), .A2(m4stg_exp[10]), .Y(n80) );
  NAND2X0_RVT U57 ( .A1(m6stg_step), .A2(m4stg_exp[4]), .Y(n91) );
  NAND2X0_RVT U58 ( .A1(m6stg_step), .A2(m4stg_exp[6]), .Y(n88) );
  NAND2X0_RVT U59 ( .A1(m6stg_step), .A2(m4stg_exp[8]), .Y(n84) );
  INVX1_RVT U60 ( .A(\intadd_7/SUM[0] ), .Y(m2stg_expadd[10]) );
  INVX1_RVT U61 ( .A(\intadd_7/SUM[1] ), .Y(m2stg_expadd[11]) );
  OR2X1_RVT U62 ( .A1(m3stg_ld0_inv[0]), .A2(m3stg_expa[0]), .Y(\intadd_6/CI )
         );
  HADDX1_RVT U63 ( .A0(m3stg_exp[5]), .B0(m3stg_ld0_inv[5]), .SO(n3) );
  NOR4X1_RVT U64 ( .A1(m3stg_exp[9]), .A2(m3stg_exp[10]), .A3(m3stg_exp[11]), 
        .A4(m3stg_exp[12]), .Y(n2) );
  NAND2X0_RVT U65 ( .A1(n3), .A2(n2), .Y(n11) );
  AOI22X1_RVT U66 ( .A1(m3stg_exp[3]), .A2(m3stg_ld0_inv[3]), .A3(m3stg_exp[6]), .A4(m3stg_ld0_inv[6]), .Y(n4) );
  OA221X1_RVT U67 ( .A1(m3stg_exp[3]), .A2(m3stg_ld0_inv[3]), .A3(m3stg_exp[6]), .A4(m3stg_ld0_inv[6]), .A5(n4), .Y(n9) );
  AOI22X1_RVT U68 ( .A1(m3stg_ld0_inv[0]), .A2(m3stg_exp[0]), .A3(
        m3stg_ld0_inv[4]), .A4(m3stg_exp[4]), .Y(n5) );
  OA221X1_RVT U69 ( .A1(m3stg_ld0_inv[0]), .A2(m3stg_exp[0]), .A3(
        m3stg_ld0_inv[4]), .A4(m3stg_exp[4]), .A5(n5), .Y(n8) );
  AOI22X1_RVT U70 ( .A1(m3stg_exp[2]), .A2(m3stg_ld0_inv[2]), .A3(m3stg_exp[1]), .A4(m3stg_ld0_inv[1]), .Y(n6) );
  OA221X1_RVT U71 ( .A1(m3stg_exp[2]), .A2(m3stg_ld0_inv[2]), .A3(m3stg_exp[1]), .A4(m3stg_ld0_inv[1]), .A5(n6), .Y(n7) );
  NAND3X0_RVT U72 ( .A1(n9), .A2(n8), .A3(n7), .Y(n10) );
  NOR4X1_RVT U73 ( .A1(m3stg_exp[7]), .A2(m3stg_exp[8]), .A3(n11), .A4(n10), 
        .Y(m3stg_expadd_eq_0) );
  AOI22X1_RVT U74 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[0]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in1[3]), .Y(n46) );
  AOI22X1_RVT U75 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[0]), .A3(m1stg_sngop), 
        .A4(m1stg_exp_in2[3]), .Y(n45) );
  NAND2X0_RVT U76 ( .A1(n46), .A2(n45), .Y(n47) );
  INVX1_RVT U77 ( .A(n47), .Y(\intadd_5/A[0] ) );
  AO22X1_RVT U78 ( .A1(m5stg_inc_exp_55), .A2(m5stg_shl_55), .A3(
        m5stg_inc_exp_54), .A4(m5stg_shl_54), .Y(n12) );
  OR2X1_RVT U79 ( .A1(m5stg_inc_exp_105), .A2(n12), .Y(n147) );
  INVX1_RVT U80 ( .A(n147), .Y(n148) );
  AO221X1_RVT U81 ( .A1(n148), .A2(m5stg_exp_pre2[8]), .A3(n147), .A4(
        m5stg_exp_pre1[8]), .A5(m5stg_exp_pre3[8]), .Y(m5stg_exp[8]) );
  AO221X1_RVT U82 ( .A1(n148), .A2(m5stg_exp_pre2[0]), .A3(n147), .A4(
        m5stg_exp_pre1[0]), .A5(m5stg_exp_pre3[0]), .Y(m5stg_exp[0]) );
  AO221X1_RVT U83 ( .A1(n148), .A2(m5stg_exp_pre2[1]), .A3(n147), .A4(
        m5stg_exp_pre1[1]), .A5(m5stg_exp_pre3[1]), .Y(m5stg_exp[1]) );
  AO221X1_RVT U84 ( .A1(n148), .A2(m5stg_exp_pre2[6]), .A3(n147), .A4(
        m5stg_exp_pre1[6]), .A5(m5stg_exp_pre3[6]), .Y(m5stg_exp[6]) );
  AO221X1_RVT U85 ( .A1(n148), .A2(m5stg_exp_pre2[4]), .A3(n147), .A4(
        m5stg_exp_pre1[4]), .A5(m5stg_exp_pre3[4]), .Y(m5stg_exp[4]) );
  AO221X1_RVT U86 ( .A1(n148), .A2(m5stg_exp_pre2[2]), .A3(n147), .A4(
        m5stg_exp_pre1[2]), .A5(m5stg_exp_pre3[2]), .Y(m5stg_exp[2]) );
  AO221X1_RVT U87 ( .A1(n148), .A2(m5stg_exp_pre2[5]), .A3(n147), .A4(
        m5stg_exp_pre1[5]), .A5(m5stg_exp_pre3[5]), .Y(m5stg_exp[5]) );
  AO221X1_RVT U88 ( .A1(n148), .A2(m5stg_exp_pre2[3]), .A3(n147), .A4(
        m5stg_exp_pre1[3]), .A5(m5stg_exp_pre3[3]), .Y(m5stg_exp[3]) );
  AO221X1_RVT U89 ( .A1(n148), .A2(m5stg_exp_pre2[7]), .A3(n147), .A4(
        m5stg_exp_pre1[7]), .A5(m5stg_exp_pre3[7]), .Y(m5stg_exp[7]) );
  AO221X1_RVT U90 ( .A1(n148), .A2(m5stg_exp_pre2[10]), .A3(n147), .A4(
        m5stg_exp_pre1[10]), .A5(m5stg_exp_pre3[10]), .Y(m5stg_exp[10]) );
  AO221X1_RVT U91 ( .A1(n148), .A2(m5stg_exp_pre2[9]), .A3(n147), .A4(
        m5stg_exp_pre1[9]), .A5(m5stg_exp_pre3[9]), .Y(m5stg_exp[9]) );
  AND2X1_RVT U92 ( .A1(m1stg_fsmuld), .A2(m2stg_exp_zero), .Y(m2stg_exp_in[12]) );
  INVX1_RVT U93 ( .A(m2stg_exp_0bff), .Y(n22) );
  INVX1_RVT U94 ( .A(\intadd_5/SUM[7] ), .Y(n13) );
  NAND2X0_RVT U95 ( .A1(m2stg_exp_expadd), .A2(n13), .Y(n14) );
  NAND3X0_RVT U96 ( .A1(n15), .A2(n22), .A3(n14), .Y(m2stg_exp_in[8]) );
  INVX1_RVT U97 ( .A(m2stg_exp_in[12]), .Y(n21) );
  INVX1_RVT U98 ( .A(\intadd_5/SUM[9] ), .Y(n16) );
  NAND2X0_RVT U99 ( .A1(m2stg_exp_expadd), .A2(n16), .Y(n17) );
  NAND3X0_RVT U100 ( .A1(n18), .A2(n21), .A3(n17), .Y(m2stg_exp_in[10]) );
  INVX1_RVT U101 ( .A(\intadd_5/n1 ), .Y(n19) );
  NAND2X0_RVT U102 ( .A1(m2stg_exp_expadd), .A2(n19), .Y(n20) );
  NAND3X0_RVT U103 ( .A1(n22), .A2(n21), .A3(n20), .Y(m2stg_exp_in[11]) );
  NAND4X0_RVT U104 ( .A1(m4stg_exp[3]), .A2(m4stg_exp[2]), .A3(m4stg_exp[0]), 
        .A4(m4stg_exp[1]), .Y(n27) );
  AND2X1_RVT U105 ( .A1(n27), .A2(m6stg_step), .Y(n26) );
  NAND3X0_RVT U106 ( .A1(m4stg_exp[2]), .A2(m4stg_exp[0]), .A3(m4stg_exp[1]), 
        .Y(n23) );
  NAND2X0_RVT U107 ( .A1(n24), .A2(n23), .Y(n25) );
  AND2X1_RVT U108 ( .A1(n26), .A2(n25), .Y(m5stg_exp_pre1_in[3]) );
  INVX1_RVT U109 ( .A(n27), .Y(n92) );
  AND2X1_RVT U110 ( .A1(m4stg_exp[4]), .A2(n92), .Y(n86) );
  NAND2X0_RVT U111 ( .A1(m4stg_exp[5]), .A2(n86), .Y(n32) );
  AND2X1_RVT U112 ( .A1(n32), .A2(m6stg_step), .Y(n31) );
  NAND2X0_RVT U113 ( .A1(n29), .A2(n28), .Y(n30) );
  AND2X1_RVT U114 ( .A1(n31), .A2(n30), .Y(m5stg_exp_pre1_in[5]) );
  INVX1_RVT U115 ( .A(n32), .Y(n89) );
  AND2X1_RVT U116 ( .A1(m4stg_exp[6]), .A2(n89), .Y(n82) );
  NAND2X0_RVT U117 ( .A1(m4stg_exp[7]), .A2(n82), .Y(n37) );
  AND2X1_RVT U118 ( .A1(n37), .A2(m6stg_step), .Y(n36) );
  NAND2X0_RVT U119 ( .A1(n34), .A2(n33), .Y(n35) );
  AND2X1_RVT U120 ( .A1(n36), .A2(n35), .Y(m5stg_exp_pre1_in[7]) );
  INVX1_RVT U121 ( .A(n37), .Y(n85) );
  AND2X1_RVT U122 ( .A1(m4stg_exp[8]), .A2(n85), .Y(n78) );
  NAND2X0_RVT U123 ( .A1(m4stg_exp[9]), .A2(n78), .Y(n74) );
  AND2X1_RVT U124 ( .A1(n74), .A2(m6stg_step), .Y(n41) );
  NAND2X0_RVT U125 ( .A1(n39), .A2(n38), .Y(n40) );
  AND2X1_RVT U126 ( .A1(n41), .A2(n40), .Y(m5stg_exp_pre1_in[9]) );
  AO21X1_RVT U127 ( .A1(m5stg_exp_pre1[12]), .A2(n147), .A3(m5stg_exp_pre3[12]), .Y(m5stg_exp[12]) );
  NAND2X0_RVT U129 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[8]), .Y(
        \intadd_5/A[7] ) );
  NAND2X0_RVT U130 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[8]), .Y(
        \intadd_5/B[7] ) );
  NAND2X0_RVT U131 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[9]), .Y(
        \intadd_5/A[8] ) );
  NAND2X0_RVT U132 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[9]), .Y(
        \intadd_5/B[8] ) );
  NAND2X0_RVT U133 ( .A1(m1stg_dblop), .A2(m1stg_exp_in1[10]), .Y(
        \intadd_5/A[9] ) );
  NAND2X0_RVT U134 ( .A1(m1stg_dblop), .A2(m1stg_exp_in2[10]), .Y(
        \intadd_5/B[9] ) );
  INVX1_RVT U135 ( .A(m2stg_exp_expadd), .Y(n44) );
  NOR2X0_RVT U136 ( .A1(m2stg_exp_04ff), .A2(m2stg_exp_0bff), .Y(n42) );
  OAI21X1_RVT U137 ( .A1(\intadd_5/SUM[6] ), .A2(n44), .A3(n42), .Y(
        m2stg_exp_in[7]) );
  INVX1_RVT U138 ( .A(\intadd_5/SUM[8] ), .Y(n43) );
  AO21X1_RVT U139 ( .A1(n43), .A2(m2stg_exp_expadd), .A3(m2stg_exp_0bff), .Y(
        m2stg_exp_in[9]) );
  NOR3X0_RVT U140 ( .A1(m2stg_exp_017f), .A2(m2stg_exp_04ff), .A3(
        m2stg_exp_0bff), .Y(n49) );
  OAI21X1_RVT U141 ( .A1(\intadd_5/SUM[5] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[6]) );
  OAI21X1_RVT U142 ( .A1(\intadd_5/SUM[4] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[5]) );
  OAI21X1_RVT U143 ( .A1(\intadd_5/SUM[3] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[4]) );
  OAI21X1_RVT U144 ( .A1(\intadd_5/SUM[2] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[3]) );
  OAI21X1_RVT U145 ( .A1(\intadd_5/SUM[1] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[2]) );
  OAI21X1_RVT U146 ( .A1(\intadd_5/SUM[0] ), .A2(n44), .A3(n49), .Y(
        m2stg_exp_in[1]) );
  AO221X1_RVT U147 ( .A1(n47), .A2(n46), .A3(n47), .A4(n45), .A5(n44), .Y(n48)
         );
  NAND2X0_RVT U148 ( .A1(n49), .A2(n48), .Y(m2stg_exp_in[0]) );
  OR2X1_RVT U149 ( .A1(m3stg_expa[9]), .A2(n56), .Y(n54) );
  OR2X1_RVT U150 ( .A1(m3stg_expa[10]), .A2(n54), .Y(n52) );
  OR2X1_RVT U151 ( .A1(m3stg_expa[11]), .A2(n52), .Y(n50) );
  XOR2X1_RVT U152 ( .A1(m3stg_expa[12]), .A2(n50), .Y(n151) );
  OA221X1_RVT U153 ( .A1(n51), .A2(m3stg_expa[11]), .A3(n51), .A4(n52), .A5(
        n151), .Y(m4stg_exp_in[11]) );
  OA221X1_RVT U154 ( .A1(n53), .A2(m3stg_expa[10]), .A3(n53), .A4(n54), .A5(
        n151), .Y(m4stg_exp_in[10]) );
  OA221X1_RVT U155 ( .A1(n55), .A2(m3stg_expa[9]), .A3(n55), .A4(n56), .A5(
        n151), .Y(m4stg_exp_in[9]) );
  OR2X1_RVT U156 ( .A1(m3stg_expa[7]), .A2(\intadd_6/n1 ), .Y(n71) );
  OA221X1_RVT U157 ( .A1(n70), .A2(m3stg_expa[8]), .A3(n70), .A4(n71), .A5(
        n151), .Y(m4stg_exp_in[8]) );
  INVX1_RVT U158 ( .A(n71), .Y(n72) );
  OA221X1_RVT U159 ( .A1(n72), .A2(\intadd_6/n1 ), .A3(n72), .A4(m3stg_expa[7]), .A5(n151), .Y(m4stg_exp_in[7]) );
  AND2X1_RVT U160 ( .A1(\intadd_6/SUM[5] ), .A2(n151), .Y(m4stg_exp_in[6]) );
  AND2X1_RVT U161 ( .A1(\intadd_6/SUM[4] ), .A2(n151), .Y(m4stg_exp_in[5]) );
  AND2X1_RVT U162 ( .A1(\intadd_6/SUM[3] ), .A2(n151), .Y(m4stg_exp_in[4]) );
  AND2X1_RVT U163 ( .A1(\intadd_6/SUM[2] ), .A2(n151), .Y(m4stg_exp_in[3]) );
  AND2X1_RVT U164 ( .A1(\intadd_6/SUM[1] ), .A2(n151), .Y(m4stg_exp_in[2]) );
  AND2X1_RVT U165 ( .A1(\intadd_6/SUM[0] ), .A2(n151), .Y(m4stg_exp_in[1]) );
  INVX1_RVT U166 ( .A(\intadd_6/CI ), .Y(n73) );
  OA221X1_RVT U167 ( .A1(n73), .A2(m3stg_ld0_inv[0]), .A3(n73), .A4(
        m3stg_expa[0]), .A5(n151), .Y(m4stg_exp_in[0]) );
  AND2X1_RVT U168 ( .A1(m6stg_step), .A2(m4stg_exp[11]), .Y(
        m5stg_exp_pre2_in[11]) );
  INVX1_RVT U169 ( .A(n74), .Y(n81) );
  NAND2X0_RVT U170 ( .A1(m4stg_exp[10]), .A2(n81), .Y(n75) );
  INVX1_RVT U171 ( .A(n75), .Y(n77) );
  AND2X1_RVT U172 ( .A1(m5stg_exp_pre2_in[11]), .A2(n77), .Y(
        m5stg_exp_pre1_in[12]) );
  OA221X1_RVT U173 ( .A1(m4stg_exp[11]), .A2(n77), .A3(n76), .A4(n75), .A5(
        m6stg_step), .Y(m5stg_exp_pre1_in[11]) );
  AND2X1_RVT U174 ( .A1(m6stg_step), .A2(m4stg_exp[9]), .Y(
        m5stg_exp_pre2_in[9]) );
  NAND2X0_RVT U175 ( .A1(n78), .A2(m5stg_exp_pre2_in[9]), .Y(n79) );
  OAI22X1_RVT U176 ( .A1(n81), .A2(n80), .A3(m4stg_exp[10]), .A4(n79), .Y(
        m5stg_exp_pre1_in[10]) );
  AND2X1_RVT U177 ( .A1(m6stg_step), .A2(m4stg_exp[7]), .Y(
        m5stg_exp_pre2_in[7]) );
  NAND2X0_RVT U178 ( .A1(n82), .A2(m5stg_exp_pre2_in[7]), .Y(n83) );
  OAI22X1_RVT U179 ( .A1(n85), .A2(n84), .A3(m4stg_exp[8]), .A4(n83), .Y(
        m5stg_exp_pre1_in[8]) );
  AND2X1_RVT U180 ( .A1(m6stg_step), .A2(m4stg_exp[5]), .Y(
        m5stg_exp_pre2_in[5]) );
  NAND2X0_RVT U181 ( .A1(n86), .A2(m5stg_exp_pre2_in[5]), .Y(n87) );
  OAI22X1_RVT U182 ( .A1(n89), .A2(n88), .A3(m4stg_exp[6]), .A4(n87), .Y(
        m5stg_exp_pre1_in[6]) );
  AND2X1_RVT U183 ( .A1(m6stg_step), .A2(m4stg_exp[3]), .Y(
        m5stg_exp_pre2_in[3]) );
  NAND4X0_RVT U184 ( .A1(m4stg_exp[2]), .A2(m4stg_exp[0]), .A3(m4stg_exp[1]), 
        .A4(m5stg_exp_pre2_in[3]), .Y(n90) );
  OAI22X1_RVT U185 ( .A1(n92), .A2(n91), .A3(m4stg_exp[4]), .A4(n90), .Y(
        m5stg_exp_pre1_in[4]) );
  AND2X1_RVT U186 ( .A1(m6stg_step), .A2(m4stg_exp[2]), .Y(
        m5stg_exp_pre2_in[2]) );
  AND2X1_RVT U187 ( .A1(m6stg_step), .A2(m4stg_exp[0]), .Y(
        m5stg_exp_pre2_in[0]) );
  NAND2X0_RVT U188 ( .A1(m4stg_exp[0]), .A2(m4stg_exp[1]), .Y(n95) );
  AND2X1_RVT U189 ( .A1(m4stg_exp[1]), .A2(m5stg_exp_pre2_in[0]), .Y(n94) );
  AO22X1_RVT U190 ( .A1(m5stg_exp_pre2_in[2]), .A2(n95), .A3(n94), .A4(n93), 
        .Y(m5stg_exp_pre1_in[2]) );
  AND2X1_RVT U191 ( .A1(m6stg_step), .A2(m4stg_exp[1]), .Y(
        m5stg_exp_pre2_in[1]) );
  INVX1_RVT U192 ( .A(m4stg_exp[0]), .Y(n97) );
  AO22X1_RVT U193 ( .A1(m5stg_exp_pre2_in[0]), .A2(n96), .A3(
        m5stg_exp_pre2_in[1]), .A4(n97), .Y(m5stg_exp_pre1_in[1]) );
  AND2X1_RVT U194 ( .A1(m6stg_step), .A2(n97), .Y(m5stg_exp_pre1_in[0]) );
  NAND2X0_RVT U195 ( .A1(m5stg_in_of), .A2(m5stg_fmuld), .Y(n109) );
  AND3X1_RVT U196 ( .A1(m5stg_exp[2]), .A2(m5stg_exp[0]), .A3(m5stg_exp[1]), 
        .Y(n128) );
  AND3X1_RVT U197 ( .A1(n128), .A2(m5stg_exp[3]), .A3(m5stg_exp[4]), .Y(n120)
         );
  NAND3X0_RVT U198 ( .A1(n120), .A2(m5stg_exp[5]), .A3(m5stg_exp[6]), .Y(n112)
         );
  INVX1_RVT U199 ( .A(n112), .Y(n110) );
  AND3X1_RVT U200 ( .A1(n110), .A2(m5stg_exp[8]), .A3(m5stg_exp[7]), .Y(n98)
         );
  NAND2X0_RVT U201 ( .A1(m5stg_fracadd_cout), .A2(mul_exp_out_exp_plus1), .Y(
        n138) );
  INVX1_RVT U202 ( .A(mul_exp_out_exp), .Y(n111) );
  OA21X1_RVT U203 ( .A1(m5stg_in_of), .A2(m5stg_fracadd_cout), .A3(n111), .Y(
        n142) );
  OA21X1_RVT U204 ( .A1(n98), .A2(n138), .A3(n142), .Y(n102) );
  AO221X1_RVT U205 ( .A1(n102), .A2(n138), .A3(n102), .A4(m5stg_exp[9]), .A5(
        n99), .Y(n101) );
  INVX1_RVT U206 ( .A(n138), .Y(n146) );
  NAND4X0_RVT U207 ( .A1(n146), .A2(n110), .A3(m5stg_exp[7]), .A4(m5stg_exp[8]), .Y(n104) );
  NAND3X0_RVT U208 ( .A1(n109), .A2(n101), .A3(n100), .Y(mul_exp_out_in[10])
         );
  OAI221X1_RVT U209 ( .A1(m5stg_exp[9]), .A2(n104), .A3(n103), .A4(n102), .A5(
        n109), .Y(mul_exp_out_in[9]) );
  AND2X1_RVT U210 ( .A1(n110), .A2(m5stg_exp[7]), .Y(n105) );
  AO221X1_RVT U211 ( .A1(n142), .A2(n105), .A3(n142), .A4(n138), .A5(n106), 
        .Y(n108) );
  NAND4X0_RVT U212 ( .A1(n106), .A2(n146), .A3(n110), .A4(m5stg_exp[7]), .Y(
        n107) );
  NAND3X0_RVT U213 ( .A1(n109), .A2(n108), .A3(n107), .Y(mul_exp_out_in[8]) );
  AND2X1_RVT U214 ( .A1(n146), .A2(n110), .Y(n114) );
  NAND2X0_RVT U215 ( .A1(m5stg_fracadd_cout), .A2(n111), .Y(n116) );
  AO21X1_RVT U216 ( .A1(n146), .A2(n112), .A3(n116), .Y(n113) );
  AO221X1_RVT U217 ( .A1(n115), .A2(n114), .A3(m5stg_exp[7]), .A4(n113), .A5(
        m5stg_in_of), .Y(mul_exp_out_in[7]) );
  INVX1_RVT U218 ( .A(n116), .Y(n133) );
  OA21X1_RVT U219 ( .A1(n120), .A2(n138), .A3(n133), .Y(n121) );
  AO221X1_RVT U220 ( .A1(n121), .A2(m5stg_exp[5]), .A3(n121), .A4(n138), .A5(
        n117), .Y(n119) );
  NAND4X0_RVT U221 ( .A1(n146), .A2(n117), .A3(n120), .A4(m5stg_exp[5]), .Y(
        n118) );
  NAND3X0_RVT U222 ( .A1(n140), .A2(n119), .A3(n118), .Y(mul_exp_out_in[6]) );
  AND2X1_RVT U223 ( .A1(n146), .A2(n120), .Y(n123) );
  INVX1_RVT U224 ( .A(n121), .Y(n122) );
  AO221X1_RVT U225 ( .A1(n124), .A2(n123), .A3(m5stg_exp[5]), .A4(n122), .A5(
        m5stg_in_of), .Y(mul_exp_out_in[5]) );
  OA21X1_RVT U226 ( .A1(n128), .A2(n138), .A3(n133), .Y(n129) );
  AO221X1_RVT U227 ( .A1(n129), .A2(m5stg_exp[3]), .A3(n129), .A4(n138), .A5(
        n125), .Y(n127) );
  NAND4X0_RVT U228 ( .A1(n146), .A2(n125), .A3(n128), .A4(m5stg_exp[3]), .Y(
        n126) );
  NAND3X0_RVT U229 ( .A1(n140), .A2(n127), .A3(n126), .Y(mul_exp_out_in[4]) );
  AND2X1_RVT U230 ( .A1(n146), .A2(n128), .Y(n131) );
  INVX1_RVT U231 ( .A(n129), .Y(n130) );
  AO221X1_RVT U232 ( .A1(n132), .A2(n131), .A3(m5stg_exp[3]), .A4(n130), .A5(
        m5stg_in_of), .Y(mul_exp_out_in[3]) );
  OA21X1_RVT U233 ( .A1(n138), .A2(m5stg_exp[0]), .A3(n133), .Y(n137) );
  AO221X1_RVT U234 ( .A1(n137), .A2(n138), .A3(n137), .A4(m5stg_exp[1]), .A5(
        n134), .Y(n136) );
  NAND4X0_RVT U235 ( .A1(n134), .A2(n146), .A3(m5stg_exp[0]), .A4(m5stg_exp[1]), .Y(n135) );
  NAND3X0_RVT U236 ( .A1(n140), .A2(n136), .A3(n135), .Y(mul_exp_out_in[2]) );
  AO222X1_RVT U237 ( .A1(n139), .A2(n145), .A3(n139), .A4(n138), .A5(n137), 
        .A6(m5stg_exp[1]), .Y(n141) );
  NAND2X0_RVT U238 ( .A1(n141), .A2(n140), .Y(mul_exp_out_in[1]) );
  AO22X1_RVT U239 ( .A1(m5stg_in_of), .A2(m5stg_to_0_inv), .A3(n143), .A4(
        m5stg_exp[0]), .Y(n144) );
  AO21X1_RVT U240 ( .A1(n146), .A2(n145), .A3(n144), .Y(mul_exp_out_in[0]) );
  NAND2X0_RVT U241 ( .A1(n149), .A2(m5stg_exp[12]), .Y(n69) );
  AO221X1_RVT U242 ( .A1(n148), .A2(m5stg_exp_pre2[11]), .A3(n147), .A4(
        m5stg_exp_pre1[11]), .A5(m5stg_exp_pre3[11]), .Y(m5stg_exp[11]) );
  NAND2X0_RVT U243 ( .A1(n149), .A2(m5stg_exp[11]), .Y(n68) );
  NAND2X0_RVT U244 ( .A1(m5stg_exp[10]), .A2(n149), .Y(n67) );
  NAND2X0_RVT U245 ( .A1(m5stg_exp[9]), .A2(n149), .Y(n66) );
  NAND2X0_RVT U246 ( .A1(m5stg_exp[8]), .A2(n149), .Y(n65) );
  NAND2X0_RVT U247 ( .A1(m5stg_exp[7]), .A2(n149), .Y(n64) );
  INVX1_RVT U248 ( .A(m6stg_step), .Y(n149) );
  NAND2X0_RVT U249 ( .A1(m5stg_exp[6]), .A2(n149), .Y(n63) );
  NAND2X0_RVT U250 ( .A1(m5stg_exp[5]), .A2(n149), .Y(n62) );
  NAND2X0_RVT U251 ( .A1(m5stg_exp[4]), .A2(n149), .Y(n61) );
  NAND2X0_RVT U252 ( .A1(m5stg_exp[3]), .A2(n149), .Y(n60) );
  NAND2X0_RVT U253 ( .A1(m5stg_exp[2]), .A2(n149), .Y(n59) );
  NAND2X0_RVT U254 ( .A1(m5stg_exp[1]), .A2(n149), .Y(n58) );
  NAND2X0_RVT U255 ( .A1(m5stg_exp[0]), .A2(n149), .Y(n57) );
  INVX1_RVT U256 ( .A(m3stg_expadd_eq_0), .Y(n150) );
  AND2X1_RVT U257 ( .A1(n151), .A2(n150), .Y(m3stg_expadd_lte_0_inv) );
  OR2X1_RVT U258 ( .A1(m2stg_fmuls), .A2(m2stg_fsmuld), .Y(n155) );
  AO22X1_RVT U259 ( .A1(m2stg_fmuls), .A2(m2stg_exp[7]), .A3(m2stg_exp[8]), 
        .A4(n155), .Y(n154) );
  AOI21X1_RVT U260 ( .A1(m2stg_exp[9]), .A2(n155), .A3(n154), .Y(
        \intadd_7/B[0] ) );
  NAND2X0_RVT U261 ( .A1(m2stg_fmuls), .A2(m2stg_exp[7]), .Y(n152) );
  OA21X1_RVT U262 ( .A1(m2stg_fmuls), .A2(m2stg_exp[7]), .A3(n152), .Y(
        m2stg_expadd[7]) );
  AND2X1_RVT U263 ( .A1(n155), .A2(n152), .Y(n153) );
  HADDX1_RVT U264 ( .A0(n153), .B0(m2stg_exp[8]), .SO(m2stg_expadd[8]) );
  FADDX1_RVT U265 ( .A(m2stg_exp[9]), .B(n155), .CI(n154), .S(m2stg_expadd[9])
         );
endmodule


module fpu_cnt_lead0_lvl4_5 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX1_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_24_eq_0), .A2(n1), .Y(lead0_32b_3) );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl4_6 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_16_eq_0), .A2(din_15_0_eq_0), .Y(din_31_0_eq_0)
         );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(din_15_8_eq_0), .A3(n1), .A4(
        din_31_24_eq_0), .Y(lead0_32b_3) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U6 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl3_7 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_8 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_9 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl1_27 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_28 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_29 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_30 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_31 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_32 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_33 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_34 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_35 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_36 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_37 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_38 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_39 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl2_13 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_14 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_15 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_16 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_17 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_18 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_53b_0 ( din, lead0 );
  input [52:0] din;
  output [5:0] lead0;
  wire   din_52_49_eq_0, din_52_51_eq_0, lead0_52_49_0, din_48_45_eq_0,
         din_48_47_eq_0, lead0_48_45_0, din_44_41_eq_0, din_44_43_eq_0,
         lead0_44_41_0, din_40_37_eq_0, din_40_39_eq_0, lead0_40_37_0,
         din_36_33_eq_0, din_36_35_eq_0, lead0_36_33_0, din_32_29_eq_0,
         din_32_31_eq_0, lead0_32_29_0, din_28_25_eq_0, din_28_27_eq_0,
         lead0_28_25_0, din_24_21_eq_0, din_24_23_eq_0, lead0_24_21_0,
         din_20_17_eq_0, din_20_19_eq_0, lead0_20_17_0, din_16_13_eq_0,
         din_16_15_eq_0, lead0_16_13_0, din_12_9_eq_0, din_12_11_eq_0,
         lead0_12_9_0, din_8_5_eq_0, din_8_7_eq_0, lead0_8_5_0, din_4_1_eq_0,
         din_4_3_eq_0, lead0_4_1_0, din_52_45_eq_0, lead0_52_45_1,
         lead0_52_45_0, din_44_37_eq_0, lead0_44_37_1, lead0_44_37_0,
         din_36_29_eq_0, lead0_36_29_1, lead0_36_29_0, din_28_21_eq_0,
         lead0_28_21_1, lead0_28_21_0, din_20_13_eq_0, lead0_20_13_1,
         lead0_20_13_0, din_12_5_eq_0, lead0_12_5_1, lead0_12_5_0, lead0_4_0_1,
         lead0_4_0_0, din_52_37_eq_0, lead0_52_37_2, lead0_52_37_1,
         lead0_52_37_0, din_36_21_eq_0, lead0_36_21_2, lead0_36_21_1,
         lead0_36_21_0, din_20_5_eq_0, lead0_20_5_2, lead0_20_5_1,
         lead0_20_5_0, lead0_52_21_3, lead0_52_21_2, lead0_52_21_1,
         lead0_52_21_0, lead0_20_0_3, lead0_20_0_2, lead0_20_0_1, lead0_20_0_0,
         n1, n2;

  fpu_cnt_lead0_lvl1_39 i_fpu_cnt_lead0_lvl1_52_49 ( .din(din[52:49]), 
        .din_3_0_eq_0(din_52_49_eq_0), .din_3_2_eq_0(din_52_51_eq_0), 
        .lead0_4b_0(lead0_52_49_0) );
  fpu_cnt_lead0_lvl1_38 i_fpu_cnt_lead0_lvl1_48_45 ( .din(din[48:45]), 
        .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(din_48_47_eq_0), 
        .lead0_4b_0(lead0_48_45_0) );
  fpu_cnt_lead0_lvl1_37 i_fpu_cnt_lead0_lvl1_44_41 ( .din(din[44:41]), 
        .din_3_0_eq_0(din_44_41_eq_0), .din_3_2_eq_0(din_44_43_eq_0), 
        .lead0_4b_0(lead0_44_41_0) );
  fpu_cnt_lead0_lvl1_36 i_fpu_cnt_lead0_lvl1_40_37 ( .din(din[40:37]), 
        .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(din_40_39_eq_0), 
        .lead0_4b_0(lead0_40_37_0) );
  fpu_cnt_lead0_lvl1_35 i_fpu_cnt_lead0_lvl1_36_33 ( .din(din[36:33]), 
        .din_3_0_eq_0(din_36_33_eq_0), .din_3_2_eq_0(din_36_35_eq_0), 
        .lead0_4b_0(lead0_36_33_0) );
  fpu_cnt_lead0_lvl1_34 i_fpu_cnt_lead0_lvl1_32_29 ( .din(din[32:29]), 
        .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(din_32_31_eq_0), 
        .lead0_4b_0(lead0_32_29_0) );
  fpu_cnt_lead0_lvl1_33 i_fpu_cnt_lead0_lvl1_28_25 ( .din(din[28:25]), 
        .din_3_0_eq_0(din_28_25_eq_0), .din_3_2_eq_0(din_28_27_eq_0), 
        .lead0_4b_0(lead0_28_25_0) );
  fpu_cnt_lead0_lvl1_32 i_fpu_cnt_lead0_lvl1_24_21 ( .din(din[24:21]), 
        .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(din_24_23_eq_0), 
        .lead0_4b_0(lead0_24_21_0) );
  fpu_cnt_lead0_lvl1_31 i_fpu_cnt_lead0_lvl1_20_17 ( .din(din[20:17]), 
        .din_3_0_eq_0(din_20_17_eq_0), .din_3_2_eq_0(din_20_19_eq_0), 
        .lead0_4b_0(lead0_20_17_0) );
  fpu_cnt_lead0_lvl1_30 i_fpu_cnt_lead0_lvl1_16_13 ( .din(din[16:13]), 
        .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(din_16_15_eq_0), 
        .lead0_4b_0(lead0_16_13_0) );
  fpu_cnt_lead0_lvl1_29 i_fpu_cnt_lead0_lvl1_12_9 ( .din(din[12:9]), 
        .din_3_0_eq_0(din_12_9_eq_0), .din_3_2_eq_0(din_12_11_eq_0), 
        .lead0_4b_0(lead0_12_9_0) );
  fpu_cnt_lead0_lvl1_28 i_fpu_cnt_lead0_lvl1_8_5 ( .din(din[8:5]), 
        .din_3_0_eq_0(din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0(
        lead0_8_5_0) );
  fpu_cnt_lead0_lvl1_27 i_fpu_cnt_lead0_lvl1_4_1 ( .din(din[4:1]), 
        .din_3_0_eq_0(din_4_1_eq_0), .din_3_2_eq_0(din_4_3_eq_0), .lead0_4b_0(
        lead0_4_1_0) );
  fpu_cnt_lead0_lvl2_18 i_fpu_cnt_lead0_lvl2_52_45 ( .din_7_4_eq_0(
        din_52_49_eq_0), .din_7_6_eq_0(din_52_51_eq_0), .lead0_4b_0_hi(
        lead0_52_49_0), .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(
        din_48_47_eq_0), .lead0_4b_0_lo(lead0_48_45_0), .din_7_0_eq_0(
        din_52_45_eq_0), .lead0_8b_1(lead0_52_45_1), .lead0_8b_0(lead0_52_45_0) );
  fpu_cnt_lead0_lvl2_17 i_fpu_cnt_lead0_lvl2_44_37 ( .din_7_4_eq_0(
        din_44_41_eq_0), .din_7_6_eq_0(din_44_43_eq_0), .lead0_4b_0_hi(
        lead0_44_41_0), .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(
        din_40_39_eq_0), .lead0_4b_0_lo(lead0_40_37_0), .din_7_0_eq_0(
        din_44_37_eq_0), .lead0_8b_1(lead0_44_37_1), .lead0_8b_0(lead0_44_37_0) );
  fpu_cnt_lead0_lvl2_16 i_fpu_cnt_lead0_lvl2_36_29 ( .din_7_4_eq_0(
        din_36_33_eq_0), .din_7_6_eq_0(din_36_35_eq_0), .lead0_4b_0_hi(
        lead0_36_33_0), .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(
        din_32_31_eq_0), .lead0_4b_0_lo(lead0_32_29_0), .din_7_0_eq_0(
        din_36_29_eq_0), .lead0_8b_1(lead0_36_29_1), .lead0_8b_0(lead0_36_29_0) );
  fpu_cnt_lead0_lvl2_15 i_fpu_cnt_lead0_lvl2_28_21 ( .din_7_4_eq_0(
        din_28_25_eq_0), .din_7_6_eq_0(din_28_27_eq_0), .lead0_4b_0_hi(
        lead0_28_25_0), .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(
        din_24_23_eq_0), .lead0_4b_0_lo(lead0_24_21_0), .din_7_0_eq_0(
        din_28_21_eq_0), .lead0_8b_1(lead0_28_21_1), .lead0_8b_0(lead0_28_21_0) );
  fpu_cnt_lead0_lvl2_14 i_fpu_cnt_lead0_lvl2_20_13 ( .din_7_4_eq_0(
        din_20_17_eq_0), .din_7_6_eq_0(din_20_19_eq_0), .lead0_4b_0_hi(
        lead0_20_17_0), .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(
        din_16_15_eq_0), .lead0_4b_0_lo(lead0_16_13_0), .din_7_0_eq_0(
        din_20_13_eq_0), .lead0_8b_1(lead0_20_13_1), .lead0_8b_0(lead0_20_13_0) );
  fpu_cnt_lead0_lvl2_13 i_fpu_cnt_lead0_lvl2_12_5 ( .din_7_4_eq_0(
        din_12_9_eq_0), .din_7_6_eq_0(din_12_11_eq_0), .lead0_4b_0_hi(
        lead0_12_9_0), .din_3_0_eq_0(din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0_lo(lead0_8_5_0), .din_7_0_eq_0(din_12_5_eq_0), .lead0_8b_1(
        lead0_12_5_1), .lead0_8b_0(lead0_12_5_0) );
  fpu_cnt_lead0_lvl3_9 i_fpu_cnt_lead0_lvl3_52_37 ( .din_15_8_eq_0(
        din_52_45_eq_0), .din_15_12_eq_0(din_52_49_eq_0), .lead0_8b_1_hi(
        lead0_52_45_1), .lead0_8b_0_hi(lead0_52_45_0), .din_7_0_eq_0(
        din_44_37_eq_0), .din_7_4_eq_0(din_44_41_eq_0), .lead0_8b_1_lo(
        lead0_44_37_1), .lead0_8b_0_lo(lead0_44_37_0), .din_15_0_eq_0(
        din_52_37_eq_0), .lead0_16b_2(lead0_52_37_2), .lead0_16b_1(
        lead0_52_37_1), .lead0_16b_0(lead0_52_37_0) );
  fpu_cnt_lead0_lvl3_8 i_fpu_cnt_lead0_lvl3_36_21 ( .din_15_8_eq_0(
        din_36_29_eq_0), .din_15_12_eq_0(din_36_33_eq_0), .lead0_8b_1_hi(
        lead0_36_29_1), .lead0_8b_0_hi(lead0_36_29_0), .din_7_0_eq_0(
        din_28_21_eq_0), .din_7_4_eq_0(din_28_25_eq_0), .lead0_8b_1_lo(
        lead0_28_21_1), .lead0_8b_0_lo(lead0_28_21_0), .din_15_0_eq_0(
        din_36_21_eq_0), .lead0_16b_2(lead0_36_21_2), .lead0_16b_1(
        lead0_36_21_1), .lead0_16b_0(lead0_36_21_0) );
  fpu_cnt_lead0_lvl3_7 i_fpu_cnt_lead0_lvl3_20_5 ( .din_15_8_eq_0(
        din_20_13_eq_0), .din_15_12_eq_0(din_20_17_eq_0), .lead0_8b_1_hi(
        lead0_20_13_1), .lead0_8b_0_hi(lead0_20_13_0), .din_7_0_eq_0(
        din_12_5_eq_0), .din_7_4_eq_0(din_12_9_eq_0), .lead0_8b_1_lo(
        lead0_12_5_1), .lead0_8b_0_lo(lead0_12_5_0), .din_15_0_eq_0(
        din_20_5_eq_0), .lead0_16b_2(lead0_20_5_2), .lead0_16b_1(lead0_20_5_1), 
        .lead0_16b_0(lead0_20_5_0) );
  fpu_cnt_lead0_lvl4_6 i_fpu_cnt_lead0_lvl4_52_21 ( .din_31_16_eq_0(
        din_52_37_eq_0), .din_31_24_eq_0(din_52_45_eq_0), .lead0_16b_2_hi(
        lead0_52_37_2), .lead0_16b_1_hi(lead0_52_37_1), .lead0_16b_0_hi(
        lead0_52_37_0), .din_15_0_eq_0(din_36_21_eq_0), .din_15_8_eq_0(
        din_36_29_eq_0), .lead0_16b_2_lo(lead0_36_21_2), .lead0_16b_1_lo(
        lead0_36_21_1), .lead0_16b_0_lo(lead0_36_21_0), .din_31_0_eq_0(
        lead0[5]), .lead0_32b_3(lead0_52_21_3), .lead0_32b_2(lead0_52_21_2), 
        .lead0_32b_1(lead0_52_21_1), .lead0_32b_0(lead0_52_21_0) );
  fpu_cnt_lead0_lvl4_5 i_fpu_cnt_lead0_lvl4_20_0 ( .din_31_16_eq_0(
        din_20_5_eq_0), .din_31_24_eq_0(din_20_13_eq_0), .lead0_16b_2_hi(
        lead0_20_5_2), .lead0_16b_1_hi(lead0_20_5_1), .lead0_16b_0_hi(
        lead0_20_5_0), .din_15_0_eq_0(1'b0), .din_15_8_eq_0(1'b0), 
        .lead0_16b_2_lo(din_4_1_eq_0), .lead0_16b_1_lo(lead0_4_0_1), 
        .lead0_16b_0_lo(lead0_4_0_0), .lead0_32b_3(lead0_20_0_3), 
        .lead0_32b_2(lead0_20_0_2), .lead0_32b_1(lead0_20_0_1), .lead0_32b_0(
        lead0_20_0_0) );
  INVX0_RVT U2 ( .A(din_4_1_eq_0), .Y(n1) );
  OR2X1_RVT U3 ( .A1(din_4_1_eq_0), .A2(lead0_4_1_0), .Y(lead0_4_0_0) );
  AND2X1_RVT U5 ( .A1(din_4_3_eq_0), .A2(n1), .Y(lead0_4_0_1) );
  INVX1_RVT U6 ( .A(lead0[5]), .Y(n2) );
  AO22X1_RVT U7 ( .A1(lead0[5]), .A2(din_20_5_eq_0), .A3(n2), .A4(
        din_52_37_eq_0), .Y(lead0[4]) );
  AO22X1_RVT U8 ( .A1(lead0[5]), .A2(lead0_20_0_3), .A3(n2), .A4(lead0_52_21_3), .Y(lead0[3]) );
  AO22X1_RVT U9 ( .A1(lead0[5]), .A2(lead0_20_0_2), .A3(n2), .A4(lead0_52_21_2), .Y(lead0[2]) );
  AO22X1_RVT U10 ( .A1(lead0[5]), .A2(lead0_20_0_1), .A3(n2), .A4(
        lead0_52_21_1), .Y(lead0[1]) );
  AO22X1_RVT U11 ( .A1(lead0[5]), .A2(lead0_20_0_0), .A3(n2), .A4(
        lead0_52_21_0), .Y(lead0[0]) );
endmodule


module clken_buf_8 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module fpu_cnt_lead0_lvl4_3 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX1_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_24_eq_0), .A2(n1), .Y(lead0_32b_3) );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl4_4 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  AND2X1_RVT U1 ( .A1(din_31_16_eq_0), .A2(din_15_0_eq_0), .Y(din_31_0_eq_0)
         );
  INVX1_RVT U2 ( .A(din_31_16_eq_0), .Y(n1) );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(din_15_8_eq_0), .A3(n1), .A4(
        din_31_24_eq_0), .Y(lead0_32b_3) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U6 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl3_4 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_5 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_6 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl1_14 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_15 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_16 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_17 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_18 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_19 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_20 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_21 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_22 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_23 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_24 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_25 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_26 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl2_7 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_8 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_9 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_10 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_11 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_12 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_53b_2 ( din, lead0 );
  input [52:0] din;
  output [5:0] lead0;
  wire   din_52_49_eq_0, din_52_51_eq_0, lead0_52_49_0, din_48_45_eq_0,
         din_48_47_eq_0, lead0_48_45_0, din_44_41_eq_0, din_44_43_eq_0,
         lead0_44_41_0, din_40_37_eq_0, din_40_39_eq_0, lead0_40_37_0,
         din_36_33_eq_0, din_36_35_eq_0, lead0_36_33_0, din_32_29_eq_0,
         din_32_31_eq_0, lead0_32_29_0, din_28_25_eq_0, din_28_27_eq_0,
         lead0_28_25_0, din_24_21_eq_0, din_24_23_eq_0, lead0_24_21_0,
         din_20_17_eq_0, din_20_19_eq_0, lead0_20_17_0, din_16_13_eq_0,
         din_16_15_eq_0, lead0_16_13_0, din_12_9_eq_0, din_12_11_eq_0,
         lead0_12_9_0, din_8_5_eq_0, din_8_7_eq_0, lead0_8_5_0, din_4_1_eq_0,
         din_4_3_eq_0, lead0_4_1_0, din_52_45_eq_0, lead0_52_45_1,
         lead0_52_45_0, din_44_37_eq_0, lead0_44_37_1, lead0_44_37_0,
         din_36_29_eq_0, lead0_36_29_1, lead0_36_29_0, din_28_21_eq_0,
         lead0_28_21_1, lead0_28_21_0, din_20_13_eq_0, lead0_20_13_1,
         lead0_20_13_0, din_12_5_eq_0, lead0_12_5_1, lead0_12_5_0, lead0_4_0_1,
         lead0_4_0_0, din_52_37_eq_0, lead0_52_37_2, lead0_52_37_1,
         lead0_52_37_0, din_36_21_eq_0, lead0_36_21_2, lead0_36_21_1,
         lead0_36_21_0, din_20_5_eq_0, lead0_20_5_2, lead0_20_5_1,
         lead0_20_5_0, lead0_52_21_3, lead0_52_21_2, lead0_52_21_1,
         lead0_52_21_0, lead0_20_0_3, lead0_20_0_2, lead0_20_0_1, lead0_20_0_0,
         n1, n2;

  fpu_cnt_lead0_lvl1_26 i_fpu_cnt_lead0_lvl1_52_49 ( .din(din[52:49]), 
        .din_3_0_eq_0(din_52_49_eq_0), .din_3_2_eq_0(din_52_51_eq_0), 
        .lead0_4b_0(lead0_52_49_0) );
  fpu_cnt_lead0_lvl1_25 i_fpu_cnt_lead0_lvl1_48_45 ( .din(din[48:45]), 
        .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(din_48_47_eq_0), 
        .lead0_4b_0(lead0_48_45_0) );
  fpu_cnt_lead0_lvl1_24 i_fpu_cnt_lead0_lvl1_44_41 ( .din(din[44:41]), 
        .din_3_0_eq_0(din_44_41_eq_0), .din_3_2_eq_0(din_44_43_eq_0), 
        .lead0_4b_0(lead0_44_41_0) );
  fpu_cnt_lead0_lvl1_23 i_fpu_cnt_lead0_lvl1_40_37 ( .din(din[40:37]), 
        .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(din_40_39_eq_0), 
        .lead0_4b_0(lead0_40_37_0) );
  fpu_cnt_lead0_lvl1_22 i_fpu_cnt_lead0_lvl1_36_33 ( .din(din[36:33]), 
        .din_3_0_eq_0(din_36_33_eq_0), .din_3_2_eq_0(din_36_35_eq_0), 
        .lead0_4b_0(lead0_36_33_0) );
  fpu_cnt_lead0_lvl1_21 i_fpu_cnt_lead0_lvl1_32_29 ( .din(din[32:29]), 
        .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(din_32_31_eq_0), 
        .lead0_4b_0(lead0_32_29_0) );
  fpu_cnt_lead0_lvl1_20 i_fpu_cnt_lead0_lvl1_28_25 ( .din(din[28:25]), 
        .din_3_0_eq_0(din_28_25_eq_0), .din_3_2_eq_0(din_28_27_eq_0), 
        .lead0_4b_0(lead0_28_25_0) );
  fpu_cnt_lead0_lvl1_19 i_fpu_cnt_lead0_lvl1_24_21 ( .din(din[24:21]), 
        .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(din_24_23_eq_0), 
        .lead0_4b_0(lead0_24_21_0) );
  fpu_cnt_lead0_lvl1_18 i_fpu_cnt_lead0_lvl1_20_17 ( .din(din[20:17]), 
        .din_3_0_eq_0(din_20_17_eq_0), .din_3_2_eq_0(din_20_19_eq_0), 
        .lead0_4b_0(lead0_20_17_0) );
  fpu_cnt_lead0_lvl1_17 i_fpu_cnt_lead0_lvl1_16_13 ( .din(din[16:13]), 
        .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(din_16_15_eq_0), 
        .lead0_4b_0(lead0_16_13_0) );
  fpu_cnt_lead0_lvl1_16 i_fpu_cnt_lead0_lvl1_12_9 ( .din(din[12:9]), 
        .din_3_0_eq_0(din_12_9_eq_0), .din_3_2_eq_0(din_12_11_eq_0), 
        .lead0_4b_0(lead0_12_9_0) );
  fpu_cnt_lead0_lvl1_15 i_fpu_cnt_lead0_lvl1_8_5 ( .din(din[8:5]), 
        .din_3_0_eq_0(din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0(
        lead0_8_5_0) );
  fpu_cnt_lead0_lvl1_14 i_fpu_cnt_lead0_lvl1_4_1 ( .din(din[4:1]), 
        .din_3_0_eq_0(din_4_1_eq_0), .din_3_2_eq_0(din_4_3_eq_0), .lead0_4b_0(
        lead0_4_1_0) );
  fpu_cnt_lead0_lvl2_12 i_fpu_cnt_lead0_lvl2_52_45 ( .din_7_4_eq_0(
        din_52_49_eq_0), .din_7_6_eq_0(din_52_51_eq_0), .lead0_4b_0_hi(
        lead0_52_49_0), .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(
        din_48_47_eq_0), .lead0_4b_0_lo(lead0_48_45_0), .din_7_0_eq_0(
        din_52_45_eq_0), .lead0_8b_1(lead0_52_45_1), .lead0_8b_0(lead0_52_45_0) );
  fpu_cnt_lead0_lvl2_11 i_fpu_cnt_lead0_lvl2_44_37 ( .din_7_4_eq_0(
        din_44_41_eq_0), .din_7_6_eq_0(din_44_43_eq_0), .lead0_4b_0_hi(
        lead0_44_41_0), .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(
        din_40_39_eq_0), .lead0_4b_0_lo(lead0_40_37_0), .din_7_0_eq_0(
        din_44_37_eq_0), .lead0_8b_1(lead0_44_37_1), .lead0_8b_0(lead0_44_37_0) );
  fpu_cnt_lead0_lvl2_10 i_fpu_cnt_lead0_lvl2_36_29 ( .din_7_4_eq_0(
        din_36_33_eq_0), .din_7_6_eq_0(din_36_35_eq_0), .lead0_4b_0_hi(
        lead0_36_33_0), .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(
        din_32_31_eq_0), .lead0_4b_0_lo(lead0_32_29_0), .din_7_0_eq_0(
        din_36_29_eq_0), .lead0_8b_1(lead0_36_29_1), .lead0_8b_0(lead0_36_29_0) );
  fpu_cnt_lead0_lvl2_9 i_fpu_cnt_lead0_lvl2_28_21 ( .din_7_4_eq_0(
        din_28_25_eq_0), .din_7_6_eq_0(din_28_27_eq_0), .lead0_4b_0_hi(
        lead0_28_25_0), .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(
        din_24_23_eq_0), .lead0_4b_0_lo(lead0_24_21_0), .din_7_0_eq_0(
        din_28_21_eq_0), .lead0_8b_1(lead0_28_21_1), .lead0_8b_0(lead0_28_21_0) );
  fpu_cnt_lead0_lvl2_8 i_fpu_cnt_lead0_lvl2_20_13 ( .din_7_4_eq_0(
        din_20_17_eq_0), .din_7_6_eq_0(din_20_19_eq_0), .lead0_4b_0_hi(
        lead0_20_17_0), .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(
        din_16_15_eq_0), .lead0_4b_0_lo(lead0_16_13_0), .din_7_0_eq_0(
        din_20_13_eq_0), .lead0_8b_1(lead0_20_13_1), .lead0_8b_0(lead0_20_13_0) );
  fpu_cnt_lead0_lvl2_7 i_fpu_cnt_lead0_lvl2_12_5 ( .din_7_4_eq_0(din_12_9_eq_0), .din_7_6_eq_0(din_12_11_eq_0), .lead0_4b_0_hi(lead0_12_9_0), .din_3_0_eq_0(
        din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0_lo(lead0_8_5_0), .din_7_0_eq_0(din_12_5_eq_0), .lead0_8b_1(lead0_12_5_1), .lead0_8b_0(
        lead0_12_5_0) );
  fpu_cnt_lead0_lvl3_6 i_fpu_cnt_lead0_lvl3_52_37 ( .din_15_8_eq_0(
        din_52_45_eq_0), .din_15_12_eq_0(din_52_49_eq_0), .lead0_8b_1_hi(
        lead0_52_45_1), .lead0_8b_0_hi(lead0_52_45_0), .din_7_0_eq_0(
        din_44_37_eq_0), .din_7_4_eq_0(din_44_41_eq_0), .lead0_8b_1_lo(
        lead0_44_37_1), .lead0_8b_0_lo(lead0_44_37_0), .din_15_0_eq_0(
        din_52_37_eq_0), .lead0_16b_2(lead0_52_37_2), .lead0_16b_1(
        lead0_52_37_1), .lead0_16b_0(lead0_52_37_0) );
  fpu_cnt_lead0_lvl3_5 i_fpu_cnt_lead0_lvl3_36_21 ( .din_15_8_eq_0(
        din_36_29_eq_0), .din_15_12_eq_0(din_36_33_eq_0), .lead0_8b_1_hi(
        lead0_36_29_1), .lead0_8b_0_hi(lead0_36_29_0), .din_7_0_eq_0(
        din_28_21_eq_0), .din_7_4_eq_0(din_28_25_eq_0), .lead0_8b_1_lo(
        lead0_28_21_1), .lead0_8b_0_lo(lead0_28_21_0), .din_15_0_eq_0(
        din_36_21_eq_0), .lead0_16b_2(lead0_36_21_2), .lead0_16b_1(
        lead0_36_21_1), .lead0_16b_0(lead0_36_21_0) );
  fpu_cnt_lead0_lvl3_4 i_fpu_cnt_lead0_lvl3_20_5 ( .din_15_8_eq_0(
        din_20_13_eq_0), .din_15_12_eq_0(din_20_17_eq_0), .lead0_8b_1_hi(
        lead0_20_13_1), .lead0_8b_0_hi(lead0_20_13_0), .din_7_0_eq_0(
        din_12_5_eq_0), .din_7_4_eq_0(din_12_9_eq_0), .lead0_8b_1_lo(
        lead0_12_5_1), .lead0_8b_0_lo(lead0_12_5_0), .din_15_0_eq_0(
        din_20_5_eq_0), .lead0_16b_2(lead0_20_5_2), .lead0_16b_1(lead0_20_5_1), 
        .lead0_16b_0(lead0_20_5_0) );
  fpu_cnt_lead0_lvl4_4 i_fpu_cnt_lead0_lvl4_52_21 ( .din_31_16_eq_0(
        din_52_37_eq_0), .din_31_24_eq_0(din_52_45_eq_0), .lead0_16b_2_hi(
        lead0_52_37_2), .lead0_16b_1_hi(lead0_52_37_1), .lead0_16b_0_hi(
        lead0_52_37_0), .din_15_0_eq_0(din_36_21_eq_0), .din_15_8_eq_0(
        din_36_29_eq_0), .lead0_16b_2_lo(lead0_36_21_2), .lead0_16b_1_lo(
        lead0_36_21_1), .lead0_16b_0_lo(lead0_36_21_0), .din_31_0_eq_0(
        lead0[5]), .lead0_32b_3(lead0_52_21_3), .lead0_32b_2(lead0_52_21_2), 
        .lead0_32b_1(lead0_52_21_1), .lead0_32b_0(lead0_52_21_0) );
  fpu_cnt_lead0_lvl4_3 i_fpu_cnt_lead0_lvl4_20_0 ( .din_31_16_eq_0(
        din_20_5_eq_0), .din_31_24_eq_0(din_20_13_eq_0), .lead0_16b_2_hi(
        lead0_20_5_2), .lead0_16b_1_hi(lead0_20_5_1), .lead0_16b_0_hi(
        lead0_20_5_0), .din_15_0_eq_0(1'b0), .din_15_8_eq_0(1'b0), 
        .lead0_16b_2_lo(din_4_1_eq_0), .lead0_16b_1_lo(lead0_4_0_1), 
        .lead0_16b_0_lo(lead0_4_0_0), .lead0_32b_3(lead0_20_0_3), 
        .lead0_32b_2(lead0_20_0_2), .lead0_32b_1(lead0_20_0_1), .lead0_32b_0(
        lead0_20_0_0) );
  INVX0_RVT U2 ( .A(din_4_1_eq_0), .Y(n1) );
  OR2X1_RVT U3 ( .A1(din_4_1_eq_0), .A2(lead0_4_1_0), .Y(lead0_4_0_0) );
  AND2X1_RVT U5 ( .A1(din_4_3_eq_0), .A2(n1), .Y(lead0_4_0_1) );
  INVX1_RVT U6 ( .A(lead0[5]), .Y(n2) );
  AO22X1_RVT U7 ( .A1(lead0[5]), .A2(din_20_5_eq_0), .A3(n2), .A4(
        din_52_37_eq_0), .Y(lead0[4]) );
  AO22X1_RVT U8 ( .A1(lead0[5]), .A2(lead0_20_0_3), .A3(n2), .A4(lead0_52_21_3), .Y(lead0[3]) );
  AO22X1_RVT U9 ( .A1(lead0[5]), .A2(lead0_20_0_2), .A3(n2), .A4(lead0_52_21_2), .Y(lead0[2]) );
  AO22X1_RVT U10 ( .A1(lead0[5]), .A2(lead0_20_0_1), .A3(n2), .A4(
        lead0_52_21_1), .Y(lead0[1]) );
  AO22X1_RVT U11 ( .A1(lead0[5]), .A2(lead0_20_0_0), .A3(n2), .A4(
        lead0_52_21_0), .Y(lead0[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_9 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_9 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_8 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_8 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE56 ( din, en, clk, q, se, si, so );
  input [55:0] din;
  output [55:0] q;
  input [55:0] si;
  output [55:0] so;
  input en, clk, se;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         net24354, n3, n1;
  assign q[50] = q[43];

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE56 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24354), .TE(1'b0) );
  DFFX1_RVT \q_reg[50]  ( .D(N47), .CLK(net24354), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24354), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24354), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24354), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24354), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24354), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24354), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24354), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24354), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24354), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24354), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24354), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24354), .Q(q[31]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[31]), .A2(n1), .Y(N35) );
  AND2X1_RVT U4 ( .A1(din[32]), .A2(n1), .Y(N36) );
  AND2X1_RVT U5 ( .A1(din[33]), .A2(n1), .Y(N37) );
  AND2X1_RVT U6 ( .A1(din[34]), .A2(n1), .Y(N38) );
  AND2X1_RVT U7 ( .A1(din[35]), .A2(n1), .Y(N39) );
  AND2X1_RVT U8 ( .A1(din[36]), .A2(n1), .Y(N40) );
  AND2X1_RVT U9 ( .A1(din[37]), .A2(n1), .Y(N41) );
  AND2X1_RVT U10 ( .A1(din[38]), .A2(n1), .Y(N42) );
  AND2X1_RVT U11 ( .A1(din[39]), .A2(n1), .Y(N43) );
  AND2X1_RVT U12 ( .A1(din[40]), .A2(n1), .Y(N44) );
  AND2X1_RVT U13 ( .A1(din[41]), .A2(n1), .Y(N45) );
  AND2X1_RVT U14 ( .A1(din[42]), .A2(n1), .Y(N46) );
  AND2X1_RVT U15 ( .A1(din[43]), .A2(n1), .Y(N47) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module dff_SIZE55_0 ( din, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, n1, n2,
         n3, n4;

  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n3), .Y(N57) );
endmodule


module dff_SIZE55_3 ( din, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, n1, n2, n3, n4
;

  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n1), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  INVX1_RVT U4 ( .A(se), .Y(n2) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n2), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n2), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n2), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n2), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n2), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n2), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n2), .Y(N10) );
  INVX1_RVT U12 ( .A(se), .Y(n3) );
  AND2X1_RVT U13 ( .A1(din[8]), .A2(n3), .Y(N11) );
  AND2X1_RVT U14 ( .A1(din[9]), .A2(n3), .Y(N12) );
  AND2X1_RVT U15 ( .A1(din[10]), .A2(n3), .Y(N13) );
  AND2X1_RVT U16 ( .A1(din[11]), .A2(n3), .Y(N14) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n3), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n3), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n3), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n3), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n3), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n3), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n3), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n3), .Y(N22) );
  INVX1_RVT U25 ( .A(se), .Y(n4) );
  AND2X1_RVT U26 ( .A1(din[20]), .A2(n4), .Y(N23) );
  AND2X1_RVT U27 ( .A1(din[21]), .A2(n4), .Y(N24) );
  AND2X1_RVT U28 ( .A1(din[22]), .A2(n4), .Y(N25) );
  AND2X1_RVT U29 ( .A1(din[23]), .A2(n4), .Y(N26) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n4), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n4), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n4), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n4), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n4), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n4), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n4), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n4), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n2), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n2), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n2), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n2), .Y(N38) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n2), .Y(N39) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n2), .Y(N40) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n3), .Y(N41) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n2), .Y(N44) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n3), .Y(N45) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n1), .Y(N57) );
endmodule


module dff_SIZE55_2 ( din, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, n1, n2,
         n3, n4;

  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n2), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n3), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U60 ( .A1(din[53]), .A2(n2), .Y(N56) );
  AND2X1_RVT U61 ( .A1(din[54]), .A2(n3), .Y(N57) );
endmodule


module dff_SIZE55_1 ( din, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, n1, n2, n3, n4
;

  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n1), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  INVX1_RVT U4 ( .A(se), .Y(n2) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n2), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n2), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n2), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n2), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n2), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n2), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n2), .Y(N10) );
  INVX1_RVT U12 ( .A(se), .Y(n3) );
  AND2X1_RVT U13 ( .A1(din[8]), .A2(n3), .Y(N11) );
  AND2X1_RVT U14 ( .A1(din[9]), .A2(n3), .Y(N12) );
  AND2X1_RVT U15 ( .A1(din[10]), .A2(n3), .Y(N13) );
  AND2X1_RVT U16 ( .A1(din[11]), .A2(n3), .Y(N14) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n3), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n3), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n3), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n3), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n3), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n3), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n3), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n3), .Y(N22) );
  INVX1_RVT U25 ( .A(se), .Y(n4) );
  AND2X1_RVT U26 ( .A1(din[20]), .A2(n4), .Y(N23) );
  AND2X1_RVT U27 ( .A1(din[21]), .A2(n4), .Y(N24) );
  AND2X1_RVT U28 ( .A1(din[22]), .A2(n4), .Y(N25) );
  AND2X1_RVT U29 ( .A1(din[23]), .A2(n4), .Y(N26) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n4), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n4), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n4), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n4), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n4), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n4), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n4), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n4), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n2), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n2), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n2), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n2), .Y(N38) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n2), .Y(N39) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n2), .Y(N40) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n3), .Y(N41) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n2), .Y(N44) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n3), .Y(N45) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n1), .Y(N57) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE52 ( din, en, clk, q, se, si, so );
  input [51:0] din;
  output [51:0] q;
  input [51:0] si;
  output [51:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, net24336, n3, n1, n2, n4,
         n5;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE52 clk_gate_q_reg ( .CLK(clk), .EN(n3), 
        .ENCLK(net24336), .TE(1'b0) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24336), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24336), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24336), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24336), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24336), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24336), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24336), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24336), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24336), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24336), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24336), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24336), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24336), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24336), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24336), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24336), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24336), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24336), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24336), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24336), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24336), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24336), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24336), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24336), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24336), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24336), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24336), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24336), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24336), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24336), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24336), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24336), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24336), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24336), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24336), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24336), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24336), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24336), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24336), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24336), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24336), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24336), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24336), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24336), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24336), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24336), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24336), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24336), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24336), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24336), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24336), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24336), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  OR2X1_RVT U59 ( .A1(se), .A2(en), .Y(n3) );
endmodule


module fpu_mul_frac_dp ( inq_in1, inq_in2, m6stg_step, m2stg_frac1_dbl_norm, 
        m2stg_frac1_dbl_dnrm, m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, 
        m2stg_frac1_inf, m1stg_snan_dbl_in1, m1stg_snan_sng_in1, 
        m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, 
        m2stg_frac2_sng_dnrm, m2stg_frac2_inf, m1stg_snan_dbl_in2, 
        m1stg_snan_sng_in2, m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, 
        m1stg_dblop, m1stg_dblop_inv, m4stg_frac, m4stg_sh_cnt_in, 
        m3bstg_ld0_inv, m4stg_left_shift_step, m4stg_right_shift_step, 
        m5stg_fmuls, m5stg_fmulda, mul_frac_out_fracadd, mul_frac_out_frac, 
        m5stg_in_of, m5stg_to_0, fmul_clken_l, rclk, m2stg_frac1_array_in, 
        m2stg_frac2_array_in, m1stg_ld0_1, m1stg_ld0_2, m4stg_frac_105, 
        m3stg_ld0_inv, m4stg_shl_54, m4stg_shl_55, m5stg_frac_32_0, 
        m5stg_frac_dbl_nx, m5stg_frac_sng_nx, m5stg_frac_neq_0, 
        m5stg_fracadd_cout, mul_frac_out, se, si, so );
  input [54:0] inq_in1;
  input [54:0] inq_in2;
  input [105:0] m4stg_frac;
  input [5:0] m4stg_sh_cnt_in;
  input [6:0] m3bstg_ld0_inv;
  output [52:0] m2stg_frac1_array_in;
  output [52:0] m2stg_frac2_array_in;
  output [5:0] m1stg_ld0_1;
  output [5:0] m1stg_ld0_2;
  output [6:0] m3stg_ld0_inv;
  output [32:0] m5stg_frac_32_0;
  output [51:0] mul_frac_out;
  input m6stg_step, m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm,
         m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, m2stg_frac1_inf,
         m1stg_snan_dbl_in1, m1stg_snan_sng_in1, m2stg_frac2_dbl_norm,
         m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, m2stg_frac2_sng_dnrm,
         m2stg_frac2_inf, m1stg_snan_dbl_in2, m1stg_snan_sng_in2,
         m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, m1stg_dblop,
         m1stg_dblop_inv, m4stg_left_shift_step, m4stg_right_shift_step,
         m5stg_fmuls, m5stg_fmulda, mul_frac_out_fracadd, mul_frac_out_frac,
         m5stg_in_of, m5stg_to_0, fmul_clken_l, rclk, se, si;
  output m4stg_frac_105, m4stg_shl_54, m4stg_shl_55, m5stg_frac_dbl_nx,
         m5stg_frac_sng_nx, m5stg_frac_neq_0, m5stg_fracadd_cout, so;
  wire   clk, \m4stg_sh_cnt_5[0] , n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, \add_x_3/A[29] , \add_x_3/A[28] , \add_x_3/A[27] ,
         \add_x_3/A[26] , \add_x_3/A[25] , \add_x_3/A[24] , \add_x_3/A[23] ,
         \add_x_3/A[22] , \add_x_3/A[21] , \add_x_3/A[20] , \add_x_3/A[19] ,
         \add_x_3/A[18] , \add_x_3/A[15] , \add_x_3/A[14] , \add_x_3/A[13] ,
         \add_x_3/A[12] , \add_x_3/A[11] , \add_x_3/A[10] , \add_x_3/A[9] ,
         \add_x_3/A[8] , \add_x_3/A[7] , \add_x_3/A[6] , \add_x_3/A[5] ,
         \add_x_3/A[4] , \add_x_3/A[3] , \add_x_3/A[2] , \add_x_3/A[1] ,
         \add_x_3/A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
  wire   [54:0] mul_frac_in1;
  wire   [54:0] mul_frac_in2;
  wire   [52:1] m1stg_ld0_1_din;
  wire   [52:1] m1stg_ld0_2_din;
  wire   [5:0] m4stg_sh_cnt;
  wire   [54:0] m5stg_frac_pre1;
  wire   [54:0] m5stg_frac_pre2;
  wire   [54:0] m5stg_frac_pre3;
  wire   [54:0] m5stg_frac_pre4;
  wire   [51:0] mul_frac_out_in;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41;
  assign m4stg_frac_105 = m4stg_frac[105];
  assign m5stg_frac_32_0[32] = \add_x_3/A[29] ;
  assign m5stg_frac_32_0[31] = \add_x_3/A[28] ;
  assign m5stg_frac_32_0[30] = \add_x_3/A[27] ;
  assign m5stg_frac_32_0[29] = \add_x_3/A[26] ;
  assign m5stg_frac_32_0[28] = \add_x_3/A[25] ;
  assign m5stg_frac_32_0[27] = \add_x_3/A[24] ;
  assign m5stg_frac_32_0[26] = \add_x_3/A[23] ;
  assign m5stg_frac_32_0[25] = \add_x_3/A[22] ;
  assign m5stg_frac_32_0[24] = \add_x_3/A[21] ;
  assign m5stg_frac_32_0[23] = \add_x_3/A[20] ;
  assign m5stg_frac_32_0[22] = \add_x_3/A[19] ;
  assign m5stg_frac_32_0[21] = \add_x_3/A[18] ;
  assign m5stg_frac_32_0[18] = \add_x_3/A[15] ;
  assign m5stg_frac_32_0[17] = \add_x_3/A[14] ;
  assign m5stg_frac_32_0[16] = \add_x_3/A[13] ;
  assign m5stg_frac_32_0[15] = \add_x_3/A[12] ;
  assign m5stg_frac_32_0[14] = \add_x_3/A[11] ;
  assign m5stg_frac_32_0[13] = \add_x_3/A[10] ;
  assign m5stg_frac_32_0[12] = \add_x_3/A[9] ;
  assign m5stg_frac_32_0[11] = \add_x_3/A[8] ;
  assign m5stg_frac_32_0[10] = \add_x_3/A[7] ;
  assign m5stg_frac_32_0[9] = \add_x_3/A[6] ;
  assign m5stg_frac_32_0[8] = \add_x_3/A[5] ;
  assign m5stg_frac_32_0[7] = \add_x_3/A[4] ;
  assign m5stg_frac_32_0[6] = \add_x_3/A[3] ;
  assign m5stg_frac_32_0[5] = \add_x_3/A[2] ;
  assign m5stg_frac_32_0[4] = \add_x_3/A[1] ;
  assign m5stg_frac_32_0[3] = \add_x_3/A[0] ;
  assign so = 1'b0;

  clken_buf_8 ckbuf_mul_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fmul_clken_l), 
        .tmb_l(n2148) );
  dffe_SIZE55_9 i_mul_frac_in1 ( .din(inq_in1), .en(m6stg_step), .clk(clk), 
        .q(mul_frac_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE55_8 i_mul_frac_in2 ( .din(inq_in2), .en(m6stg_step), .clk(clk), 
        .q(mul_frac_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  fpu_cnt_lead0_53b_0 i_m1stg_ld0_1 ( .din({m1stg_ld0_1_din, 1'b0}), .lead0(
        m1stg_ld0_1) );
  fpu_cnt_lead0_53b_2 i_m1stg_ld0_2 ( .din({m1stg_ld0_2_din, 1'b0}), .lead0(
        m1stg_ld0_2) );
  dffe_SIZE56 i_mstg_xtra_regs ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        m4stg_sh_cnt_in[5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        m4stg_sh_cnt_in, m3bstg_ld0_inv, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .en(m6stg_step), .clk(clk), .q({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, \m4stg_sh_cnt_5[0] , 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, m4stg_sh_cnt, 
        m3stg_ld0_inv, SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE55_0 i_m5stg_frac_pre1 ( .din({n1878, n1877, n1876, n1875, n1874, 
        n1873, n1872, n1871, n1870, n1869, n1868, n1867, n1866, n1865, n1864, 
        n1863, n1862, n1861, n1860, n1859, n1858, n1857, n1856, n1855, n1854, 
        n1853, n1852, n1851, n1850, n1849, n1848, n1847, n1846, n1845, n1844, 
        n1843, n1842, n1841, n1840, n1839, n1838, n1837, n1836, n1835, n1834, 
        n1833, n1832, n1831, n1830, n1829, n1828, n1827, n1826, n1825, n1824}), 
        .clk(clk), .q(m5stg_frac_pre1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE55_3 i_m5stg_frac_pre2 ( .din({n1770, n1771, n1772, n1773, n1774, 
        n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
        n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
        n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
        n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
        n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 1'b1}), 
        .clk(clk), .q(m5stg_frac_pre2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE55_2 i_m5stg_frac_pre3 ( .din({n1769, n1768, n1767, n1766, n1765, 
        n1764, n1763, n1762, n1761, n1760, n1759, n1758, n1757, n1756, n1755, 
        n1754, n1753, n1752, n1751, n1750, n1749, n1748, n1747, n1746, n1745, 
        n1744, n1743, n1742, n1741, n1740, n1739, n1738, n1737, n1736, n1735, 
        n1734, n1733, n1732, n1731, n1730, n1729, n1728, n1727, n1726, n1725, 
        n1724, n1723, n1722, n1721, n1720, n1719, n1718, n1717, n1716, n1715}), 
        .clk(clk), .q(m5stg_frac_pre3), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dff_SIZE55_1 i_m5stg_frac_pre4 ( .din({n1661, n1662, n1663, n1664, n1665, 
        n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
        n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
        n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
        n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
        n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 1'b1}), 
        .clk(clk), .q(m5stg_frac_pre4), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE52 i_mul_frac_out ( .din(mul_frac_out_in), .en(m6stg_step), .clk(
        clk), .q(mul_frac_out), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  INVX0_RVT U3 ( .A(n661), .Y(n664) );
  INVX0_RVT U4 ( .A(n679), .Y(n676) );
  INVX0_RVT U5 ( .A(n1933), .Y(n1943) );
  INVX0_RVT U6 ( .A(m4stg_shl_55), .Y(n1974) );
  INVX0_RVT U7 ( .A(n1955), .Y(n1287) );
  INVX0_RVT U8 ( .A(n1954), .Y(n1309) );
  INVX0_RVT U9 ( .A(n1961), .Y(n1333) );
  INVX0_RVT U10 ( .A(n421), .Y(n383) );
  INVX0_RVT U11 ( .A(n2073), .Y(n408) );
  OR3X1_RVT U12 ( .A1(n393), .A2(n392), .A3(n391), .Y(n400) );
  INVX0_RVT U13 ( .A(n1469), .Y(n1630) );
  INVX0_RVT U14 ( .A(n1442), .Y(n1615) );
  INVX0_RVT U15 ( .A(n381), .Y(n288) );
  INVX0_RVT U16 ( .A(n1940), .Y(n1586) );
  INVX0_RVT U17 ( .A(n2076), .Y(n449) );
  INVX0_RVT U18 ( .A(n1941), .Y(n1567) );
  INVX0_RVT U19 ( .A(n1944), .Y(n1660) );
  INVX0_RVT U20 ( .A(n390), .Y(n108) );
  OR3X1_RVT U21 ( .A1(n333), .A2(n332), .A3(n331), .Y(n389) );
  INVX0_RVT U22 ( .A(n1901), .Y(n1572) );
  INVX0_RVT U23 ( .A(n1887), .Y(n1634) );
  INVX0_RVT U24 ( .A(n1429), .Y(n1430) );
  INVX0_RVT U25 ( .A(n177), .Y(n157) );
  INVX0_RVT U26 ( .A(n1509), .Y(n1412) );
  INVX0_RVT U27 ( .A(n273), .Y(n277) );
  INVX0_RVT U28 ( .A(n1617), .Y(n1583) );
  INVX0_RVT U29 ( .A(n194), .Y(n143) );
  INVX0_RVT U30 ( .A(n1218), .Y(n1220) );
  INVX0_RVT U31 ( .A(n1175), .Y(n1075) );
  INVX0_RVT U32 ( .A(n1217), .Y(n1222) );
  INVX0_RVT U33 ( .A(n351), .Y(n310) );
  INVX0_RVT U34 ( .A(n1602), .Y(n1564) );
  INVX0_RVT U35 ( .A(n305), .Y(n231) );
  INVX0_RVT U36 ( .A(n290), .Y(n309) );
  INVX0_RVT U37 ( .A(n262), .Y(n276) );
  INVX0_RVT U38 ( .A(n340), .Y(n320) );
  INVX0_RVT U39 ( .A(n360), .Y(n285) );
  INVX0_RVT U40 ( .A(n203), .Y(n132) );
  INVX0_RVT U41 ( .A(n1325), .Y(n1191) );
  INVX0_RVT U42 ( .A(n186), .Y(n151) );
  INVX0_RVT U43 ( .A(n417), .Y(n172) );
  INVX0_RVT U44 ( .A(n1302), .Y(n1132) );
  INVX0_RVT U45 ( .A(n1109), .Y(n1214) );
  INVX0_RVT U46 ( .A(n1111), .Y(n1216) );
  INVX0_RVT U47 ( .A(n1068), .Y(n1167) );
  INVX0_RVT U48 ( .A(n1046), .Y(n1126) );
  INVX0_RVT U49 ( .A(n178), .Y(n138) );
  OR3X1_RVT U50 ( .A1(n412), .A2(n359), .A3(n350), .Y(n339) );
  INVX0_RVT U51 ( .A(n195), .Y(n114) );
  INVX0_RVT U52 ( .A(n291), .Y(n280) );
  INVX0_RVT U53 ( .A(n198), .Y(n162) );
  INVX0_RVT U54 ( .A(n298), .Y(n239) );
  INVX0_RVT U55 ( .A(n418), .Y(n292) );
  INVX0_RVT U56 ( .A(n1388), .Y(n1435) );
  INVX0_RVT U57 ( .A(n295), .Y(n249) );
  INVX0_RVT U58 ( .A(n1400), .Y(n1355) );
  INVX0_RVT U59 ( .A(n181), .Y(n169) );
  INVX0_RVT U60 ( .A(n1378), .Y(n1330) );
  INVX0_RVT U61 ( .A(n1897), .Y(n1900) );
  INVX1_RVT U62 ( .A(n70), .Y(n154) );
  INVX0_RVT U63 ( .A(n1004), .Y(n1005) );
  INVX0_RVT U64 ( .A(n1899), .Y(n1885) );
  INVX0_RVT U65 ( .A(n437), .Y(n2087) );
  INVX0_RVT U66 ( .A(n621), .Y(n1246) );
  INVX0_RVT U67 ( .A(n591), .Y(n1086) );
  INVX0_RVT U68 ( .A(n641), .Y(n1298) );
  INVX0_RVT U69 ( .A(\add_x_3/A[15] ), .Y(n1515) );
  INVX0_RVT U70 ( .A(\add_x_3/A[14] ), .Y(n1526) );
  INVX0_RVT U71 ( .A(\add_x_3/A[21] ), .Y(n1440) );
  INVX0_RVT U72 ( .A(\add_x_3/A[20] ), .Y(n1456) );
  INVX0_RVT U73 ( .A(\add_x_3/A[19] ), .Y(n1467) );
  INVX0_RVT U74 ( .A(\add_x_3/A[18] ), .Y(n1484) );
  INVX0_RVT U75 ( .A(\add_x_3/A[24] ), .Y(n1405) );
  INVX0_RVT U76 ( .A(\add_x_3/A[25] ), .Y(n1392) );
  INVX0_RVT U77 ( .A(n836), .Y(n553) );
  INVX0_RVT U78 ( .A(\add_x_3/A[26] ), .Y(n1383) );
  INVX0_RVT U79 ( .A(\add_x_3/A[13] ), .Y(n1536) );
  INVX0_RVT U80 ( .A(\add_x_3/A[12] ), .Y(n1548) );
  INVX0_RVT U81 ( .A(\add_x_3/A[27] ), .Y(n1370) );
  INVX0_RVT U82 ( .A(n631), .Y(n1276) );
  INVX0_RVT U83 ( .A(\add_x_3/A[28] ), .Y(n1361) );
  INVX0_RVT U84 ( .A(\add_x_3/A[0] ), .Y(n1644) );
  INVX0_RVT U85 ( .A(m5stg_frac_32_0[20]), .Y(n1492) );
  INVX0_RVT U86 ( .A(n636), .Y(n1290) );
  INVX0_RVT U87 ( .A(n566), .Y(n996) );
  INVX0_RVT U88 ( .A(n650), .Y(n1321) );
  INVX0_RVT U89 ( .A(n611), .Y(n1183) );
  INVX0_RVT U90 ( .A(n561), .Y(n982) );
  INVX0_RVT U91 ( .A(n606), .Y(n1153) );
  INVX0_RVT U92 ( .A(\add_x_3/A[29] ), .Y(n1346) );
  INVX0_RVT U93 ( .A(n601), .Y(n1124) );
  INVX0_RVT U94 ( .A(n555), .Y(n913) );
  INVX0_RVT U95 ( .A(n596), .Y(n1108) );
  INVX0_RVT U96 ( .A(n646), .Y(n1312) );
  INVX0_RVT U97 ( .A(n586), .Y(n1064) );
  INVX0_RVT U98 ( .A(n626), .Y(n1261) );
  INVX0_RVT U99 ( .A(n581), .Y(n1044) );
  INVX0_RVT U100 ( .A(n571), .Y(n1013) );
  INVX0_RVT U101 ( .A(n655), .Y(n1336) );
  INVX0_RVT U102 ( .A(n616), .Y(n1212) );
  INVX0_RVT U103 ( .A(n576), .Y(n1028) );
  INVX0_RVT U104 ( .A(\add_x_3/A[23] ), .Y(n1420) );
  INVX0_RVT U105 ( .A(\add_x_3/A[22] ), .Y(n1431) );
  INVX0_RVT U106 ( .A(m5stg_frac_32_0[2]), .Y(n1649) );
  INVX0_RVT U107 ( .A(m5stg_frac_32_0[1]), .Y(n1653) );
  INVX0_RVT U108 ( .A(m4stg_frac[97]), .Y(n843) );
  INVX0_RVT U109 ( .A(m4stg_frac[98]), .Y(n841) );
  INVX0_RVT U110 ( .A(m6stg_step), .Y(n1972) );
  AOI22X1_RVT U111 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[32]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[29]), .Y(n1) );
  AOI22X1_RVT U112 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[33]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[30]), .Y(n2) );
  AOI22X1_RVT U113 ( .A1(m2stg_frac2_inf), .A2(m1stg_inf_zero_in), .A3(
        mul_frac_in2[50]), .A4(m2stg_frac2_dbl_norm), .Y(n3) );
  AOI22X1_RVT U114 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[50]), .A3(
        m2stg_frac2_sng_norm), .A4(n503), .Y(n4) );
  NAND2X0_RVT U115 ( .A1(m5stg_to_0), .A2(m5stg_in_of), .Y(n5) );
  AND2X1_RVT U116 ( .A1(m4stg_sh_cnt[2]), .A2(m4stg_sh_cnt[3]), .Y(n6) );
  AOI22X1_RVT U117 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[29]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n7) );
  AOI221X1_RVT U118 ( .A1(m4stg_sh_cnt[5]), .A2(n2070), .A3(m4stg_sh_cnt[5]), 
        .A4(n441), .A5(n440), .Y(n8) );
  NAND2X0_RVT U119 ( .A1(m2stg_frac2_inf), .A2(m1stg_inf_zero_in), .Y(n9) );
  AOI22X1_RVT U120 ( .A1(m4stg_sh_cnt[5]), .A2(n431), .A3(n430), .A4(n429), 
        .Y(n10) );
  AOI22X1_RVT U121 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[34]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n11) );
  AOI22X1_RVT U122 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[35]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n12) );
  AOI22X1_RVT U123 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[36]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n13) );
  AOI22X1_RVT U124 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[37]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n14) );
  AOI22X1_RVT U125 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[38]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n15) );
  AOI22X1_RVT U126 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[39]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n16) );
  AOI22X1_RVT U127 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[40]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n17) );
  AOI22X1_RVT U128 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[41]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n18) );
  AOI22X1_RVT U129 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[42]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n19) );
  AOI22X1_RVT U130 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[43]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n20) );
  AOI22X1_RVT U131 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[44]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n21) );
  AOI22X1_RVT U132 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[45]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n22) );
  AOI22X1_RVT U133 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[46]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n23) );
  AOI22X1_RVT U134 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[47]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n24) );
  AOI22X1_RVT U135 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[48]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n25) );
  AOI22X1_RVT U136 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[50]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n26) );
  AOI22X1_RVT U137 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[51]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n27) );
  AOI22X1_RVT U138 ( .A1(m2stg_frac2_sng_norm), .A2(mul_frac_in2[52]), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n28) );
  AOI22X1_RVT U139 ( .A1(mul_frac_in2[53]), .A2(m2stg_frac2_sng_norm), .A3(
        mul_frac_in2[52]), .A4(m2stg_frac2_sng_dnrm), .Y(n29) );
  INVX1_RVT U140 ( .A(m4stg_sh_cnt[1]), .Y(n975) );
  NAND2X0_RVT U141 ( .A1(m4stg_sh_cnt[0]), .A2(n975), .Y(n842) );
  INVX1_RVT U142 ( .A(n842), .Y(n1579) );
  INVX1_RVT U143 ( .A(m4stg_sh_cnt[0]), .Y(n778) );
  NAND2X0_RVT U144 ( .A1(n975), .A2(n778), .Y(n772) );
  INVX1_RVT U145 ( .A(n772), .Y(n1593) );
  AO22X1_RVT U146 ( .A1(n1579), .A2(m4stg_frac[44]), .A3(n1593), .A4(
        m4stg_frac[45]), .Y(n31) );
  NAND2X0_RVT U147 ( .A1(m4stg_sh_cnt[1]), .A2(n778), .Y(n844) );
  INVX1_RVT U148 ( .A(n844), .Y(n1573) );
  NAND2X0_RVT U149 ( .A1(m4stg_sh_cnt[1]), .A2(m4stg_sh_cnt[0]), .Y(n779) );
  INVX1_RVT U150 ( .A(n779), .Y(n1422) );
  AO22X1_RVT U151 ( .A1(n1573), .A2(m4stg_frac[43]), .A3(n1422), .A4(
        m4stg_frac[42]), .Y(n30) );
  OR2X1_RVT U152 ( .A1(n31), .A2(n30), .Y(n1129) );
  INVX1_RVT U153 ( .A(n1129), .Y(n1053) );
  INVX1_RVT U154 ( .A(m4stg_sh_cnt[2]), .Y(n1908) );
  AO22X1_RVT U155 ( .A1(n1579), .A2(m4stg_frac[48]), .A3(n1593), .A4(
        m4stg_frac[49]), .Y(n33) );
  AO22X1_RVT U156 ( .A1(n1573), .A2(m4stg_frac[47]), .A3(n1422), .A4(
        m4stg_frac[46]), .Y(n32) );
  OR2X1_RVT U157 ( .A1(n33), .A2(n32), .Y(n1047) );
  INVX1_RVT U158 ( .A(n1047), .Y(n1138) );
  NAND2X0_RVT U159 ( .A1(m4stg_sh_cnt[3]), .A2(n1908), .Y(n1616) );
  OA22X1_RVT U160 ( .A1(n1053), .A2(n1095), .A3(n1138), .A4(n1616), .Y(n37) );
  NAND2X0_RVT U161 ( .A1(n1593), .A2(m4stg_frac[53]), .Y(n211) );
  NAND2X0_RVT U162 ( .A1(n1579), .A2(m4stg_frac[52]), .Y(n119) );
  NAND2X0_RVT U163 ( .A1(n1573), .A2(m4stg_frac[51]), .Y(n410) );
  NAND2X0_RVT U164 ( .A1(n1422), .A2(m4stg_frac[50]), .Y(n34) );
  AND4X1_RVT U165 ( .A1(n211), .A2(n119), .A3(n410), .A4(n34), .Y(n1137) );
  INVX1_RVT U166 ( .A(m4stg_sh_cnt[3]), .Y(n1636) );
  NAND2X0_RVT U167 ( .A1(m4stg_sh_cnt[2]), .A2(n1636), .Y(n35) );
  INVX1_RVT U168 ( .A(n35), .Y(n1582) );
  NAND2X0_RVT U169 ( .A1(n1593), .A2(m4stg_frac[57]), .Y(n171) );
  NAND2X0_RVT U170 ( .A1(n1579), .A2(m4stg_frac[56]), .Y(n124) );
  NAND2X0_RVT U171 ( .A1(n1573), .A2(m4stg_frac[55]), .Y(n210) );
  NAND2X0_RVT U172 ( .A1(n1422), .A2(m4stg_frac[54]), .Y(n118) );
  AND4X1_RVT U173 ( .A1(n171), .A2(n124), .A3(n210), .A4(n118), .Y(n1140) );
  AND2X1_RVT U174 ( .A1(n1908), .A2(n1636), .Y(n1539) );
  INVX1_RVT U175 ( .A(n1539), .Y(n1623) );
  OA22X1_RVT U176 ( .A1(n1137), .A2(n35), .A3(n1140), .A4(n1623), .Y(n36) );
  NAND2X0_RVT U177 ( .A1(n37), .A2(n36), .Y(n1442) );
  INVX1_RVT U178 ( .A(m4stg_sh_cnt[4]), .Y(n1879) );
  NAND2X0_RVT U179 ( .A1(\m4stg_sh_cnt_5[0] ), .A2(m4stg_sh_cnt[4]), .Y(n1625)
         );
  INVX1_RVT U180 ( .A(n1625), .Y(n1647) );
  NAND2X0_RVT U181 ( .A1(n1593), .A2(m4stg_frac[65]), .Y(n75) );
  NAND2X0_RVT U182 ( .A1(n1579), .A2(m4stg_frac[64]), .Y(n102) );
  NAND2X0_RVT U183 ( .A1(n1573), .A2(m4stg_frac[63]), .Y(n78) );
  NAND2X0_RVT U184 ( .A1(n1422), .A2(m4stg_frac[62]), .Y(n105) );
  AND4X1_RVT U185 ( .A1(n75), .A2(n102), .A3(n78), .A4(n105), .Y(n1143) );
  NAND2X0_RVT U186 ( .A1(n1593), .A2(m4stg_frac[61]), .Y(n77) );
  NAND2X0_RVT U187 ( .A1(n1579), .A2(m4stg_frac[60]), .Y(n104) );
  NAND2X0_RVT U188 ( .A1(n1573), .A2(m4stg_frac[59]), .Y(n170) );
  NAND2X0_RVT U189 ( .A1(n1422), .A2(m4stg_frac[58]), .Y(n123) );
  AND4X1_RVT U190 ( .A1(n77), .A2(n104), .A3(n170), .A4(n123), .Y(n1139) );
  OA22X1_RVT U191 ( .A1(n1143), .A2(n1616), .A3(n1139), .A4(n1095), .Y(n39) );
  NAND2X0_RVT U192 ( .A1(n1593), .A2(m4stg_frac[69]), .Y(n72) );
  NAND2X0_RVT U193 ( .A1(n1579), .A2(m4stg_frac[68]), .Y(n99) );
  NAND2X0_RVT U194 ( .A1(n1573), .A2(m4stg_frac[67]), .Y(n76) );
  NAND2X0_RVT U195 ( .A1(n1422), .A2(m4stg_frac[66]), .Y(n103) );
  AND4X1_RVT U196 ( .A1(n72), .A2(n99), .A3(n76), .A4(n103), .Y(n1144) );
  NAND2X0_RVT U197 ( .A1(n1593), .A2(m4stg_frac[73]), .Y(n73) );
  NAND2X0_RVT U198 ( .A1(n1579), .A2(m4stg_frac[72]), .Y(n100) );
  NAND2X0_RVT U199 ( .A1(n1573), .A2(m4stg_frac[71]), .Y(n71) );
  NAND2X0_RVT U200 ( .A1(n1422), .A2(m4stg_frac[70]), .Y(n98) );
  AND4X1_RVT U201 ( .A1(n73), .A2(n100), .A3(n71), .A4(n98), .Y(n1145) );
  OA22X1_RVT U202 ( .A1(n1144), .A2(n35), .A3(n1145), .A4(n1623), .Y(n38) );
  NAND2X0_RVT U203 ( .A1(n39), .A2(n38), .Y(n1441) );
  AND2X1_RVT U204 ( .A1(\m4stg_sh_cnt_5[0] ), .A2(n1879), .Y(n1916) );
  NAND2X0_RVT U205 ( .A1(n1593), .A2(m4stg_frac[105]), .Y(n70) );
  NAND2X0_RVT U206 ( .A1(n1579), .A2(m4stg_frac[104]), .Y(n59) );
  NAND2X0_RVT U207 ( .A1(n1573), .A2(m4stg_frac[103]), .Y(n53) );
  NAND2X0_RVT U208 ( .A1(n1422), .A2(m4stg_frac[102]), .Y(n63) );
  NAND4X0_RVT U209 ( .A1(n70), .A2(n59), .A3(n53), .A4(n63), .Y(n41) );
  NAND2X0_RVT U210 ( .A1(n1593), .A2(m4stg_frac[101]), .Y(n52) );
  NAND2X0_RVT U211 ( .A1(n1579), .A2(m4stg_frac[100]), .Y(n62) );
  NAND2X0_RVT U212 ( .A1(n1573), .A2(m4stg_frac[99]), .Y(n54) );
  NAND2X0_RVT U213 ( .A1(n1422), .A2(m4stg_frac[98]), .Y(n40) );
  NAND4X0_RVT U214 ( .A1(n52), .A2(n62), .A3(n54), .A4(n40), .Y(n983) );
  NAND2X0_RVT U215 ( .A1(n1879), .A2(n1636), .Y(n1906) );
  INVX1_RVT U216 ( .A(n1906), .Y(n2101) );
  OAI221X1_RVT U217 ( .A1(m4stg_sh_cnt[2]), .A2(n41), .A3(n1908), .A4(n983), 
        .A5(n2101), .Y(n47) );
  AND2X1_RVT U218 ( .A1(n6), .A2(n1879), .Y(n857) );
  NAND2X0_RVT U219 ( .A1(n1593), .A2(m4stg_frac[93]), .Y(n57) );
  NAND2X0_RVT U220 ( .A1(n1579), .A2(m4stg_frac[92]), .Y(n68) );
  NAND2X0_RVT U221 ( .A1(n1573), .A2(m4stg_frac[91]), .Y(n81) );
  NAND2X0_RVT U222 ( .A1(n1422), .A2(m4stg_frac[90]), .Y(n89) );
  NAND4X0_RVT U223 ( .A1(n57), .A2(n68), .A3(n81), .A4(n89), .Y(n1046) );
  INVX1_RVT U224 ( .A(n1616), .Y(n1268) );
  AND2X1_RVT U225 ( .A1(n1268), .A2(n1879), .Y(n858) );
  NAND2X0_RVT U226 ( .A1(n1579), .A2(m4stg_frac[96]), .Y(n64) );
  NAND2X0_RVT U227 ( .A1(n1573), .A2(m4stg_frac[95]), .Y(n58) );
  NAND2X0_RVT U228 ( .A1(n1422), .A2(m4stg_frac[94]), .Y(n69) );
  NAND2X0_RVT U229 ( .A1(n1593), .A2(m4stg_frac[97]), .Y(n42) );
  NAND4X0_RVT U230 ( .A1(n64), .A2(n58), .A3(n69), .A4(n42), .Y(n1045) );
  AOI22X1_RVT U231 ( .A1(n857), .A2(n1046), .A3(n858), .A4(n1045), .Y(n46) );
  NAND2X0_RVT U232 ( .A1(n1593), .A2(m4stg_frac[81]), .Y(n85) );
  NAND2X0_RVT U233 ( .A1(n1579), .A2(m4stg_frac[80]), .Y(n93) );
  NAND2X0_RVT U234 ( .A1(n1573), .A2(m4stg_frac[79]), .Y(n88) );
  NAND2X0_RVT U235 ( .A1(n1422), .A2(m4stg_frac[78]), .Y(n96) );
  AND4X1_RVT U236 ( .A1(n85), .A2(n93), .A3(n88), .A4(n96), .Y(n1128) );
  NAND2X0_RVT U237 ( .A1(n1593), .A2(m4stg_frac[77]), .Y(n87) );
  NAND2X0_RVT U238 ( .A1(n1579), .A2(m4stg_frac[76]), .Y(n95) );
  NAND2X0_RVT U239 ( .A1(n1573), .A2(m4stg_frac[75]), .Y(n74) );
  NAND2X0_RVT U240 ( .A1(n1422), .A2(m4stg_frac[74]), .Y(n101) );
  AND4X1_RVT U241 ( .A1(n87), .A2(n95), .A3(n74), .A4(n101), .Y(n1146) );
  OA22X1_RVT U242 ( .A1(n1128), .A2(n1616), .A3(n1146), .A4(n1095), .Y(n44) );
  NAND2X0_RVT U243 ( .A1(n1593), .A2(m4stg_frac[85]), .Y(n84) );
  NAND2X0_RVT U244 ( .A1(n1579), .A2(m4stg_frac[84]), .Y(n92) );
  NAND2X0_RVT U245 ( .A1(n1573), .A2(m4stg_frac[83]), .Y(n86) );
  NAND2X0_RVT U246 ( .A1(n1422), .A2(m4stg_frac[82]), .Y(n94) );
  AND4X1_RVT U247 ( .A1(n84), .A2(n92), .A3(n86), .A4(n94), .Y(n1127) );
  NAND2X0_RVT U248 ( .A1(n1593), .A2(m4stg_frac[89]), .Y(n82) );
  NAND2X0_RVT U249 ( .A1(n1579), .A2(m4stg_frac[88]), .Y(n90) );
  NAND2X0_RVT U250 ( .A1(n1573), .A2(m4stg_frac[87]), .Y(n83) );
  NAND2X0_RVT U251 ( .A1(n1422), .A2(m4stg_frac[86]), .Y(n91) );
  AND4X1_RVT U252 ( .A1(n82), .A2(n90), .A3(n83), .A4(n91), .Y(n1125) );
  OA22X1_RVT U253 ( .A1(n1127), .A2(n35), .A3(n1125), .A4(n1623), .Y(n43) );
  NAND2X0_RVT U254 ( .A1(n44), .A2(n43), .Y(n1247) );
  NAND2X0_RVT U255 ( .A1(m4stg_sh_cnt[4]), .A2(n1247), .Y(n45) );
  NAND3X0_RVT U256 ( .A1(n47), .A2(n46), .A3(n45), .Y(n48) );
  INVX1_RVT U257 ( .A(m4stg_sh_cnt[5]), .Y(n2069) );
  AO222X1_RVT U258 ( .A1(n1442), .A2(n1647), .A3(n1441), .A4(n1916), .A5(n48), 
        .A6(n2069), .Y(m4stg_shl_55) );
  AO22X1_RVT U259 ( .A1(m2stg_frac1_dbl_dnrm), .A2(mul_frac_in1[50]), .A3(
        m2stg_frac1_sng_dnrm), .A4(mul_frac_in1[53]), .Y(n49) );
  AO221X1_RVT U260 ( .A1(m2stg_frac1_sng_norm), .A2(m1stg_snan_sng_in1), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[54]), .A5(n49), .Y(n50) );
  AOI221X1_RVT U261 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[51]), .A3(
        m2stg_frac1_dbl_norm), .A4(m1stg_snan_dbl_in1), .A5(n50), .Y(
        m2stg_frac1_array_in[51]) );
  NAND4X0_RVT U262 ( .A1(m5stg_frac_pre2[10]), .A2(m5stg_frac_pre1[10]), .A3(
        m5stg_frac_pre4[10]), .A4(m5stg_frac_pre3[10]), .Y(\add_x_3/A[7] ) );
  NAND4X0_RVT U263 ( .A1(m5stg_frac_pre2[9]), .A2(m5stg_frac_pre1[9]), .A3(
        m5stg_frac_pre4[9]), .A4(m5stg_frac_pre3[9]), .Y(\add_x_3/A[6] ) );
  INVX1_RVT U264 ( .A(se), .Y(n2148) );
  NAND4X0_RVT U265 ( .A1(m5stg_frac_pre2[30]), .A2(m5stg_frac_pre1[30]), .A3(
        m5stg_frac_pre4[30]), .A4(m5stg_frac_pre3[30]), .Y(\add_x_3/A[27] ) );
  NAND4X0_RVT U266 ( .A1(m5stg_frac_pre2[17]), .A2(m5stg_frac_pre1[17]), .A3(
        m5stg_frac_pre4[17]), .A4(m5stg_frac_pre3[17]), .Y(\add_x_3/A[14] ) );
  NAND4X0_RVT U267 ( .A1(m5stg_frac_pre2[26]), .A2(m5stg_frac_pre1[26]), .A3(
        m5stg_frac_pre4[26]), .A4(m5stg_frac_pre3[26]), .Y(\add_x_3/A[23] ) );
  NAND4X0_RVT U268 ( .A1(m5stg_frac_pre2[28]), .A2(m5stg_frac_pre1[28]), .A3(
        m5stg_frac_pre4[28]), .A4(m5stg_frac_pre3[28]), .Y(\add_x_3/A[25] ) );
  NAND4X0_RVT U269 ( .A1(m5stg_frac_pre2[3]), .A2(m5stg_frac_pre1[3]), .A3(
        m5stg_frac_pre4[3]), .A4(m5stg_frac_pre3[3]), .Y(\add_x_3/A[0] ) );
  NAND4X0_RVT U270 ( .A1(m5stg_frac_pre2[21]), .A2(m5stg_frac_pre1[21]), .A3(
        m5stg_frac_pre4[21]), .A4(m5stg_frac_pre3[21]), .Y(\add_x_3/A[18] ) );
  NAND4X0_RVT U271 ( .A1(m5stg_frac_pre2[23]), .A2(m5stg_frac_pre1[23]), .A3(
        m5stg_frac_pre4[23]), .A4(m5stg_frac_pre3[23]), .Y(\add_x_3/A[20] ) );
  NAND4X0_RVT U272 ( .A1(m5stg_frac_pre2[0]), .A2(m5stg_frac_pre1[0]), .A3(
        m5stg_frac_pre4[0]), .A4(m5stg_frac_pre3[0]), .Y(m5stg_frac_32_0[0])
         );
  NAND4X0_RVT U273 ( .A1(m5stg_frac_pre2[2]), .A2(m5stg_frac_pre1[2]), .A3(
        m5stg_frac_pre4[2]), .A4(m5stg_frac_pre3[2]), .Y(m5stg_frac_32_0[2])
         );
  NAND4X0_RVT U274 ( .A1(m5stg_frac_pre2[1]), .A2(m5stg_frac_pre1[1]), .A3(
        m5stg_frac_pre4[1]), .A4(m5stg_frac_pre3[1]), .Y(m5stg_frac_32_0[1])
         );
  OR3X2_RVT U275 ( .A1(m5stg_frac_32_0[0]), .A2(m5stg_frac_32_0[2]), .A3(
        m5stg_frac_32_0[1]), .Y(m5stg_frac_dbl_nx) );
  NAND4X0_RVT U276 ( .A1(m5stg_frac_pre2[29]), .A2(m5stg_frac_pre1[29]), .A3(
        m5stg_frac_pre4[29]), .A4(m5stg_frac_pre3[29]), .Y(\add_x_3/A[26] ) );
  NAND4X0_RVT U277 ( .A1(m5stg_frac_pre2[27]), .A2(m5stg_frac_pre1[27]), .A3(
        m5stg_frac_pre4[27]), .A4(m5stg_frac_pre3[27]), .Y(\add_x_3/A[24] ) );
  NAND2X0_RVT U278 ( .A1(n1879), .A2(n2069), .Y(n437) );
  AND4X1_RVT U279 ( .A1(n1539), .A2(n154), .A3(n2087), .A4(
        m4stg_right_shift_step), .Y(n2043) );
  AO22X1_RVT U280 ( .A1(n1579), .A2(m4stg_frac[105]), .A3(n1593), .A4(
        m4stg_frac[104]), .Y(n234) );
  NAND2X0_RVT U281 ( .A1(n2043), .A2(n234), .Y(n1769) );
  INVX1_RVT U282 ( .A(n234), .Y(n284) );
  AO22X1_RVT U283 ( .A1(m4stg_sh_cnt[0]), .A2(m4stg_frac[101]), .A3(n778), 
        .A4(m4stg_frac[100]), .Y(n223) );
  AOI222X1_RVT U284 ( .A1(n223), .A2(n975), .A3(n1573), .A4(m4stg_frac[102]), 
        .A5(m4stg_frac[103]), .A6(n1422), .Y(n246) );
  AO22X1_RVT U285 ( .A1(m4stg_sh_cnt[2]), .A2(n284), .A3(n1908), .A4(n246), 
        .Y(n316) );
  INVX1_RVT U286 ( .A(n316), .Y(n2098) );
  NAND2X0_RVT U287 ( .A1(n2043), .A2(n2098), .Y(n1765) );
  NAND2X0_RVT U288 ( .A1(n1422), .A2(m4stg_frac[104]), .Y(n51) );
  NAND2X0_RVT U289 ( .A1(n1579), .A2(m4stg_frac[102]), .Y(n838) );
  AND4X1_RVT U290 ( .A1(n53), .A2(n52), .A3(n51), .A4(n838), .Y(n147) );
  AO22X1_RVT U291 ( .A1(m4stg_sh_cnt[2]), .A2(n70), .A3(n1908), .A4(n147), .Y(
        n2036) );
  NAND2X0_RVT U292 ( .A1(n1422), .A2(m4stg_frac[100]), .Y(n839) );
  AND2X1_RVT U293 ( .A1(n54), .A2(n839), .Y(n56) );
  AOI22X1_RVT U294 ( .A1(m4stg_sh_cnt[0]), .A2(n841), .A3(n778), .A4(n843), 
        .Y(n65) );
  NAND2X0_RVT U295 ( .A1(n975), .A2(n65), .Y(n55) );
  AND2X1_RVT U296 ( .A1(n56), .A2(n55), .Y(n148) );
  NAND2X0_RVT U297 ( .A1(n1422), .A2(m4stg_frac[96]), .Y(n845) );
  NAND2X0_RVT U298 ( .A1(n1579), .A2(m4stg_frac[94]), .Y(n849) );
  AND4X1_RVT U299 ( .A1(n58), .A2(n57), .A3(n845), .A4(n849), .Y(n186) );
  OAI222X1_RVT U300 ( .A1(n1636), .A2(n2036), .A3(n35), .A4(n148), .A5(n1623), 
        .A6(n186), .Y(n2091) );
  NAND2X0_RVT U301 ( .A1(n2043), .A2(n2091), .Y(n1758) );
  NAND2X0_RVT U302 ( .A1(n1593), .A2(m4stg_frac[103]), .Y(n837) );
  AND2X1_RVT U303 ( .A1(n837), .A2(n59), .Y(n61) );
  NAND2X0_RVT U304 ( .A1(m4stg_frac[105]), .A2(n1573), .Y(n60) );
  AND2X1_RVT U305 ( .A1(n61), .A2(n60), .Y(n127) );
  NAND2X0_RVT U306 ( .A1(n1573), .A2(m4stg_frac[101]), .Y(n840) );
  NAND2X0_RVT U307 ( .A1(n1593), .A2(m4stg_frac[99]), .Y(n846) );
  AND4X1_RVT U308 ( .A1(n63), .A2(n62), .A3(n840), .A4(n846), .Y(n128) );
  AO22X1_RVT U309 ( .A1(m4stg_sh_cnt[2]), .A2(n127), .A3(n1908), .A4(n128), 
        .Y(n2037) );
  NAND2X0_RVT U310 ( .A1(n1593), .A2(m4stg_frac[95]), .Y(n851) );
  AND2X1_RVT U311 ( .A1(n851), .A2(n64), .Y(n67) );
  NAND2X0_RVT U312 ( .A1(n65), .A2(m4stg_sh_cnt[1]), .Y(n66) );
  AND2X1_RVT U313 ( .A1(n67), .A2(n66), .Y(n129) );
  NAND2X0_RVT U314 ( .A1(n1573), .A2(m4stg_frac[93]), .Y(n852) );
  NAND2X0_RVT U315 ( .A1(n1593), .A2(m4stg_frac[91]), .Y(n856) );
  AND4X1_RVT U316 ( .A1(n69), .A2(n68), .A3(n852), .A4(n856), .Y(n203) );
  OA222X1_RVT U317 ( .A1(n1636), .A2(n2037), .A3(n35), .A4(n129), .A5(n1623), 
        .A6(n203), .Y(n448) );
  INVX1_RVT U318 ( .A(n448), .Y(n2089) );
  NAND2X0_RVT U319 ( .A1(n2043), .A2(n2089), .Y(n1756) );
  OA222X1_RVT U320 ( .A1(n35), .A2(n128), .A3(n1623), .A4(n129), .A5(n1616), 
        .A6(n127), .Y(n407) );
  INVX1_RVT U321 ( .A(n407), .Y(n2093) );
  NAND2X0_RVT U322 ( .A1(n2043), .A2(n2093), .Y(n1760) );
  OA222X1_RVT U323 ( .A1(n1616), .A2(n70), .A3(n1623), .A4(n148), .A5(n35), 
        .A6(n147), .Y(n404) );
  INVX1_RVT U324 ( .A(n404), .Y(n2095) );
  NAND2X0_RVT U325 ( .A1(n2043), .A2(n2095), .Y(n1762) );
  NAND2X0_RVT U326 ( .A1(n1422), .A2(m4stg_frac[72]), .Y(n866) );
  NAND2X0_RVT U327 ( .A1(n1579), .A2(m4stg_frac[70]), .Y(n908) );
  NAND4X0_RVT U328 ( .A1(n72), .A2(n71), .A3(n866), .A4(n908), .Y(n181) );
  NAND2X0_RVT U329 ( .A1(n1422), .A2(m4stg_frac[76]), .Y(n862) );
  NAND2X0_RVT U330 ( .A1(n1579), .A2(m4stg_frac[74]), .Y(n865) );
  AND4X1_RVT U331 ( .A1(n74), .A2(n73), .A3(n862), .A4(n865), .Y(n178) );
  OA22X1_RVT U332 ( .A1(n169), .A2(n1616), .A3(n178), .A4(n1095), .Y(n80) );
  NAND2X0_RVT U333 ( .A1(n1422), .A2(m4stg_frac[68]), .Y(n909) );
  NAND2X0_RVT U334 ( .A1(n1579), .A2(m4stg_frac[66]), .Y(n905) );
  NAND4X0_RVT U335 ( .A1(n76), .A2(n75), .A3(n909), .A4(n905), .Y(n176) );
  INVX1_RVT U336 ( .A(n176), .Y(n213) );
  NAND2X0_RVT U337 ( .A1(n1422), .A2(m4stg_frac[64]), .Y(n904) );
  NAND2X0_RVT U338 ( .A1(n1579), .A2(m4stg_frac[62]), .Y(n897) );
  NAND4X0_RVT U339 ( .A1(n78), .A2(n77), .A3(n904), .A4(n897), .Y(n363) );
  INVX1_RVT U340 ( .A(n363), .Y(n212) );
  OA22X1_RVT U341 ( .A1(n213), .A2(n35), .A3(n212), .A4(n1623), .Y(n79) );
  NAND2X0_RVT U342 ( .A1(n80), .A2(n79), .Y(n373) );
  NAND2X0_RVT U343 ( .A1(m4stg_sh_cnt[5]), .A2(n1879), .Y(n257) );
  NAND2X0_RVT U344 ( .A1(m4stg_sh_cnt[4]), .A2(n2069), .Y(n397) );
  NAND2X0_RVT U345 ( .A1(n1422), .A2(m4stg_frac[92]), .Y(n850) );
  NAND2X0_RVT U346 ( .A1(n1579), .A2(m4stg_frac[90]), .Y(n854) );
  NAND4X0_RVT U347 ( .A1(n82), .A2(n81), .A3(n850), .A4(n854), .Y(n184) );
  NAND2X0_RVT U348 ( .A1(n1422), .A2(m4stg_frac[88]), .Y(n853) );
  NAND2X0_RVT U349 ( .A1(n1579), .A2(m4stg_frac[86]), .Y(n873) );
  NAND4X0_RVT U350 ( .A1(n84), .A2(n83), .A3(n853), .A4(n873), .Y(n189) );
  OAI22X1_RVT U351 ( .A1(n1908), .A2(n184), .A3(m4stg_sh_cnt[2]), .A4(n189), 
        .Y(n135) );
  NAND2X0_RVT U352 ( .A1(n1422), .A2(m4stg_frac[84]), .Y(n871) );
  NAND2X0_RVT U353 ( .A1(n1579), .A2(m4stg_frac[82]), .Y(n867) );
  AND4X1_RVT U354 ( .A1(n86), .A2(n85), .A3(n871), .A4(n867), .Y(n185) );
  NAND2X0_RVT U355 ( .A1(n1422), .A2(m4stg_frac[80]), .Y(n870) );
  NAND2X0_RVT U356 ( .A1(n1579), .A2(m4stg_frac[78]), .Y(n861) );
  AND4X1_RVT U357 ( .A1(n88), .A2(n87), .A3(n870), .A4(n861), .Y(n177) );
  OA222X1_RVT U358 ( .A1(n1636), .A2(n135), .A3(n35), .A4(n185), .A5(n1623), 
        .A6(n177), .Y(n380) );
  INVX1_RVT U359 ( .A(n380), .Y(n405) );
  AO222X1_RVT U360 ( .A1(n2087), .A2(n373), .A3(n1916), .A4(n2091), .A5(n1651), 
        .A6(n405), .Y(n2056) );
  NAND2X0_RVT U361 ( .A1(n2043), .A2(n2056), .Y(n1726) );
  NAND2X0_RVT U362 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .Y(n375) );
  NAND2X0_RVT U363 ( .A1(n1573), .A2(m4stg_frac[89]), .Y(n855) );
  NAND2X0_RVT U364 ( .A1(n1593), .A2(m4stg_frac[87]), .Y(n874) );
  NAND4X0_RVT U365 ( .A1(n90), .A2(n89), .A3(n855), .A4(n874), .Y(n201) );
  NAND2X0_RVT U366 ( .A1(n1573), .A2(m4stg_frac[85]), .Y(n872) );
  NAND2X0_RVT U367 ( .A1(n1593), .A2(m4stg_frac[83]), .Y(n869) );
  NAND4X0_RVT U368 ( .A1(n92), .A2(n91), .A3(n872), .A4(n869), .Y(n206) );
  OAI22X1_RVT U369 ( .A1(n1908), .A2(n201), .A3(m4stg_sh_cnt[2]), .A4(n206), 
        .Y(n111) );
  NAND2X0_RVT U370 ( .A1(n1573), .A2(m4stg_frac[81]), .Y(n868) );
  NAND2X0_RVT U371 ( .A1(n1593), .A2(m4stg_frac[79]), .Y(n859) );
  AND4X1_RVT U372 ( .A1(n94), .A2(n93), .A3(n868), .A4(n859), .Y(n202) );
  NAND2X0_RVT U373 ( .A1(n1573), .A2(m4stg_frac[77]), .Y(n860) );
  NAND2X0_RVT U374 ( .A1(n1593), .A2(m4stg_frac[75]), .Y(n863) );
  AND4X1_RVT U375 ( .A1(n96), .A2(n95), .A3(n860), .A4(n863), .Y(n194) );
  OA222X1_RVT U376 ( .A1(n1636), .A2(n111), .A3(n35), .A4(n202), .A5(n1623), 
        .A6(n194), .Y(n447) );
  AOI22X1_RVT U377 ( .A1(m4stg_sh_cnt[4]), .A2(n447), .A3(m4stg_sh_cnt[5]), 
        .A4(n448), .Y(n97) );
  AND2X1_RVT U378 ( .A1(n375), .A2(n97), .Y(n110) );
  NAND2X0_RVT U379 ( .A1(n1573), .A2(m4stg_frac[69]), .Y(n907) );
  NAND2X0_RVT U380 ( .A1(n1593), .A2(m4stg_frac[67]), .Y(n902) );
  NAND4X0_RVT U381 ( .A1(n99), .A2(n98), .A3(n907), .A4(n902), .Y(n198) );
  NAND2X0_RVT U382 ( .A1(n1573), .A2(m4stg_frac[73]), .Y(n864) );
  NAND2X0_RVT U383 ( .A1(n1593), .A2(m4stg_frac[71]), .Y(n906) );
  AND4X1_RVT U384 ( .A1(n101), .A2(n100), .A3(n864), .A4(n906), .Y(n195) );
  OA22X1_RVT U385 ( .A1(n162), .A2(n1616), .A3(n195), .A4(n1095), .Y(n107) );
  NAND2X0_RVT U386 ( .A1(n1573), .A2(m4stg_frac[65]), .Y(n903) );
  NAND2X0_RVT U387 ( .A1(n1593), .A2(m4stg_frac[63]), .Y(n895) );
  NAND4X0_RVT U388 ( .A1(n103), .A2(n102), .A3(n903), .A4(n895), .Y(n193) );
  INVX1_RVT U389 ( .A(n193), .Y(n163) );
  NAND2X0_RVT U390 ( .A1(n1573), .A2(m4stg_frac[61]), .Y(n894) );
  NAND2X0_RVT U391 ( .A1(n1593), .A2(m4stg_frac[59]), .Y(n900) );
  NAND4X0_RVT U392 ( .A1(n105), .A2(n104), .A3(n894), .A4(n900), .Y(n362) );
  INVX1_RVT U393 ( .A(n362), .Y(n120) );
  OA22X1_RVT U394 ( .A1(n163), .A2(n35), .A3(n120), .A4(n1623), .Y(n106) );
  NAND2X0_RVT U395 ( .A1(n107), .A2(n106), .Y(n390) );
  NAND2X0_RVT U396 ( .A1(n108), .A2(n2087), .Y(n109) );
  AND2X1_RVT U397 ( .A1(n110), .A2(n109), .Y(n2054) );
  NAND2X0_RVT U398 ( .A1(n2043), .A2(n2054), .Y(n1724) );
  INVX1_RVT U399 ( .A(n6), .Y(n1095) );
  OA222X1_RVT U400 ( .A1(n1095), .A2(n129), .A3(n1616), .A4(n203), .A5(n111), 
        .A6(m4stg_sh_cnt[3]), .Y(n394) );
  NAND2X0_RVT U401 ( .A1(m4stg_sh_cnt[4]), .A2(n1636), .Y(n317) );
  OAI22X1_RVT U402 ( .A1(m4stg_sh_cnt[4]), .A2(n394), .A3(n2037), .A4(n317), 
        .Y(n2079) );
  NAND2X0_RVT U403 ( .A1(n2043), .A2(n2079), .Y(n1748) );
  NAND2X0_RVT U404 ( .A1(n2101), .A2(m4stg_sh_cnt[5]), .Y(n283) );
  NAND2X0_RVT U405 ( .A1(n1539), .A2(n198), .Y(n113) );
  OA22X1_RVT U406 ( .A1(n194), .A2(n1616), .A3(n202), .A4(n1095), .Y(n112) );
  AND2X1_RVT U407 ( .A1(n113), .A2(n112), .Y(n116) );
  NAND2X0_RVT U408 ( .A1(n114), .A2(n1582), .Y(n115) );
  AND2X1_RVT U409 ( .A1(n116), .A2(n115), .Y(n117) );
  OAI222X1_RVT U410 ( .A1(n2037), .A2(n283), .A3(n397), .A4(n394), .A5(n437), 
        .A6(n117), .Y(n2062) );
  NAND2X0_RVT U411 ( .A1(n2043), .A2(n2062), .Y(n1732) );
  INVX1_RVT U412 ( .A(n117), .Y(n391) );
  NAND2X0_RVT U413 ( .A1(n1573), .A2(m4stg_frac[53]), .Y(n890) );
  NAND2X0_RVT U414 ( .A1(n1593), .A2(m4stg_frac[51]), .Y(n885) );
  NAND4X0_RVT U415 ( .A1(n119), .A2(n118), .A3(n890), .A4(n885), .Y(n355) );
  NAND2X0_RVT U416 ( .A1(n1539), .A2(n355), .Y(n122) );
  OA22X1_RVT U417 ( .A1(n163), .A2(n1095), .A3(n120), .A4(n1616), .Y(n121) );
  AND2X1_RVT U418 ( .A1(n122), .A2(n121), .Y(n126) );
  NAND2X0_RVT U419 ( .A1(n1573), .A2(m4stg_frac[57]), .Y(n898) );
  NAND2X0_RVT U420 ( .A1(n1593), .A2(m4stg_frac[55]), .Y(n889) );
  NAND4X0_RVT U421 ( .A1(n124), .A2(n123), .A3(n898), .A4(n889), .Y(n357) );
  NAND2X0_RVT U422 ( .A1(n357), .A2(n1582), .Y(n125) );
  AND2X1_RVT U423 ( .A1(n126), .A2(n125), .Y(n426) );
  INVX1_RVT U424 ( .A(n426), .Y(n420) );
  AO222X1_RVT U425 ( .A1(n1651), .A2(n391), .A3(n2087), .A4(n420), .A5(
        m4stg_sh_cnt[5]), .A6(n2079), .Y(n2046) );
  NAND2X0_RVT U426 ( .A1(n2043), .A2(n2046), .Y(n1716) );
  INVX1_RVT U427 ( .A(n127), .Y(n2103) );
  NAND2X0_RVT U428 ( .A1(n1539), .A2(n2103), .Y(n146) );
  NAND2X0_RVT U429 ( .A1(n1539), .A2(n201), .Y(n131) );
  OA22X1_RVT U430 ( .A1(n129), .A2(n1616), .A3(n128), .A4(n1095), .Y(n130) );
  AND2X1_RVT U431 ( .A1(n131), .A2(n130), .Y(n134) );
  NAND2X0_RVT U432 ( .A1(n132), .A2(n1582), .Y(n133) );
  AND2X1_RVT U433 ( .A1(n134), .A2(n133), .Y(n379) );
  AO22X1_RVT U434 ( .A1(m4stg_sh_cnt[4]), .A2(n146), .A3(n1879), .A4(n379), 
        .Y(n168) );
  INVX1_RVT U435 ( .A(n168), .Y(n2083) );
  NAND2X0_RVT U436 ( .A1(n2043), .A2(n2083), .Y(n1752) );
  OA222X1_RVT U437 ( .A1(n1095), .A2(n148), .A3(n1616), .A4(n186), .A5(n135), 
        .A6(m4stg_sh_cnt[3]), .Y(n377) );
  NAND2X0_RVT U438 ( .A1(n1539), .A2(n181), .Y(n137) );
  OA22X1_RVT U439 ( .A1(n177), .A2(n1616), .A3(n185), .A4(n1095), .Y(n136) );
  AND2X1_RVT U440 ( .A1(n137), .A2(n136), .Y(n140) );
  NAND2X0_RVT U441 ( .A1(n138), .A2(n1582), .Y(n139) );
  AND2X1_RVT U442 ( .A1(n140), .A2(n139), .Y(n423) );
  OAI222X1_RVT U443 ( .A1(n283), .A2(n2036), .A3(n397), .A4(n377), .A5(n437), 
        .A6(n423), .Y(n2064) );
  NAND2X0_RVT U444 ( .A1(n2043), .A2(n2064), .Y(n1734) );
  NAND2X0_RVT U445 ( .A1(n6), .A2(n206), .Y(n142) );
  OA22X1_RVT U446 ( .A1(n195), .A2(n1623), .A3(n202), .A4(n1616), .Y(n141) );
  AND2X1_RVT U447 ( .A1(n142), .A2(n141), .Y(n145) );
  NAND2X0_RVT U448 ( .A1(n143), .A2(n1582), .Y(n144) );
  AND2X1_RVT U449 ( .A1(n145), .A2(n144), .Y(n425) );
  OAI222X1_RVT U450 ( .A1(n146), .A2(n257), .A3(n437), .A4(n425), .A5(n397), 
        .A6(n379), .Y(n2066) );
  NAND2X0_RVT U451 ( .A1(n2043), .A2(n2066), .Y(n1736) );
  NAND2X0_RVT U452 ( .A1(n1539), .A2(n184), .Y(n150) );
  OA22X1_RVT U453 ( .A1(n148), .A2(n1616), .A3(n147), .A4(n1095), .Y(n149) );
  AND2X1_RVT U454 ( .A1(n150), .A2(n149), .Y(n153) );
  NAND2X0_RVT U455 ( .A1(n151), .A2(n1582), .Y(n152) );
  AND2X1_RVT U456 ( .A1(n153), .A2(n152), .Y(n428) );
  INVX1_RVT U457 ( .A(n428), .Y(n161) );
  OA222X1_RVT U458 ( .A1(n1879), .A2(n1539), .A3(n1879), .A4(n154), .A5(
        m4stg_sh_cnt[4]), .A6(n161), .Y(n2085) );
  NAND2X0_RVT U459 ( .A1(n2043), .A2(n2085), .Y(n1754) );
  NAND2X0_RVT U460 ( .A1(n6), .A2(n189), .Y(n156) );
  OA22X1_RVT U461 ( .A1(n178), .A2(n1623), .A3(n185), .A4(n1616), .Y(n155) );
  AND2X1_RVT U462 ( .A1(n156), .A2(n155), .Y(n159) );
  NAND2X0_RVT U463 ( .A1(n157), .A2(n1582), .Y(n158) );
  AND2X1_RVT U464 ( .A1(n159), .A2(n158), .Y(n382) );
  INVX1_RVT U465 ( .A(n382), .Y(n175) );
  AND3X1_RVT U466 ( .A1(n1593), .A2(n1539), .A3(m4stg_frac[105]), .Y(n160) );
  AO222X1_RVT U467 ( .A1(n161), .A2(n1651), .A3(n175), .A4(n2087), .A5(n160), 
        .A6(n1916), .Y(n2068) );
  NAND2X0_RVT U468 ( .A1(n2043), .A2(n2068), .Y(n1738) );
  NAND2X0_RVT U469 ( .A1(n1539), .A2(n357), .Y(n165) );
  OA22X1_RVT U470 ( .A1(n163), .A2(n1616), .A3(n162), .A4(n1095), .Y(n164) );
  AND2X1_RVT U471 ( .A1(n165), .A2(n164), .Y(n167) );
  NAND2X0_RVT U472 ( .A1(n362), .A2(n1582), .Y(n166) );
  AND2X1_RVT U473 ( .A1(n167), .A2(n166), .Y(n435) );
  OAI222X1_RVT U474 ( .A1(n168), .A2(n2069), .A3(n437), .A4(n435), .A5(n397), 
        .A6(n425), .Y(n2050) );
  NAND2X0_RVT U475 ( .A1(n2043), .A2(n2050), .Y(n1720) );
  OA22X1_RVT U476 ( .A1(n213), .A2(n1616), .A3(n169), .A4(n1095), .Y(n174) );
  NAND2X0_RVT U477 ( .A1(n1422), .A2(m4stg_frac[60]), .Y(n896) );
  NAND2X0_RVT U478 ( .A1(n1579), .A2(m4stg_frac[58]), .Y(n901) );
  NAND4X0_RVT U479 ( .A1(n171), .A2(n170), .A3(n896), .A4(n901), .Y(n417) );
  OA22X1_RVT U480 ( .A1(n212), .A2(n35), .A3(n172), .A4(n1623), .Y(n173) );
  NAND2X0_RVT U481 ( .A1(n174), .A2(n173), .Y(n332) );
  AO222X1_RVT U482 ( .A1(n175), .A2(n1651), .A3(n332), .A4(n2087), .A5(n2085), 
        .A6(m4stg_sh_cnt[5]), .Y(n2052) );
  NAND2X0_RVT U483 ( .A1(n2043), .A2(n2052), .Y(n1722) );
  NAND2X0_RVT U484 ( .A1(n1539), .A2(n176), .Y(n180) );
  OA22X1_RVT U485 ( .A1(n178), .A2(n1616), .A3(n177), .A4(n1095), .Y(n179) );
  AND2X1_RVT U486 ( .A1(n180), .A2(n179), .Y(n183) );
  NAND2X0_RVT U487 ( .A1(n181), .A2(n1582), .Y(n182) );
  AND2X1_RVT U488 ( .A1(n183), .A2(n182), .Y(n326) );
  NAND2X0_RVT U489 ( .A1(n1268), .A2(n184), .Y(n188) );
  OA22X1_RVT U490 ( .A1(n186), .A2(n1095), .A3(n185), .A4(n1623), .Y(n187) );
  AND2X1_RVT U491 ( .A1(n188), .A2(n187), .Y(n191) );
  NAND2X0_RVT U492 ( .A1(n189), .A2(n1582), .Y(n190) );
  AND2X1_RVT U493 ( .A1(n191), .A2(n190), .Y(n403) );
  AO222X1_RVT U494 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .A3(
        m4stg_sh_cnt[4]), .A4(n403), .A5(m4stg_sh_cnt[5]), .A6(n404), .Y(n192)
         );
  AOI21X1_RVT U495 ( .A1(n326), .A2(n2087), .A3(n192), .Y(n2060) );
  NAND2X0_RVT U496 ( .A1(n2043), .A2(n2060), .Y(n1730) );
  NAND2X0_RVT U497 ( .A1(n1539), .A2(n193), .Y(n197) );
  OA22X1_RVT U498 ( .A1(n195), .A2(n1616), .A3(n194), .A4(n1095), .Y(n196) );
  AND2X1_RVT U499 ( .A1(n197), .A2(n196), .Y(n200) );
  NAND2X0_RVT U500 ( .A1(n198), .A2(n1582), .Y(n199) );
  AND2X1_RVT U501 ( .A1(n200), .A2(n199), .Y(n330) );
  NAND2X0_RVT U502 ( .A1(n1268), .A2(n201), .Y(n205) );
  OA22X1_RVT U503 ( .A1(n203), .A2(n1095), .A3(n202), .A4(n1623), .Y(n204) );
  AND2X1_RVT U504 ( .A1(n205), .A2(n204), .Y(n208) );
  NAND2X0_RVT U505 ( .A1(n206), .A2(n1582), .Y(n207) );
  AND2X1_RVT U506 ( .A1(n208), .A2(n207), .Y(n406) );
  AO222X1_RVT U507 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .A3(
        m4stg_sh_cnt[4]), .A4(n406), .A5(m4stg_sh_cnt[5]), .A6(n407), .Y(n209)
         );
  AOI21X1_RVT U508 ( .A1(n330), .A2(n2087), .A3(n209), .Y(n2058) );
  NAND2X0_RVT U509 ( .A1(n2043), .A2(n2058), .Y(n1728) );
  OA22X1_RVT U510 ( .A1(m4stg_sh_cnt[4]), .A2(n377), .A3(n2036), .A4(n317), 
        .Y(n218) );
  INVX1_RVT U511 ( .A(n218), .Y(n2081) );
  NAND2X0_RVT U512 ( .A1(n2043), .A2(n2081), .Y(n1750) );
  NAND2X0_RVT U513 ( .A1(n1422), .A2(m4stg_frac[56]), .Y(n899) );
  NAND2X0_RVT U514 ( .A1(n1579), .A2(m4stg_frac[54]), .Y(n891) );
  NAND4X0_RVT U515 ( .A1(n211), .A2(n210), .A3(n899), .A4(n891), .Y(n359) );
  NAND2X0_RVT U516 ( .A1(n1539), .A2(n359), .Y(n215) );
  OA22X1_RVT U517 ( .A1(n213), .A2(n1095), .A3(n212), .A4(n1616), .Y(n214) );
  AND2X1_RVT U518 ( .A1(n215), .A2(n214), .Y(n217) );
  NAND2X0_RVT U519 ( .A1(n417), .A2(n1582), .Y(n216) );
  AND2X1_RVT U520 ( .A1(n217), .A2(n216), .Y(n433) );
  OAI222X1_RVT U521 ( .A1(n397), .A2(n423), .A3(n437), .A4(n433), .A5(n2069), 
        .A6(n218), .Y(n2048) );
  NAND2X0_RVT U522 ( .A1(n2043), .A2(n2048), .Y(n1718) );
  NAND4X0_RVT U523 ( .A1(m5stg_frac_pre2[32]), .A2(m5stg_frac_pre1[32]), .A3(
        m5stg_frac_pre4[32]), .A4(m5stg_frac_pre3[32]), .Y(\add_x_3/A[29] ) );
  NAND4X0_RVT U524 ( .A1(m5stg_frac_pre2[25]), .A2(m5stg_frac_pre1[25]), .A3(
        m5stg_frac_pre4[25]), .A4(m5stg_frac_pre3[25]), .Y(\add_x_3/A[22] ) );
  NAND4X0_RVT U525 ( .A1(m5stg_frac_pre2[18]), .A2(m5stg_frac_pre1[18]), .A3(
        m5stg_frac_pre4[18]), .A4(m5stg_frac_pre3[18]), .Y(\add_x_3/A[15] ) );
  NAND4X0_RVT U526 ( .A1(m5stg_frac_pre2[24]), .A2(m5stg_frac_pre1[24]), .A3(
        m5stg_frac_pre4[24]), .A4(m5stg_frac_pre3[24]), .Y(\add_x_3/A[21] ) );
  NAND4X0_RVT U527 ( .A1(m5stg_frac_pre2[22]), .A2(m5stg_frac_pre1[22]), .A3(
        m5stg_frac_pre4[22]), .A4(m5stg_frac_pre3[22]), .Y(\add_x_3/A[19] ) );
  NAND4X0_RVT U528 ( .A1(m5stg_frac_pre2[16]), .A2(m5stg_frac_pre1[16]), .A3(
        m5stg_frac_pre4[16]), .A4(m5stg_frac_pre3[16]), .Y(\add_x_3/A[13] ) );
  NAND4X0_RVT U529 ( .A1(m5stg_frac_pre2[15]), .A2(m5stg_frac_pre1[15]), .A3(
        m5stg_frac_pre4[15]), .A4(m5stg_frac_pre3[15]), .Y(\add_x_3/A[12] ) );
  NAND4X0_RVT U530 ( .A1(m5stg_frac_pre2[14]), .A2(m5stg_frac_pre1[14]), .A3(
        m5stg_frac_pre4[14]), .A4(m5stg_frac_pre3[14]), .Y(\add_x_3/A[11] ) );
  NAND4X0_RVT U531 ( .A1(m5stg_frac_pre2[13]), .A2(m5stg_frac_pre1[13]), .A3(
        m5stg_frac_pre4[13]), .A4(m5stg_frac_pre3[13]), .Y(\add_x_3/A[10] ) );
  NAND4X0_RVT U532 ( .A1(m5stg_frac_pre2[12]), .A2(m5stg_frac_pre1[12]), .A3(
        m5stg_frac_pre4[12]), .A4(m5stg_frac_pre3[12]), .Y(\add_x_3/A[9] ) );
  NAND4X0_RVT U533 ( .A1(m5stg_frac_pre2[8]), .A2(m5stg_frac_pre1[8]), .A3(
        m5stg_frac_pre4[8]), .A4(m5stg_frac_pre3[8]), .Y(\add_x_3/A[5] ) );
  NAND4X0_RVT U534 ( .A1(m5stg_frac_pre2[5]), .A2(m5stg_frac_pre1[5]), .A3(
        m5stg_frac_pre4[5]), .A4(m5stg_frac_pre3[5]), .Y(\add_x_3/A[2] ) );
  NAND4X0_RVT U535 ( .A1(m5stg_frac_pre2[11]), .A2(m5stg_frac_pre1[11]), .A3(
        m5stg_frac_pre4[11]), .A4(m5stg_frac_pre3[11]), .Y(\add_x_3/A[8] ) );
  NAND4X0_RVT U536 ( .A1(m5stg_frac_pre2[7]), .A2(m5stg_frac_pre1[7]), .A3(
        m5stg_frac_pre4[7]), .A4(m5stg_frac_pre3[7]), .Y(\add_x_3/A[4] ) );
  NAND4X0_RVT U537 ( .A1(m5stg_frac_pre2[6]), .A2(m5stg_frac_pre1[6]), .A3(
        m5stg_frac_pre4[6]), .A4(m5stg_frac_pre3[6]), .Y(\add_x_3/A[3] ) );
  NAND4X0_RVT U538 ( .A1(m5stg_frac_pre2[31]), .A2(m5stg_frac_pre1[31]), .A3(
        m5stg_frac_pre4[31]), .A4(m5stg_frac_pre3[31]), .Y(\add_x_3/A[28] ) );
  NAND4X0_RVT U539 ( .A1(m5stg_frac_pre2[4]), .A2(m5stg_frac_pre1[4]), .A3(
        m5stg_frac_pre4[4]), .A4(m5stg_frac_pre3[4]), .Y(\add_x_3/A[1] ) );
  AOI22X1_RVT U540 ( .A1(n1422), .A2(m4stg_frac[97]), .A3(n1579), .A4(
        m4stg_frac[95]), .Y(n219) );
  NAND2X0_RVT U541 ( .A1(n1573), .A2(m4stg_frac[96]), .Y(n972) );
  NAND2X0_RVT U542 ( .A1(n1593), .A2(m4stg_frac[94]), .Y(n916) );
  NAND3X0_RVT U543 ( .A1(n219), .A2(n972), .A3(n916), .Y(n273) );
  NAND2X0_RVT U544 ( .A1(n1573), .A2(m4stg_frac[92]), .Y(n917) );
  NAND2X0_RVT U545 ( .A1(n1422), .A2(m4stg_frac[93]), .Y(n220) );
  NAND2X0_RVT U546 ( .A1(n1579), .A2(m4stg_frac[91]), .Y(n771) );
  NAND2X0_RVT U547 ( .A1(n1593), .A2(m4stg_frac[90]), .Y(n921) );
  NAND4X0_RVT U548 ( .A1(n917), .A2(n220), .A3(n771), .A4(n921), .Y(n262) );
  AOI22X1_RVT U549 ( .A1(n1422), .A2(m4stg_frac[105]), .A3(n1593), .A4(
        m4stg_frac[102]), .Y(n222) );
  NAND2X0_RVT U550 ( .A1(n1579), .A2(m4stg_frac[103]), .Y(n777) );
  NAND2X0_RVT U551 ( .A1(m4stg_frac[104]), .A2(n1573), .Y(n221) );
  NAND3X0_RVT U552 ( .A1(n222), .A2(n777), .A3(n221), .Y(n2102) );
  AO22X1_RVT U553 ( .A1(m4stg_sh_cnt[1]), .A2(n223), .A3(n1593), .A4(
        m4stg_frac[98]), .Y(n224) );
  AO21X1_RVT U554 ( .A1(n1579), .A2(m4stg_frac[99]), .A3(n224), .Y(n252) );
  AO22X1_RVT U555 ( .A1(m4stg_sh_cnt[2]), .A2(n2102), .A3(n1908), .A4(n252), 
        .Y(n2096) );
  AO222X1_RVT U556 ( .A1(n273), .A2(n1582), .A3(n262), .A4(n1539), .A5(n2096), 
        .A6(m4stg_sh_cnt[3]), .Y(n2088) );
  NAND2X0_RVT U557 ( .A1(n2043), .A2(n2088), .Y(n1755) );
  AO222X1_RVT U558 ( .A1(n1582), .A2(n252), .A3(n1539), .A4(n273), .A5(n1268), 
        .A6(n2102), .Y(n2092) );
  NAND2X0_RVT U559 ( .A1(n2043), .A2(n2092), .Y(n1759) );
  NAND2X0_RVT U560 ( .A1(n1579), .A2(m4stg_frac[97]), .Y(n969) );
  AOI22X1_RVT U561 ( .A1(n1422), .A2(m4stg_frac[99]), .A3(n1593), .A4(
        m4stg_frac[96]), .Y(n225) );
  AND2X1_RVT U562 ( .A1(n969), .A2(n225), .Y(n227) );
  NAND2X0_RVT U563 ( .A1(m4stg_frac[98]), .A2(n1573), .Y(n226) );
  AND2X1_RVT U564 ( .A1(n227), .A2(n226), .Y(n245) );
  NAND2X0_RVT U565 ( .A1(n1573), .A2(m4stg_frac[94]), .Y(n228) );
  NAND2X0_RVT U566 ( .A1(n1422), .A2(m4stg_frac[95]), .Y(n970) );
  NAND2X0_RVT U567 ( .A1(n1579), .A2(m4stg_frac[93]), .Y(n914) );
  NAND2X0_RVT U568 ( .A1(n1593), .A2(m4stg_frac[92]), .Y(n768) );
  AND4X1_RVT U569 ( .A1(n228), .A2(n970), .A3(n914), .A4(n768), .Y(n244) );
  OA222X1_RVT U570 ( .A1(n1636), .A2(n316), .A3(n35), .A4(n245), .A5(n1623), 
        .A6(n244), .Y(n446) );
  INVX1_RVT U571 ( .A(n446), .Y(n2090) );
  NAND2X0_RVT U572 ( .A1(n2043), .A2(n2090), .Y(n1757) );
  NAND2X0_RVT U573 ( .A1(n1573), .A2(m4stg_frac[86]), .Y(n827) );
  NAND2X0_RVT U574 ( .A1(n1422), .A2(m4stg_frac[87]), .Y(n918) );
  NAND2X0_RVT U575 ( .A1(n1579), .A2(m4stg_frac[85]), .Y(n965) );
  NAND2X0_RVT U576 ( .A1(n1593), .A2(m4stg_frac[84]), .Y(n824) );
  NAND4X0_RVT U577 ( .A1(n827), .A2(n918), .A3(n965), .A4(n824), .Y(n242) );
  NAND2X0_RVT U578 ( .A1(n6), .A2(n242), .Y(n230) );
  NAND2X0_RVT U579 ( .A1(n1573), .A2(m4stg_frac[74]), .Y(n819) );
  NAND2X0_RVT U580 ( .A1(n1422), .A2(m4stg_frac[75]), .Y(n952) );
  NAND2X0_RVT U581 ( .A1(n1579), .A2(m4stg_frac[73]), .Y(n955) );
  NAND2X0_RVT U582 ( .A1(n1593), .A2(m4stg_frac[72]), .Y(n781) );
  AND4X1_RVT U583 ( .A1(n819), .A2(n952), .A3(n955), .A4(n781), .Y(n298) );
  NAND2X0_RVT U584 ( .A1(n1573), .A2(m4stg_frac[82]), .Y(n822) );
  NAND2X0_RVT U585 ( .A1(n1422), .A2(m4stg_frac[83]), .Y(n963) );
  NAND2X0_RVT U586 ( .A1(n1579), .A2(m4stg_frac[81]), .Y(n959) );
  NAND2X0_RVT U587 ( .A1(n1593), .A2(m4stg_frac[80]), .Y(n814) );
  AND4X1_RVT U588 ( .A1(n822), .A2(n963), .A3(n959), .A4(n814), .Y(n306) );
  OA22X1_RVT U589 ( .A1(n298), .A2(n1623), .A3(n306), .A4(n1616), .Y(n229) );
  AND2X1_RVT U590 ( .A1(n230), .A2(n229), .Y(n233) );
  NAND2X0_RVT U591 ( .A1(n1573), .A2(m4stg_frac[78]), .Y(n815) );
  NAND2X0_RVT U592 ( .A1(n1422), .A2(m4stg_frac[79]), .Y(n961) );
  NAND2X0_RVT U593 ( .A1(n1579), .A2(m4stg_frac[77]), .Y(n951) );
  NAND2X0_RVT U594 ( .A1(n1593), .A2(m4stg_frac[76]), .Y(n818) );
  AND4X1_RVT U595 ( .A1(n815), .A2(n961), .A3(n951), .A4(n818), .Y(n305) );
  NAND2X0_RVT U596 ( .A1(n231), .A2(n1582), .Y(n232) );
  AND2X1_RVT U597 ( .A1(n233), .A2(n232), .Y(n381) );
  NAND2X0_RVT U598 ( .A1(n1573), .A2(m4stg_frac[90]), .Y(n769) );
  NAND2X0_RVT U599 ( .A1(n1422), .A2(m4stg_frac[91]), .Y(n915) );
  NAND2X0_RVT U600 ( .A1(n1579), .A2(m4stg_frac[89]), .Y(n919) );
  NAND2X0_RVT U601 ( .A1(n1593), .A2(m4stg_frac[88]), .Y(n828) );
  AND4X1_RVT U602 ( .A1(n769), .A2(n915), .A3(n919), .A4(n828), .Y(n243) );
  AO22X1_RVT U603 ( .A1(m4stg_sh_cnt[2]), .A2(n244), .A3(n1908), .A4(n243), 
        .Y(n272) );
  OA222X1_RVT U604 ( .A1(n1095), .A2(n246), .A3(n1616), .A4(n245), .A5(n272), 
        .A6(m4stg_sh_cnt[3]), .Y(n427) );
  OA22X1_RVT U605 ( .A1(n381), .A2(n437), .A3(n427), .A4(n397), .Y(n236) );
  AND2X1_RVT U606 ( .A1(n2101), .A2(n1908), .Y(n1894) );
  NAND3X0_RVT U607 ( .A1(n234), .A2(m4stg_sh_cnt[5]), .A3(n1894), .Y(n235) );
  NAND2X0_RVT U608 ( .A1(n236), .A2(n235), .Y(n2067) );
  NAND2X0_RVT U609 ( .A1(n2043), .A2(n2067), .Y(n1737) );
  NAND2X0_RVT U610 ( .A1(n1573), .A2(m4stg_frac[70]), .Y(n782) );
  NAND2X0_RVT U611 ( .A1(n1422), .A2(m4stg_frac[71]), .Y(n957) );
  NAND2X0_RVT U612 ( .A1(n1579), .A2(m4stg_frac[69]), .Y(n934) );
  NAND2X0_RVT U613 ( .A1(n1593), .A2(m4stg_frac[68]), .Y(n795) );
  NAND4X0_RVT U614 ( .A1(n782), .A2(n957), .A3(n934), .A4(n795), .Y(n268) );
  NAND2X0_RVT U615 ( .A1(n1539), .A2(n268), .Y(n238) );
  OA22X1_RVT U616 ( .A1(n305), .A2(n1616), .A3(n306), .A4(n1095), .Y(n237) );
  AND2X1_RVT U617 ( .A1(n238), .A2(n237), .Y(n241) );
  NAND2X0_RVT U618 ( .A1(n239), .A2(n1582), .Y(n240) );
  AND2X1_RVT U619 ( .A1(n241), .A2(n240), .Y(n422) );
  INVX1_RVT U620 ( .A(n242), .Y(n271) );
  AO22X1_RVT U621 ( .A1(m4stg_sh_cnt[2]), .A2(n243), .A3(n1908), .A4(n271), 
        .Y(n307) );
  OA222X1_RVT U622 ( .A1(n1095), .A2(n245), .A3(n1616), .A4(n244), .A5(n307), 
        .A6(m4stg_sh_cnt[3]), .Y(n376) );
  OAI222X1_RVT U623 ( .A1(n283), .A2(n316), .A3(n437), .A4(n422), .A5(n397), 
        .A6(n376), .Y(n2063) );
  NAND2X0_RVT U624 ( .A1(n2043), .A2(n2063), .Y(n1733) );
  OAI222X1_RVT U625 ( .A1(n35), .A2(n246), .A3(n1623), .A4(n245), .A5(n1616), 
        .A6(n284), .Y(n2094) );
  NAND2X0_RVT U626 ( .A1(n2043), .A2(n2094), .Y(n1761) );
  NAND2X0_RVT U627 ( .A1(n1539), .A2(n2102), .Y(n289) );
  NAND2X0_RVT U628 ( .A1(n1573), .A2(m4stg_frac[84]), .Y(n964) );
  NAND2X0_RVT U629 ( .A1(n1422), .A2(m4stg_frac[85]), .Y(n826) );
  NAND2X0_RVT U630 ( .A1(n1579), .A2(m4stg_frac[83]), .Y(n823) );
  NAND2X0_RVT U631 ( .A1(n1593), .A2(m4stg_frac[82]), .Y(n960) );
  NAND4X0_RVT U632 ( .A1(n964), .A2(n826), .A3(n823), .A4(n960), .Y(n274) );
  NAND2X0_RVT U633 ( .A1(n6), .A2(n274), .Y(n248) );
  NAND2X0_RVT U634 ( .A1(n1573), .A2(m4stg_frac[72]), .Y(n958) );
  NAND2X0_RVT U635 ( .A1(n1422), .A2(m4stg_frac[73]), .Y(n821) );
  NAND2X0_RVT U636 ( .A1(n1579), .A2(m4stg_frac[71]), .Y(n783) );
  NAND2X0_RVT U637 ( .A1(n1593), .A2(m4stg_frac[70]), .Y(n936) );
  AND4X1_RVT U638 ( .A1(n958), .A2(n821), .A3(n783), .A4(n936), .Y(n291) );
  NAND2X0_RVT U639 ( .A1(n1573), .A2(m4stg_frac[80]), .Y(n962) );
  NAND2X0_RVT U640 ( .A1(n1422), .A2(m4stg_frac[81]), .Y(n825) );
  NAND2X0_RVT U641 ( .A1(n1579), .A2(m4stg_frac[79]), .Y(n816) );
  NAND2X0_RVT U642 ( .A1(n1593), .A2(m4stg_frac[78]), .Y(n953) );
  AND4X1_RVT U643 ( .A1(n962), .A2(n825), .A3(n816), .A4(n953), .Y(n296) );
  OA22X1_RVT U644 ( .A1(n291), .A2(n1623), .A3(n296), .A4(n1616), .Y(n247) );
  AND2X1_RVT U645 ( .A1(n248), .A2(n247), .Y(n251) );
  NAND2X0_RVT U646 ( .A1(n1573), .A2(m4stg_frac[76]), .Y(n954) );
  NAND2X0_RVT U647 ( .A1(n1422), .A2(m4stg_frac[77]), .Y(n817) );
  NAND2X0_RVT U648 ( .A1(n1579), .A2(m4stg_frac[75]), .Y(n820) );
  NAND2X0_RVT U649 ( .A1(n1593), .A2(m4stg_frac[74]), .Y(n956) );
  AND4X1_RVT U650 ( .A1(n954), .A2(n817), .A3(n820), .A4(n956), .Y(n295) );
  NAND2X0_RVT U651 ( .A1(n249), .A2(n1582), .Y(n250) );
  AND2X1_RVT U652 ( .A1(n251), .A2(n250), .Y(n424) );
  NAND2X0_RVT U653 ( .A1(n1573), .A2(m4stg_frac[88]), .Y(n920) );
  NAND2X0_RVT U654 ( .A1(n1422), .A2(m4stg_frac[89]), .Y(n770) );
  NAND2X0_RVT U655 ( .A1(n1579), .A2(m4stg_frac[87]), .Y(n829) );
  NAND2X0_RVT U656 ( .A1(n1593), .A2(m4stg_frac[86]), .Y(n966) );
  NAND4X0_RVT U657 ( .A1(n920), .A2(n770), .A3(n829), .A4(n966), .Y(n275) );
  NAND2X0_RVT U658 ( .A1(n1539), .A2(n275), .Y(n254) );
  AOI22X1_RVT U659 ( .A1(n273), .A2(n1268), .A3(n252), .A4(n6), .Y(n253) );
  AND2X1_RVT U660 ( .A1(n254), .A2(n253), .Y(n256) );
  NAND2X0_RVT U661 ( .A1(n262), .A2(n1582), .Y(n255) );
  AND2X1_RVT U662 ( .A1(n256), .A2(n255), .Y(n378) );
  OAI222X1_RVT U663 ( .A1(n289), .A2(n257), .A3(n437), .A4(n424), .A5(n397), 
        .A6(n378), .Y(n2065) );
  NAND2X0_RVT U664 ( .A1(n2043), .A2(n2065), .Y(n1735) );
  NAND2X0_RVT U665 ( .A1(n1573), .A2(m4stg_frac[64]), .Y(n933) );
  NAND2X0_RVT U666 ( .A1(n1422), .A2(m4stg_frac[65]), .Y(n798) );
  NAND2X0_RVT U667 ( .A1(n1579), .A2(m4stg_frac[63]), .Y(n788) );
  NAND2X0_RVT U668 ( .A1(n1593), .A2(m4stg_frac[62]), .Y(n925) );
  NAND4X0_RVT U669 ( .A1(n933), .A2(n798), .A3(n788), .A4(n925), .Y(n351) );
  NAND2X0_RVT U670 ( .A1(n1539), .A2(n351), .Y(n259) );
  OA22X1_RVT U671 ( .A1(n291), .A2(n1616), .A3(n295), .A4(n1095), .Y(n258) );
  AND2X1_RVT U672 ( .A1(n259), .A2(n258), .Y(n261) );
  NAND2X0_RVT U673 ( .A1(n1573), .A2(m4stg_frac[68]), .Y(n937) );
  NAND2X0_RVT U674 ( .A1(n1422), .A2(m4stg_frac[69]), .Y(n784) );
  NAND2X0_RVT U675 ( .A1(n1579), .A2(m4stg_frac[67]), .Y(n797) );
  NAND2X0_RVT U676 ( .A1(n1593), .A2(m4stg_frac[66]), .Y(n932) );
  NAND4X0_RVT U677 ( .A1(n937), .A2(n784), .A3(n797), .A4(n932), .Y(n290) );
  NAND2X0_RVT U678 ( .A1(n290), .A2(n1582), .Y(n260) );
  AND2X1_RVT U679 ( .A1(n261), .A2(n260), .Y(n329) );
  NAND2X0_RVT U680 ( .A1(n1268), .A2(n275), .Y(n264) );
  OA22X1_RVT U681 ( .A1(n296), .A2(n1623), .A3(n276), .A4(n1095), .Y(n263) );
  AND2X1_RVT U682 ( .A1(n264), .A2(n263), .Y(n266) );
  NAND2X0_RVT U683 ( .A1(n274), .A2(n1582), .Y(n265) );
  AND2X1_RVT U684 ( .A1(n266), .A2(n265), .Y(n443) );
  INVX1_RVT U685 ( .A(n2092), .Y(n444) );
  AO222X1_RVT U686 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .A3(
        m4stg_sh_cnt[4]), .A4(n443), .A5(m4stg_sh_cnt[5]), .A6(n444), .Y(n267)
         );
  AOI21X1_RVT U687 ( .A1(n329), .A2(n2087), .A3(n267), .Y(n2057) );
  NAND2X0_RVT U688 ( .A1(n2043), .A2(n2057), .Y(n1727) );
  OA22X1_RVT U689 ( .A1(n298), .A2(n1616), .A3(n305), .A4(n1095), .Y(n270) );
  NAND2X0_RVT U690 ( .A1(n1573), .A2(m4stg_frac[66]), .Y(n796) );
  NAND2X0_RVT U691 ( .A1(n1422), .A2(m4stg_frac[67]), .Y(n935) );
  NAND2X0_RVT U692 ( .A1(n1579), .A2(m4stg_frac[65]), .Y(n930) );
  NAND2X0_RVT U693 ( .A1(n1593), .A2(m4stg_frac[64]), .Y(n785) );
  AND4X1_RVT U694 ( .A1(n796), .A2(n935), .A3(n930), .A4(n785), .Y(n319) );
  INVX1_RVT U695 ( .A(n268), .Y(n299) );
  OA22X1_RVT U696 ( .A1(n319), .A2(n1623), .A3(n299), .A4(n35), .Y(n269) );
  NAND2X0_RVT U697 ( .A1(n270), .A2(n269), .Y(n392) );
  OAI222X1_RVT U698 ( .A1(n1636), .A2(n272), .A3(n35), .A4(n271), .A5(n1623), 
        .A6(n306), .Y(n442) );
  AO222X1_RVT U699 ( .A1(n2094), .A2(n1916), .A3(n392), .A4(n2087), .A5(n442), 
        .A6(n1651), .Y(n2059) );
  NAND2X0_RVT U700 ( .A1(n2043), .A2(n2059), .Y(n1729) );
  INVX1_RVT U701 ( .A(n2096), .Y(n318) );
  OAI22X1_RVT U702 ( .A1(n1908), .A2(n275), .A3(m4stg_sh_cnt[2]), .A4(n274), 
        .Y(n297) );
  OA222X1_RVT U703 ( .A1(n1095), .A2(n277), .A3(n1616), .A4(n276), .A5(n297), 
        .A6(m4stg_sh_cnt[3]), .Y(n395) );
  NAND2X0_RVT U704 ( .A1(n1539), .A2(n290), .Y(n279) );
  OA22X1_RVT U705 ( .A1(n295), .A2(n1616), .A3(n296), .A4(n1095), .Y(n278) );
  AND2X1_RVT U706 ( .A1(n279), .A2(n278), .Y(n282) );
  NAND2X0_RVT U707 ( .A1(n280), .A2(n1582), .Y(n281) );
  AND2X1_RVT U708 ( .A1(n282), .A2(n281), .Y(n327) );
  OAI222X1_RVT U709 ( .A1(n283), .A2(n318), .A3(n397), .A4(n395), .A5(n437), 
        .A6(n327), .Y(n2061) );
  NAND2X0_RVT U710 ( .A1(n2043), .A2(n2061), .Y(n1731) );
  NAND2X0_RVT U711 ( .A1(m4stg_sh_cnt[4]), .A2(n1539), .Y(n1899) );
  OAI22X1_RVT U712 ( .A1(m4stg_sh_cnt[4]), .A2(n427), .A3(n284), .A4(n1899), 
        .Y(n2084) );
  NAND2X0_RVT U713 ( .A1(n2043), .A2(n2084), .Y(n1753) );
  OA22X1_RVT U714 ( .A1(n319), .A2(n1616), .A3(n299), .A4(n1095), .Y(n287) );
  NAND2X0_RVT U715 ( .A1(n1573), .A2(m4stg_frac[62]), .Y(n786) );
  NAND2X0_RVT U716 ( .A1(n1422), .A2(m4stg_frac[63]), .Y(n931) );
  NAND2X0_RVT U717 ( .A1(n1579), .A2(m4stg_frac[61]), .Y(n923) );
  NAND2X0_RVT U718 ( .A1(n1593), .A2(m4stg_frac[60]), .Y(n791) );
  NAND4X0_RVT U719 ( .A1(n786), .A2(n931), .A3(n923), .A4(n791), .Y(n340) );
  NAND2X0_RVT U720 ( .A1(n1573), .A2(m4stg_frac[58]), .Y(n790) );
  NAND2X0_RVT U721 ( .A1(n1422), .A2(m4stg_frac[59]), .Y(n922) );
  NAND2X0_RVT U722 ( .A1(n1579), .A2(m4stg_frac[57]), .Y(n928) );
  NAND2X0_RVT U723 ( .A1(n1593), .A2(m4stg_frac[56]), .Y(n811) );
  NAND4X0_RVT U724 ( .A1(n790), .A2(n922), .A3(n928), .A4(n811), .Y(n360) );
  OA22X1_RVT U725 ( .A1(n320), .A2(n35), .A3(n285), .A4(n1623), .Y(n286) );
  NAND2X0_RVT U726 ( .A1(n287), .A2(n286), .Y(n331) );
  AO222X1_RVT U727 ( .A1(n288), .A2(n1651), .A3(n331), .A4(n2087), .A5(n2084), 
        .A6(m4stg_sh_cnt[5]), .Y(n2051) );
  NAND2X0_RVT U728 ( .A1(n2043), .A2(n2051), .Y(n1721) );
  AO22X1_RVT U729 ( .A1(m4stg_sh_cnt[4]), .A2(n289), .A3(n1879), .A4(n378), 
        .Y(n315) );
  INVX1_RVT U730 ( .A(n315), .Y(n2082) );
  NAND2X0_RVT U731 ( .A1(n2043), .A2(n2082), .Y(n1751) );
  OA22X1_RVT U732 ( .A1(n309), .A2(n1616), .A3(n291), .A4(n1095), .Y(n294) );
  NAND2X0_RVT U733 ( .A1(n1573), .A2(m4stg_frac[60]), .Y(n924) );
  NAND2X0_RVT U734 ( .A1(n1422), .A2(m4stg_frac[61]), .Y(n787) );
  NAND2X0_RVT U735 ( .A1(n1579), .A2(m4stg_frac[59]), .Y(n792) );
  NAND2X0_RVT U736 ( .A1(n1593), .A2(m4stg_frac[58]), .Y(n929) );
  NAND4X0_RVT U737 ( .A1(n924), .A2(n787), .A3(n792), .A4(n929), .Y(n418) );
  OA22X1_RVT U738 ( .A1(n310), .A2(n35), .A3(n292), .A4(n1623), .Y(n293) );
  NAND2X0_RVT U739 ( .A1(n294), .A2(n293), .Y(n333) );
  OA222X1_RVT U740 ( .A1(n1636), .A2(n297), .A3(n35), .A4(n296), .A5(n1623), 
        .A6(n295), .Y(n384) );
  INVX1_RVT U741 ( .A(n384), .Y(n402) );
  AO222X1_RVT U742 ( .A1(n333), .A2(n2087), .A3(n2088), .A4(n1916), .A5(n402), 
        .A6(n1651), .Y(n2053) );
  NAND2X0_RVT U743 ( .A1(n2043), .A2(n2053), .Y(n1723) );
  NAND2X0_RVT U744 ( .A1(n1539), .A2(n340), .Y(n301) );
  OA22X1_RVT U745 ( .A1(n299), .A2(n1616), .A3(n298), .A4(n1095), .Y(n300) );
  AND2X1_RVT U746 ( .A1(n301), .A2(n300), .Y(n304) );
  INVX1_RVT U747 ( .A(n319), .Y(n302) );
  NAND2X0_RVT U748 ( .A1(n302), .A2(n1582), .Y(n303) );
  AND2X1_RVT U749 ( .A1(n304), .A2(n303), .Y(n328) );
  OA222X1_RVT U750 ( .A1(n1636), .A2(n307), .A3(n35), .A4(n306), .A5(n1623), 
        .A6(n305), .Y(n445) );
  AO222X1_RVT U751 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .A3(
        m4stg_sh_cnt[4]), .A4(n445), .A5(m4stg_sh_cnt[5]), .A6(n446), .Y(n308)
         );
  AOI21X1_RVT U752 ( .A1(n328), .A2(n2087), .A3(n308), .Y(n2055) );
  NAND2X0_RVT U753 ( .A1(n2043), .A2(n2055), .Y(n1725) );
  NAND2X0_RVT U754 ( .A1(n1573), .A2(m4stg_frac[56]), .Y(n927) );
  NAND2X0_RVT U755 ( .A1(n1422), .A2(m4stg_frac[57]), .Y(n789) );
  NAND2X0_RVT U756 ( .A1(n1579), .A2(m4stg_frac[55]), .Y(n810) );
  NAND2X0_RVT U757 ( .A1(n1593), .A2(m4stg_frac[54]), .Y(n947) );
  NAND4X0_RVT U758 ( .A1(n927), .A2(n789), .A3(n810), .A4(n947), .Y(n412) );
  NAND2X0_RVT U759 ( .A1(n1539), .A2(n412), .Y(n312) );
  OA22X1_RVT U760 ( .A1(n310), .A2(n1616), .A3(n309), .A4(n1095), .Y(n311) );
  AND2X1_RVT U761 ( .A1(n312), .A2(n311), .Y(n314) );
  NAND2X0_RVT U762 ( .A1(n418), .A2(n1582), .Y(n313) );
  AND2X1_RVT U763 ( .A1(n314), .A2(n313), .Y(n434) );
  OAI222X1_RVT U764 ( .A1(n315), .A2(n2069), .A3(n437), .A4(n434), .A5(n397), 
        .A6(n424), .Y(n2049) );
  NAND2X0_RVT U765 ( .A1(n2043), .A2(n2049), .Y(n1719) );
  OA22X1_RVT U766 ( .A1(m4stg_sh_cnt[4]), .A2(n376), .A3(n316), .A4(n317), .Y(
        n325) );
  INVX1_RVT U767 ( .A(n325), .Y(n2080) );
  NAND2X0_RVT U768 ( .A1(n2043), .A2(n2080), .Y(n1749) );
  OA22X1_RVT U769 ( .A1(m4stg_sh_cnt[4]), .A2(n395), .A3(n318), .A4(n317), .Y(
        n409) );
  INVX1_RVT U770 ( .A(n409), .Y(n2078) );
  NAND2X0_RVT U771 ( .A1(n2043), .A2(n2078), .Y(n1747) );
  NAND2X0_RVT U772 ( .A1(n1573), .A2(m4stg_frac[54]), .Y(n809) );
  NAND2X0_RVT U773 ( .A1(n1422), .A2(m4stg_frac[55]), .Y(n926) );
  NAND2X0_RVT U774 ( .A1(n1579), .A2(m4stg_frac[53]), .Y(n946) );
  NAND2X0_RVT U775 ( .A1(n1593), .A2(m4stg_frac[52]), .Y(n806) );
  NAND4X0_RVT U776 ( .A1(n809), .A2(n926), .A3(n946), .A4(n806), .Y(n350) );
  NAND2X0_RVT U777 ( .A1(n1539), .A2(n350), .Y(n322) );
  OA22X1_RVT U778 ( .A1(n320), .A2(n1616), .A3(n319), .A4(n1095), .Y(n321) );
  AND2X1_RVT U779 ( .A1(n322), .A2(n321), .Y(n324) );
  NAND2X0_RVT U780 ( .A1(n360), .A2(n1582), .Y(n323) );
  AND2X1_RVT U781 ( .A1(n324), .A2(n323), .Y(n432) );
  OAI222X1_RVT U782 ( .A1(n397), .A2(n422), .A3(n437), .A4(n432), .A5(n2069), 
        .A6(n325), .Y(n2047) );
  NAND2X0_RVT U783 ( .A1(n2043), .A2(n2047), .Y(n1717) );
  NAND2X0_RVT U784 ( .A1(n327), .A2(n326), .Y(n393) );
  NAND3X0_RVT U785 ( .A1(n330), .A2(n329), .A3(n328), .Y(n374) );
  AO222X1_RVT U786 ( .A1(m4stg_sh_cnt[4]), .A2(n393), .A3(m4stg_sh_cnt[4]), 
        .A4(n390), .A5(m4stg_sh_cnt[4]), .A6(n374), .Y(n456) );
  OR2X1_RVT U787 ( .A1(n373), .A2(n389), .Y(n401) );
  NOR4X1_RVT U788 ( .A1(m4stg_frac[36]), .A2(m4stg_frac[38]), .A3(
        m4stg_frac[40]), .A4(m4stg_frac[41]), .Y(n337) );
  NOR4X1_RVT U789 ( .A1(m4stg_frac[34]), .A2(m4stg_frac[33]), .A3(
        m4stg_frac[35]), .A4(m4stg_frac[37]), .Y(n336) );
  NOR4X1_RVT U790 ( .A1(m4stg_frac[30]), .A2(m4stg_frac[31]), .A3(
        m4stg_frac[32]), .A4(m4stg_frac[27]), .Y(n335) );
  NOR4X1_RVT U791 ( .A1(m4stg_frac[29]), .A2(m4stg_frac[26]), .A3(
        m4stg_frac[28]), .A4(m4stg_frac[24]), .Y(n334) );
  AND4X1_RVT U792 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .Y(n370) );
  OR4X1_RVT U793 ( .A1(m4stg_frac[49]), .A2(m4stg_frac[50]), .A3(m4stg_frac[2]), .A4(m4stg_frac[3]), .Y(n344) );
  OR4X1_RVT U794 ( .A1(m4stg_frac[44]), .A2(m4stg_frac[46]), .A3(
        m4stg_frac[48]), .A4(m4stg_frac[47]), .Y(n343) );
  OR4X1_RVT U795 ( .A1(m4stg_frac[39]), .A2(m4stg_frac[43]), .A3(
        m4stg_frac[45]), .A4(m4stg_frac[42]), .Y(n338) );
  OR4X1_RVT U796 ( .A1(n338), .A2(m4stg_frac[0]), .A3(m4stg_frac[1]), .A4(
        m4stg_frac[4]), .Y(n342) );
  AO222X1_RVT U797 ( .A1(n6), .A2(n340), .A3(n6), .A4(n360), .A5(n6), .A6(n339), .Y(n341) );
  NOR4X1_RVT U798 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .Y(n369) );
  AO22X1_RVT U799 ( .A1(n1582), .A2(n359), .A3(n1268), .A4(n417), .Y(n367) );
  AO22X1_RVT U800 ( .A1(n1582), .A2(n412), .A3(n1268), .A4(n418), .Y(n366) );
  NOR4X1_RVT U801 ( .A1(m4stg_frac[17]), .A2(m4stg_frac[16]), .A3(
        m4stg_frac[12]), .A4(m4stg_frac[14]), .Y(n348) );
  NOR4X1_RVT U802 ( .A1(m4stg_frac[13]), .A2(m4stg_frac[11]), .A3(
        m4stg_frac[9]), .A4(m4stg_frac[10]), .Y(n347) );
  NOR4X1_RVT U803 ( .A1(m4stg_frac[20]), .A2(m4stg_frac[19]), .A3(
        m4stg_frac[18]), .A4(m4stg_frac[15]), .Y(n346) );
  NOR4X1_RVT U804 ( .A1(m4stg_frac[25]), .A2(m4stg_frac[22]), .A3(
        m4stg_frac[21]), .A4(m4stg_frac[23]), .Y(n345) );
  AND4X1_RVT U805 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(n354) );
  NAND2X0_RVT U806 ( .A1(n35), .A2(n1616), .Y(n349) );
  AOI22X1_RVT U807 ( .A1(n6), .A2(n355), .A3(n350), .A4(n349), .Y(n353) );
  NAND2X0_RVT U808 ( .A1(n6), .A2(n351), .Y(n352) );
  NAND3X0_RVT U809 ( .A1(n354), .A2(n353), .A3(n352), .Y(n365) );
  HADDX1_RVT U810 ( .A0(m4stg_sh_cnt[3]), .B0(m4stg_sh_cnt[2]), .SO(n356) );
  AO22X1_RVT U811 ( .A1(m4stg_sh_cnt[3]), .A2(n357), .A3(n356), .A4(n355), .Y(
        n358) );
  AO221X1_RVT U812 ( .A1(n1268), .A2(n360), .A3(n1268), .A4(n359), .A5(n358), 
        .Y(n361) );
  AO221X1_RVT U813 ( .A1(n6), .A2(n363), .A3(n6), .A4(n362), .A5(n361), .Y(
        n364) );
  NOR4X1_RVT U814 ( .A1(n367), .A2(n366), .A3(n365), .A4(n364), .Y(n368) );
  NAND3X0_RVT U815 ( .A1(n370), .A2(n369), .A3(n368), .Y(n371) );
  AO221X1_RVT U816 ( .A1(n1651), .A2(n401), .A3(n1651), .A4(n392), .A5(n371), 
        .Y(n372) );
  AO221X1_RVT U817 ( .A1(n1916), .A2(n374), .A3(n1916), .A4(n373), .A5(n372), 
        .Y(n455) );
  INVX1_RVT U818 ( .A(n375), .Y(n430) );
  NAND4X0_RVT U819 ( .A1(n379), .A2(n378), .A3(n377), .A4(n376), .Y(n387) );
  NAND4X0_RVT U820 ( .A1(n406), .A2(n443), .A3(n380), .A4(n445), .Y(n386) );
  NAND2X0_RVT U821 ( .A1(n382), .A2(n381), .Y(n421) );
  NAND3X0_RVT U822 ( .A1(n447), .A2(n384), .A3(n383), .Y(n385) );
  AO222X1_RVT U823 ( .A1(n430), .A2(n387), .A3(n430), .A4(n386), .A5(n430), 
        .A6(n385), .Y(n388) );
  AO221X1_RVT U824 ( .A1(n1916), .A2(n390), .A3(n1916), .A4(n389), .A5(n388), 
        .Y(n454) );
  NAND4X0_RVT U825 ( .A1(n430), .A2(n395), .A3(n403), .A4(n394), .Y(n396) );
  OA22X1_RVT U826 ( .A1(n397), .A2(n420), .A3(n442), .A4(n396), .Y(n398) );
  OA221X1_RVT U827 ( .A1(m4stg_sh_cnt[4]), .A2(m4stg_sh_cnt[5]), .A3(
        m4stg_sh_cnt[4]), .A4(n400), .A5(n398), .Y(n399) );
  AOI221X1_RVT U828 ( .A1(n430), .A2(n401), .A3(n430), .A4(n400), .A5(n399), 
        .Y(n452) );
  AO22X1_RVT U829 ( .A1(m4stg_sh_cnt[4]), .A2(n2088), .A3(n1879), .A4(n402), 
        .Y(n2070) );
  AO22X1_RVT U830 ( .A1(m4stg_sh_cnt[4]), .A2(n404), .A3(n1879), .A4(n403), 
        .Y(n2038) );
  OA22X1_RVT U831 ( .A1(n1879), .A2(n2091), .A3(m4stg_sh_cnt[4]), .A4(n405), 
        .Y(n2073) );
  AO22X1_RVT U832 ( .A1(m4stg_sh_cnt[4]), .A2(n407), .A3(n1879), .A4(n406), 
        .Y(n2039) );
  NAND4X0_RVT U833 ( .A1(n409), .A2(n2038), .A3(n408), .A4(n2039), .Y(n441) );
  AOI22X1_RVT U834 ( .A1(n1573), .A2(m4stg_frac[52]), .A3(n1422), .A4(
        m4stg_frac[51]), .Y(n948) );
  NOR4X1_RVT U835 ( .A1(m4stg_frac[5]), .A2(m4stg_frac[6]), .A3(m4stg_frac[8]), 
        .A4(m4stg_frac[7]), .Y(n411) );
  NAND2X0_RVT U836 ( .A1(n1422), .A2(m4stg_frac[52]), .Y(n888) );
  AND4X1_RVT U837 ( .A1(n948), .A2(n411), .A3(n410), .A4(n888), .Y(n415) );
  AOI22X1_RVT U838 ( .A1(n1422), .A2(m4stg_frac[53]), .A3(n1579), .A4(
        m4stg_frac[51]), .Y(n414) );
  NAND2X0_RVT U839 ( .A1(n1268), .A2(n412), .Y(n413) );
  NAND3X0_RVT U840 ( .A1(n415), .A2(n414), .A3(n413), .Y(n416) );
  AO221X1_RVT U841 ( .A1(n6), .A2(n418), .A3(n6), .A4(n417), .A5(n416), .Y(
        n419) );
  AOI221X1_RVT U842 ( .A1(n1916), .A2(n421), .A3(n1916), .A4(n420), .A5(n419), 
        .Y(n439) );
  NAND4X0_RVT U843 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .Y(n431) );
  NAND3X0_RVT U844 ( .A1(n428), .A2(n427), .A3(n426), .Y(n429) );
  NAND4X0_RVT U845 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .Y(n436) );
  NAND2X0_RVT U846 ( .A1(n437), .A2(n436), .Y(n438) );
  NAND3X0_RVT U847 ( .A1(n439), .A2(n10), .A3(n438), .Y(n440) );
  OA22X1_RVT U848 ( .A1(n1879), .A2(n2094), .A3(m4stg_sh_cnt[4]), .A4(n442), 
        .Y(n2076) );
  AO22X1_RVT U849 ( .A1(m4stg_sh_cnt[4]), .A2(n444), .A3(n1879), .A4(n443), 
        .Y(n2040) );
  AO22X1_RVT U850 ( .A1(m4stg_sh_cnt[4]), .A2(n446), .A3(n1879), .A4(n445), 
        .Y(n2041) );
  AO22X1_RVT U851 ( .A1(m4stg_sh_cnt[4]), .A2(n448), .A3(n1879), .A4(n447), 
        .Y(n2042) );
  NAND4X0_RVT U852 ( .A1(n449), .A2(n2040), .A3(n2041), .A4(n2042), .Y(n450)
         );
  NAND2X0_RVT U853 ( .A1(m4stg_sh_cnt[5]), .A2(n450), .Y(n451) );
  NAND3X0_RVT U854 ( .A1(n452), .A2(n8), .A3(n451), .Y(n453) );
  OR4X1_RVT U855 ( .A1(n456), .A2(n455), .A3(n454), .A4(n453), .Y(n2045) );
  NAND2X0_RVT U856 ( .A1(n2043), .A2(n2045), .Y(n1715) );
  NAND2X0_RVT U857 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[28]), .Y(n457) );
  NAND3X0_RVT U858 ( .A1(n1), .A2(n9), .A3(n457), .Y(m2stg_frac2_array_in[29])
         );
  NAND2X0_RVT U859 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[32]), .Y(n458) );
  NAND3X0_RVT U860 ( .A1(n2), .A2(n7), .A3(n458), .Y(m2stg_frac2_array_in[30])
         );
  AOI22X1_RVT U861 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[30]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[31]), .Y(n460) );
  NAND2X0_RVT U862 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[33]), .Y(n459) );
  NAND3X0_RVT U863 ( .A1(n460), .A2(n11), .A3(n459), .Y(
        m2stg_frac2_array_in[31]) );
  AOI22X1_RVT U864 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[31]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[32]), .Y(n462) );
  NAND2X0_RVT U865 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[34]), .Y(n461) );
  NAND3X0_RVT U866 ( .A1(n462), .A2(n12), .A3(n461), .Y(
        m2stg_frac2_array_in[32]) );
  AOI22X1_RVT U867 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[32]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[33]), .Y(n464) );
  NAND2X0_RVT U868 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[35]), .Y(n463) );
  NAND3X0_RVT U869 ( .A1(n464), .A2(n13), .A3(n463), .Y(
        m2stg_frac2_array_in[33]) );
  AOI22X1_RVT U870 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[33]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[34]), .Y(n466) );
  NAND2X0_RVT U871 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[36]), .Y(n465) );
  NAND3X0_RVT U872 ( .A1(n466), .A2(n14), .A3(n465), .Y(
        m2stg_frac2_array_in[34]) );
  AOI22X1_RVT U873 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[34]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[35]), .Y(n468) );
  NAND2X0_RVT U874 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[37]), .Y(n467) );
  NAND3X0_RVT U875 ( .A1(n468), .A2(n15), .A3(n467), .Y(
        m2stg_frac2_array_in[35]) );
  AOI22X1_RVT U876 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[35]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[36]), .Y(n470) );
  NAND2X0_RVT U877 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[38]), .Y(n469) );
  NAND3X0_RVT U878 ( .A1(n470), .A2(n16), .A3(n469), .Y(
        m2stg_frac2_array_in[36]) );
  AOI22X1_RVT U879 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[36]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[37]), .Y(n472) );
  NAND2X0_RVT U880 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[39]), .Y(n471) );
  NAND3X0_RVT U881 ( .A1(n472), .A2(n17), .A3(n471), .Y(
        m2stg_frac2_array_in[37]) );
  AOI22X1_RVT U882 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[37]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[38]), .Y(n474) );
  NAND2X0_RVT U883 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[40]), .Y(n473) );
  NAND3X0_RVT U884 ( .A1(n474), .A2(n18), .A3(n473), .Y(
        m2stg_frac2_array_in[38]) );
  AOI22X1_RVT U885 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[38]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[39]), .Y(n476) );
  NAND2X0_RVT U886 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[41]), .Y(n475) );
  NAND3X0_RVT U887 ( .A1(n476), .A2(n19), .A3(n475), .Y(
        m2stg_frac2_array_in[39]) );
  AOI22X1_RVT U888 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[39]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[40]), .Y(n478) );
  NAND2X0_RVT U889 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[42]), .Y(n477) );
  NAND3X0_RVT U890 ( .A1(n478), .A2(n20), .A3(n477), .Y(
        m2stg_frac2_array_in[40]) );
  AOI22X1_RVT U891 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[40]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[41]), .Y(n480) );
  NAND2X0_RVT U892 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[43]), .Y(n479) );
  NAND3X0_RVT U893 ( .A1(n480), .A2(n21), .A3(n479), .Y(
        m2stg_frac2_array_in[41]) );
  AOI22X1_RVT U894 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[41]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[42]), .Y(n482) );
  NAND2X0_RVT U895 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[44]), .Y(n481) );
  NAND3X0_RVT U896 ( .A1(n482), .A2(n22), .A3(n481), .Y(
        m2stg_frac2_array_in[42]) );
  AOI22X1_RVT U897 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[42]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[43]), .Y(n484) );
  NAND2X0_RVT U898 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[45]), .Y(n483) );
  NAND3X0_RVT U899 ( .A1(n484), .A2(n23), .A3(n483), .Y(
        m2stg_frac2_array_in[43]) );
  AOI22X1_RVT U900 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[43]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[44]), .Y(n486) );
  NAND2X0_RVT U901 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[46]), .Y(n485) );
  NAND3X0_RVT U902 ( .A1(n486), .A2(n24), .A3(n485), .Y(
        m2stg_frac2_array_in[44]) );
  AOI22X1_RVT U903 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[44]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[45]), .Y(n488) );
  NAND2X0_RVT U904 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[47]), .Y(n487) );
  NAND3X0_RVT U905 ( .A1(n488), .A2(n25), .A3(n487), .Y(
        m2stg_frac2_array_in[45]) );
  AOI22X1_RVT U906 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[45]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[46]), .Y(n491) );
  AOI22X1_RVT U907 ( .A1(mul_frac_in2[49]), .A2(m2stg_frac2_sng_norm), .A3(
        m2stg_frac2_inf), .A4(m1stg_inf_zero_in), .Y(n490) );
  NAND2X0_RVT U908 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[48]), .Y(n489) );
  NAND3X0_RVT U909 ( .A1(n491), .A2(n490), .A3(n489), .Y(
        m2stg_frac2_array_in[46]) );
  AOI22X1_RVT U910 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[46]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[47]), .Y(n493) );
  NAND2X0_RVT U911 ( .A1(mul_frac_in2[49]), .A2(m2stg_frac2_sng_dnrm), .Y(n492) );
  NAND3X0_RVT U912 ( .A1(n493), .A2(n26), .A3(n492), .Y(
        m2stg_frac2_array_in[47]) );
  AOI22X1_RVT U913 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[47]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[48]), .Y(n495) );
  NAND2X0_RVT U914 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[50]), .Y(n494) );
  NAND3X0_RVT U915 ( .A1(n495), .A2(n27), .A3(n494), .Y(
        m2stg_frac2_array_in[48]) );
  AOI22X1_RVT U916 ( .A1(mul_frac_in2[49]), .A2(m2stg_frac2_dbl_norm), .A3(
        m2stg_frac2_dbl_dnrm), .A4(mul_frac_in2[48]), .Y(n497) );
  NAND2X0_RVT U917 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[51]), .Y(n496) );
  NAND3X0_RVT U918 ( .A1(n497), .A2(n28), .A3(n496), .Y(
        m2stg_frac2_array_in[49]) );
  NAND2X0_RVT U919 ( .A1(mul_frac_in2[49]), .A2(m2stg_frac2_dbl_dnrm), .Y(n498) );
  NAND3X0_RVT U920 ( .A1(n29), .A2(n3), .A3(n498), .Y(m2stg_frac2_array_in[50]) );
  NAND4X0_RVT U921 ( .A1(m5stg_frac_pre2[20]), .A2(m5stg_frac_pre1[20]), .A3(
        m5stg_frac_pre4[20]), .A4(m5stg_frac_pre3[20]), .Y(m5stg_frac_32_0[20]) );
  AND4X1_RVT U922 ( .A1(m5stg_frac_pre2[19]), .A2(m5stg_frac_pre1[19]), .A3(
        m5stg_frac_pre4[19]), .A4(m5stg_frac_pre3[19]), .Y(n1504) );
  NAND3X0_RVT U923 ( .A1(m5stg_fmulda), .A2(\add_x_3/A[1] ), .A3(
        \add_x_3/A[0] ), .Y(n758) );
  INVX1_RVT U924 ( .A(n758), .Y(n754) );
  NAND3X0_RVT U925 ( .A1(n754), .A2(\add_x_3/A[2] ), .A3(\add_x_3/A[3] ), .Y(
        n752) );
  INVX1_RVT U926 ( .A(n752), .Y(n748) );
  NAND3X0_RVT U927 ( .A1(n748), .A2(\add_x_3/A[4] ), .A3(\add_x_3/A[5] ), .Y(
        n746) );
  INVX1_RVT U928 ( .A(n746), .Y(n742) );
  NAND3X0_RVT U929 ( .A1(n742), .A2(\add_x_3/A[6] ), .A3(\add_x_3/A[7] ), .Y(
        n740) );
  INVX1_RVT U930 ( .A(n740), .Y(n736) );
  NAND3X0_RVT U931 ( .A1(n736), .A2(\add_x_3/A[8] ), .A3(\add_x_3/A[9] ), .Y(
        n734) );
  INVX1_RVT U932 ( .A(n734), .Y(n730) );
  NAND3X0_RVT U933 ( .A1(n730), .A2(\add_x_3/A[10] ), .A3(\add_x_3/A[11] ), 
        .Y(n723) );
  INVX1_RVT U934 ( .A(n723), .Y(n726) );
  NAND3X0_RVT U935 ( .A1(n726), .A2(\add_x_3/A[12] ), .A3(\add_x_3/A[13] ), 
        .Y(n716) );
  INVX1_RVT U936 ( .A(n716), .Y(n499) );
  NAND3X0_RVT U937 ( .A1(n499), .A2(\add_x_3/A[14] ), .A3(\add_x_3/A[15] ), 
        .Y(n708) );
  INVX1_RVT U938 ( .A(n708), .Y(n711) );
  NAND4X0_RVT U939 ( .A1(m5stg_frac_pre2[19]), .A2(m5stg_frac_pre1[19]), .A3(
        m5stg_frac_pre4[19]), .A4(m5stg_frac_pre3[19]), .Y(m5stg_frac_32_0[19]) );
  NAND3X0_RVT U940 ( .A1(n711), .A2(m5stg_frac_32_0[19]), .A3(
        m5stg_frac_32_0[20]), .Y(n700) );
  INVX1_RVT U941 ( .A(n700), .Y(n703) );
  NAND3X0_RVT U942 ( .A1(n703), .A2(\add_x_3/A[18] ), .A3(\add_x_3/A[19] ), 
        .Y(n692) );
  INVX1_RVT U943 ( .A(n692), .Y(n695) );
  NAND3X0_RVT U944 ( .A1(n695), .A2(\add_x_3/A[20] ), .A3(\add_x_3/A[21] ), 
        .Y(n684) );
  INVX1_RVT U945 ( .A(n684), .Y(n687) );
  AND3X1_RVT U946 ( .A1(n687), .A2(\add_x_3/A[22] ), .A3(\add_x_3/A[23] ), .Y(
        n679) );
  AND3X1_RVT U947 ( .A1(n679), .A2(\add_x_3/A[24] ), .A3(\add_x_3/A[25] ), .Y(
        n671) );
  AND4X1_RVT U948 ( .A1(n671), .A2(\add_x_3/A[28] ), .A3(\add_x_3/A[26] ), 
        .A4(\add_x_3/A[27] ), .Y(n661) );
  AO222X1_RVT U949 ( .A1(m5stg_fmuls), .A2(n661), .A3(m5stg_fmuls), .A4(
        \add_x_3/A[29] ), .A5(n661), .A6(\add_x_3/A[29] ), .Y(n653) );
  NAND4X0_RVT U950 ( .A1(m5stg_frac_pre2[33]), .A2(m5stg_frac_pre1[33]), .A3(
        m5stg_frac_pre4[33]), .A4(m5stg_frac_pre3[33]), .Y(n655) );
  NAND4X0_RVT U951 ( .A1(m5stg_frac_pre2[34]), .A2(m5stg_frac_pre1[34]), .A3(
        m5stg_frac_pre4[34]), .A4(m5stg_frac_pre3[34]), .Y(n650) );
  NAND3X0_RVT U952 ( .A1(n653), .A2(n655), .A3(n650), .Y(n640) );
  INVX1_RVT U953 ( .A(n640), .Y(n644) );
  NAND4X0_RVT U954 ( .A1(m5stg_frac_pre2[35]), .A2(m5stg_frac_pre1[35]), .A3(
        m5stg_frac_pre4[35]), .A4(m5stg_frac_pre3[35]), .Y(n646) );
  NAND4X0_RVT U955 ( .A1(m5stg_frac_pre2[36]), .A2(m5stg_frac_pre1[36]), .A3(
        m5stg_frac_pre4[36]), .A4(m5stg_frac_pre3[36]), .Y(n641) );
  NAND3X0_RVT U956 ( .A1(n644), .A2(n646), .A3(n641), .Y(n630) );
  INVX1_RVT U957 ( .A(n630), .Y(n634) );
  NAND4X0_RVT U958 ( .A1(m5stg_frac_pre2[37]), .A2(m5stg_frac_pre1[37]), .A3(
        m5stg_frac_pre4[37]), .A4(m5stg_frac_pre3[37]), .Y(n636) );
  NAND4X0_RVT U959 ( .A1(m5stg_frac_pre2[38]), .A2(m5stg_frac_pre1[38]), .A3(
        m5stg_frac_pre4[38]), .A4(m5stg_frac_pre3[38]), .Y(n631) );
  NAND3X0_RVT U960 ( .A1(n634), .A2(n636), .A3(n631), .Y(n620) );
  INVX1_RVT U961 ( .A(n620), .Y(n624) );
  NAND4X0_RVT U962 ( .A1(m5stg_frac_pre2[39]), .A2(m5stg_frac_pre1[39]), .A3(
        m5stg_frac_pre4[39]), .A4(m5stg_frac_pre3[39]), .Y(n626) );
  NAND4X0_RVT U963 ( .A1(m5stg_frac_pre2[40]), .A2(m5stg_frac_pre1[40]), .A3(
        m5stg_frac_pre4[40]), .A4(m5stg_frac_pre3[40]), .Y(n621) );
  NAND3X0_RVT U964 ( .A1(n624), .A2(n626), .A3(n621), .Y(n610) );
  INVX1_RVT U965 ( .A(n610), .Y(n614) );
  NAND4X0_RVT U966 ( .A1(m5stg_frac_pre2[41]), .A2(m5stg_frac_pre1[41]), .A3(
        m5stg_frac_pre4[41]), .A4(m5stg_frac_pre3[41]), .Y(n616) );
  NAND4X0_RVT U967 ( .A1(m5stg_frac_pre2[42]), .A2(m5stg_frac_pre1[42]), .A3(
        m5stg_frac_pre4[42]), .A4(m5stg_frac_pre3[42]), .Y(n611) );
  NAND3X0_RVT U968 ( .A1(n614), .A2(n616), .A3(n611), .Y(n600) );
  INVX1_RVT U969 ( .A(n600), .Y(n604) );
  NAND4X0_RVT U970 ( .A1(m5stg_frac_pre2[43]), .A2(m5stg_frac_pre1[43]), .A3(
        m5stg_frac_pre4[43]), .A4(m5stg_frac_pre3[43]), .Y(n606) );
  NAND4X0_RVT U971 ( .A1(m5stg_frac_pre2[44]), .A2(m5stg_frac_pre1[44]), .A3(
        m5stg_frac_pre4[44]), .A4(m5stg_frac_pre3[44]), .Y(n601) );
  NAND3X0_RVT U972 ( .A1(n604), .A2(n606), .A3(n601), .Y(n590) );
  INVX1_RVT U973 ( .A(n590), .Y(n594) );
  NAND4X0_RVT U974 ( .A1(m5stg_frac_pre2[45]), .A2(m5stg_frac_pre1[45]), .A3(
        m5stg_frac_pre4[45]), .A4(m5stg_frac_pre3[45]), .Y(n596) );
  NAND4X0_RVT U975 ( .A1(m5stg_frac_pre2[46]), .A2(m5stg_frac_pre1[46]), .A3(
        m5stg_frac_pre4[46]), .A4(m5stg_frac_pre3[46]), .Y(n591) );
  NAND3X0_RVT U976 ( .A1(n594), .A2(n596), .A3(n591), .Y(n580) );
  INVX1_RVT U977 ( .A(n580), .Y(n584) );
  NAND4X0_RVT U978 ( .A1(m5stg_frac_pre2[47]), .A2(m5stg_frac_pre1[47]), .A3(
        m5stg_frac_pre4[47]), .A4(m5stg_frac_pre3[47]), .Y(n586) );
  NAND4X0_RVT U979 ( .A1(m5stg_frac_pre2[48]), .A2(m5stg_frac_pre1[48]), .A3(
        m5stg_frac_pre4[48]), .A4(m5stg_frac_pre3[48]), .Y(n581) );
  NAND3X0_RVT U980 ( .A1(n584), .A2(n586), .A3(n581), .Y(n570) );
  INVX1_RVT U981 ( .A(n570), .Y(n574) );
  NAND4X0_RVT U982 ( .A1(m5stg_frac_pre2[49]), .A2(m5stg_frac_pre1[49]), .A3(
        m5stg_frac_pre4[49]), .A4(m5stg_frac_pre3[49]), .Y(n576) );
  NAND4X0_RVT U983 ( .A1(m5stg_frac_pre2[50]), .A2(m5stg_frac_pre1[50]), .A3(
        m5stg_frac_pre4[50]), .A4(m5stg_frac_pre3[50]), .Y(n571) );
  NAND3X0_RVT U984 ( .A1(n574), .A2(n576), .A3(n571), .Y(n560) );
  INVX1_RVT U985 ( .A(n560), .Y(n564) );
  NAND4X0_RVT U986 ( .A1(m5stg_frac_pre2[51]), .A2(m5stg_frac_pre1[51]), .A3(
        m5stg_frac_pre4[51]), .A4(m5stg_frac_pre3[51]), .Y(n566) );
  NAND4X0_RVT U987 ( .A1(m5stg_frac_pre2[52]), .A2(m5stg_frac_pre1[52]), .A3(
        m5stg_frac_pre4[52]), .A4(m5stg_frac_pre3[52]), .Y(n561) );
  NAND3X0_RVT U988 ( .A1(n564), .A2(n566), .A3(n561), .Y(n557) );
  INVX1_RVT U989 ( .A(n557), .Y(n551) );
  NAND4X0_RVT U990 ( .A1(m5stg_frac_pre2[53]), .A2(m5stg_frac_pre1[53]), .A3(
        m5stg_frac_pre4[53]), .A4(m5stg_frac_pre3[53]), .Y(n555) );
  NAND4X0_RVT U991 ( .A1(m5stg_frac_pre2[54]), .A2(m5stg_frac_pre1[54]), .A3(
        m5stg_frac_pre4[54]), .A4(m5stg_frac_pre3[54]), .Y(n836) );
  AND3X1_RVT U992 ( .A1(n551), .A2(n555), .A3(n836), .Y(m5stg_fracadd_cout) );
  AO22X1_RVT U995 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[51]), .A3(
        m2stg_frac2_sng_dnrm), .A4(mul_frac_in2[54]), .Y(n502) );
  OR4X1_RVT U996 ( .A1(n502), .A2(m2stg_frac2_sng_norm), .A3(m2stg_frac2_inf), 
        .A4(m2stg_frac2_dbl_norm), .Y(m2stg_frac2_array_in[52]) );
  OR2X1_RVT U997 ( .A1(mul_frac_in2[54]), .A2(m1stg_snan_sng_in2), .Y(n503) );
  NAND2X0_RVT U998 ( .A1(m2stg_frac2_sng_dnrm), .A2(mul_frac_in2[53]), .Y(n504) );
  NAND3X0_RVT U999 ( .A1(n4), .A2(n9), .A3(n504), .Y(n505) );
  AO221X1_RVT U1000 ( .A1(m2stg_frac2_dbl_norm), .A2(mul_frac_in2[51]), .A3(
        m2stg_frac2_dbl_norm), .A4(m1stg_snan_dbl_in2), .A5(n505), .Y(
        m2stg_frac2_array_in[51]) );
  AOI22X1_RVT U1001 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[27]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[28]), .Y(n506) );
  NAND2X0_RVT U1002 ( .A1(m2stg_frac2_inf), .A2(m1stg_inf_zero_in_dbl), .Y(
        n509) );
  NAND2X0_RVT U1003 ( .A1(n506), .A2(n509), .Y(m2stg_frac2_array_in[28]) );
  AOI22X1_RVT U1004 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[26]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[27]), .Y(n507) );
  NAND2X0_RVT U1005 ( .A1(n507), .A2(n509), .Y(m2stg_frac2_array_in[27]) );
  AOI22X1_RVT U1006 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[25]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[26]), .Y(n508) );
  NAND2X0_RVT U1007 ( .A1(n508), .A2(n509), .Y(m2stg_frac2_array_in[26]) );
  AOI22X1_RVT U1008 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[24]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[25]), .Y(n510) );
  NAND2X0_RVT U1009 ( .A1(n510), .A2(n509), .Y(m2stg_frac2_array_in[25]) );
  AOI22X1_RVT U1010 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[23]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[24]), .Y(n511) );
  NAND2X0_RVT U1011 ( .A1(n511), .A2(n509), .Y(m2stg_frac2_array_in[24]) );
  AOI22X1_RVT U1012 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[22]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[23]), .Y(n512) );
  NAND2X0_RVT U1013 ( .A1(n512), .A2(n509), .Y(m2stg_frac2_array_in[23]) );
  AOI22X1_RVT U1014 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[21]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[22]), .Y(n513) );
  NAND2X0_RVT U1015 ( .A1(n513), .A2(n509), .Y(m2stg_frac2_array_in[22]) );
  AOI22X1_RVT U1016 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[20]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[21]), .Y(n514) );
  NAND2X0_RVT U1017 ( .A1(n514), .A2(n509), .Y(m2stg_frac2_array_in[21]) );
  AOI22X1_RVT U1018 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[19]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[20]), .Y(n515) );
  NAND2X0_RVT U1019 ( .A1(n515), .A2(n509), .Y(m2stg_frac2_array_in[20]) );
  AOI22X1_RVT U1020 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[18]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[19]), .Y(n516) );
  NAND2X0_RVT U1021 ( .A1(n516), .A2(n509), .Y(m2stg_frac2_array_in[19]) );
  AOI22X1_RVT U1022 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[17]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[18]), .Y(n517) );
  NAND2X0_RVT U1023 ( .A1(n517), .A2(n509), .Y(m2stg_frac2_array_in[18]) );
  AOI22X1_RVT U1024 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[16]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[17]), .Y(n518) );
  NAND2X0_RVT U1025 ( .A1(n518), .A2(n509), .Y(m2stg_frac2_array_in[17]) );
  AOI22X1_RVT U1026 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[15]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[16]), .Y(n519) );
  NAND2X0_RVT U1027 ( .A1(n519), .A2(n509), .Y(m2stg_frac2_array_in[16]) );
  AOI22X1_RVT U1028 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[14]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[15]), .Y(n520) );
  NAND2X0_RVT U1029 ( .A1(n520), .A2(n509), .Y(m2stg_frac2_array_in[15]) );
  AOI22X1_RVT U1030 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[13]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[14]), .Y(n521) );
  NAND2X0_RVT U1031 ( .A1(n521), .A2(n509), .Y(m2stg_frac2_array_in[14]) );
  AOI22X1_RVT U1032 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[12]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[13]), .Y(n522) );
  NAND2X0_RVT U1033 ( .A1(n522), .A2(n509), .Y(m2stg_frac2_array_in[13]) );
  AOI22X1_RVT U1034 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[11]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[12]), .Y(n523) );
  NAND2X0_RVT U1035 ( .A1(n523), .A2(n509), .Y(m2stg_frac2_array_in[12]) );
  AOI22X1_RVT U1036 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[10]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[11]), .Y(n524) );
  NAND2X0_RVT U1037 ( .A1(n524), .A2(n509), .Y(m2stg_frac2_array_in[11]) );
  AOI22X1_RVT U1038 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[9]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[10]), .Y(n525) );
  NAND2X0_RVT U1039 ( .A1(n525), .A2(n509), .Y(m2stg_frac2_array_in[10]) );
  AOI22X1_RVT U1040 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[8]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[9]), .Y(n526) );
  NAND2X0_RVT U1041 ( .A1(n526), .A2(n509), .Y(m2stg_frac2_array_in[9]) );
  AOI22X1_RVT U1042 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[7]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[8]), .Y(n527) );
  NAND2X0_RVT U1043 ( .A1(n527), .A2(n509), .Y(m2stg_frac2_array_in[8]) );
  AOI22X1_RVT U1044 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[6]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[7]), .Y(n528) );
  NAND2X0_RVT U1045 ( .A1(n528), .A2(n509), .Y(m2stg_frac2_array_in[7]) );
  AOI22X1_RVT U1046 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[5]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[6]), .Y(n529) );
  NAND2X0_RVT U1047 ( .A1(n529), .A2(n509), .Y(m2stg_frac2_array_in[6]) );
  AOI22X1_RVT U1048 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[4]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[5]), .Y(n530) );
  NAND2X0_RVT U1049 ( .A1(n530), .A2(n509), .Y(m2stg_frac2_array_in[5]) );
  AOI22X1_RVT U1050 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[3]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[4]), .Y(n531) );
  NAND2X0_RVT U1051 ( .A1(n531), .A2(n509), .Y(m2stg_frac2_array_in[4]) );
  AOI22X1_RVT U1052 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[2]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[3]), .Y(n532) );
  NAND2X0_RVT U1053 ( .A1(n532), .A2(n509), .Y(m2stg_frac2_array_in[3]) );
  AOI22X1_RVT U1054 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[1]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[2]), .Y(n533) );
  NAND2X0_RVT U1055 ( .A1(n533), .A2(n509), .Y(m2stg_frac2_array_in[2]) );
  AOI22X1_RVT U1056 ( .A1(m2stg_frac2_dbl_dnrm), .A2(mul_frac_in2[0]), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[1]), .Y(n534) );
  NAND2X0_RVT U1057 ( .A1(n534), .A2(n509), .Y(m2stg_frac2_array_in[1]) );
  AO22X1_RVT U1058 ( .A1(m2stg_frac2_inf), .A2(m1stg_inf_zero_in_dbl), .A3(
        m2stg_frac2_dbl_norm), .A4(mul_frac_in2[0]), .Y(
        m2stg_frac2_array_in[0]) );
  AO22X1_RVT U1059 ( .A1(mul_frac_in1[51]), .A2(m1stg_dblop), .A3(
        mul_frac_in1[54]), .A4(m1stg_dblop_inv), .Y(m1stg_ld0_1_din[52]) );
  AO22X1_RVT U1060 ( .A1(mul_frac_in1[50]), .A2(m1stg_dblop), .A3(
        mul_frac_in1[53]), .A4(m1stg_dblop_inv), .Y(m1stg_ld0_1_din[51]) );
  AO22X1_RVT U1061 ( .A1(mul_frac_in1[52]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[49]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[50]) );
  AO22X1_RVT U1062 ( .A1(mul_frac_in1[51]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[48]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[49]) );
  AO22X1_RVT U1063 ( .A1(mul_frac_in1[50]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[47]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[48]) );
  AO22X1_RVT U1064 ( .A1(mul_frac_in1[49]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[46]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[47]) );
  AO22X1_RVT U1065 ( .A1(mul_frac_in1[48]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[45]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[46]) );
  AO22X1_RVT U1066 ( .A1(mul_frac_in1[47]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[44]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[45]) );
  AO22X1_RVT U1067 ( .A1(mul_frac_in1[46]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[43]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[44]) );
  AO22X1_RVT U1068 ( .A1(mul_frac_in1[45]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[42]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[43]) );
  AO22X1_RVT U1069 ( .A1(mul_frac_in1[44]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[41]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[42]) );
  AO22X1_RVT U1070 ( .A1(mul_frac_in1[43]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[40]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[41]) );
  AO22X1_RVT U1071 ( .A1(mul_frac_in1[42]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[39]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[40]) );
  AO22X1_RVT U1072 ( .A1(mul_frac_in1[41]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[38]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[39]) );
  AO22X1_RVT U1073 ( .A1(mul_frac_in1[40]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[37]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[38]) );
  AO22X1_RVT U1074 ( .A1(mul_frac_in1[39]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[36]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[37]) );
  AO22X1_RVT U1075 ( .A1(mul_frac_in1[38]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[35]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[36]) );
  AO22X1_RVT U1076 ( .A1(mul_frac_in1[37]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[34]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[35]) );
  AO22X1_RVT U1077 ( .A1(mul_frac_in1[36]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[33]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[34]) );
  AO22X1_RVT U1078 ( .A1(mul_frac_in1[35]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[32]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[33]) );
  AO22X1_RVT U1079 ( .A1(mul_frac_in1[34]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[31]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[32]) );
  AO22X1_RVT U1080 ( .A1(mul_frac_in1[33]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[30]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[31]) );
  AO22X1_RVT U1081 ( .A1(mul_frac_in1[32]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in1[29]), .A4(m1stg_dblop), .Y(m1stg_ld0_1_din[30]) );
  AND2X1_RVT U1082 ( .A1(mul_frac_in1[28]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_1_din[29]) );
  AND2X1_RVT U1083 ( .A1(m1stg_dblop), .A2(mul_frac_in1[27]), .Y(
        m1stg_ld0_1_din[28]) );
  AND2X1_RVT U1084 ( .A1(m1stg_dblop), .A2(mul_frac_in1[26]), .Y(
        m1stg_ld0_1_din[27]) );
  AND2X1_RVT U1085 ( .A1(m1stg_dblop), .A2(mul_frac_in1[25]), .Y(
        m1stg_ld0_1_din[26]) );
  AND2X1_RVT U1086 ( .A1(m1stg_dblop), .A2(mul_frac_in1[24]), .Y(
        m1stg_ld0_1_din[25]) );
  AND2X1_RVT U1087 ( .A1(m1stg_dblop), .A2(mul_frac_in1[23]), .Y(
        m1stg_ld0_1_din[24]) );
  AND2X1_RVT U1088 ( .A1(m1stg_dblop), .A2(mul_frac_in1[22]), .Y(
        m1stg_ld0_1_din[23]) );
  AND2X1_RVT U1089 ( .A1(m1stg_dblop), .A2(mul_frac_in1[21]), .Y(
        m1stg_ld0_1_din[22]) );
  AND2X1_RVT U1090 ( .A1(m1stg_dblop), .A2(mul_frac_in1[20]), .Y(
        m1stg_ld0_1_din[21]) );
  AND2X1_RVT U1091 ( .A1(m1stg_dblop), .A2(mul_frac_in1[19]), .Y(
        m1stg_ld0_1_din[20]) );
  AND2X1_RVT U1092 ( .A1(m1stg_dblop), .A2(mul_frac_in1[18]), .Y(
        m1stg_ld0_1_din[19]) );
  AND2X1_RVT U1093 ( .A1(m1stg_dblop), .A2(mul_frac_in1[17]), .Y(
        m1stg_ld0_1_din[18]) );
  AND2X1_RVT U1094 ( .A1(m1stg_dblop), .A2(mul_frac_in1[16]), .Y(
        m1stg_ld0_1_din[17]) );
  AND2X1_RVT U1095 ( .A1(m1stg_dblop), .A2(mul_frac_in1[15]), .Y(
        m1stg_ld0_1_din[16]) );
  AND2X1_RVT U1096 ( .A1(m1stg_dblop), .A2(mul_frac_in1[14]), .Y(
        m1stg_ld0_1_din[15]) );
  AND2X1_RVT U1097 ( .A1(m1stg_dblop), .A2(mul_frac_in1[13]), .Y(
        m1stg_ld0_1_din[14]) );
  AND2X1_RVT U1098 ( .A1(m1stg_dblop), .A2(mul_frac_in1[12]), .Y(
        m1stg_ld0_1_din[13]) );
  AND2X1_RVT U1099 ( .A1(m1stg_dblop), .A2(mul_frac_in1[11]), .Y(
        m1stg_ld0_1_din[12]) );
  AND2X1_RVT U1100 ( .A1(m1stg_dblop), .A2(mul_frac_in1[10]), .Y(
        m1stg_ld0_1_din[11]) );
  AND2X1_RVT U1101 ( .A1(m1stg_dblop), .A2(mul_frac_in1[9]), .Y(
        m1stg_ld0_1_din[10]) );
  AND2X1_RVT U1102 ( .A1(m1stg_dblop), .A2(mul_frac_in1[8]), .Y(
        m1stg_ld0_1_din[9]) );
  AND2X1_RVT U1103 ( .A1(m1stg_dblop), .A2(mul_frac_in1[7]), .Y(
        m1stg_ld0_1_din[8]) );
  AND2X1_RVT U1104 ( .A1(m1stg_dblop), .A2(mul_frac_in1[6]), .Y(
        m1stg_ld0_1_din[7]) );
  AND2X1_RVT U1105 ( .A1(m1stg_dblop), .A2(mul_frac_in1[5]), .Y(
        m1stg_ld0_1_din[6]) );
  AND2X1_RVT U1106 ( .A1(m1stg_dblop), .A2(mul_frac_in1[4]), .Y(
        m1stg_ld0_1_din[5]) );
  AND2X1_RVT U1107 ( .A1(m1stg_dblop), .A2(mul_frac_in1[3]), .Y(
        m1stg_ld0_1_din[4]) );
  AND2X1_RVT U1108 ( .A1(m1stg_dblop), .A2(mul_frac_in1[2]), .Y(
        m1stg_ld0_1_din[3]) );
  AND2X1_RVT U1109 ( .A1(m1stg_dblop), .A2(mul_frac_in1[1]), .Y(
        m1stg_ld0_1_din[2]) );
  AND2X1_RVT U1110 ( .A1(m1stg_dblop), .A2(mul_frac_in1[0]), .Y(
        m1stg_ld0_1_din[1]) );
  AO22X1_RVT U1111 ( .A1(mul_frac_in2[51]), .A2(m1stg_dblop), .A3(
        mul_frac_in2[54]), .A4(m1stg_dblop_inv), .Y(m1stg_ld0_2_din[52]) );
  AO22X1_RVT U1112 ( .A1(mul_frac_in2[53]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[50]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[51]) );
  AO22X1_RVT U1113 ( .A1(mul_frac_in2[49]), .A2(m1stg_dblop), .A3(
        mul_frac_in2[52]), .A4(m1stg_dblop_inv), .Y(m1stg_ld0_2_din[50]) );
  AO22X1_RVT U1114 ( .A1(mul_frac_in2[51]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[48]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[49]) );
  AO22X1_RVT U1115 ( .A1(mul_frac_in2[50]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[47]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[48]) );
  AO22X1_RVT U1116 ( .A1(mul_frac_in2[49]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[46]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[47]) );
  AO22X1_RVT U1117 ( .A1(mul_frac_in2[48]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[45]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[46]) );
  AO22X1_RVT U1118 ( .A1(mul_frac_in2[47]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[44]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[45]) );
  AO22X1_RVT U1119 ( .A1(mul_frac_in2[46]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[43]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[44]) );
  AO22X1_RVT U1120 ( .A1(mul_frac_in2[45]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[42]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[43]) );
  AO22X1_RVT U1121 ( .A1(mul_frac_in2[44]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[41]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[42]) );
  AO22X1_RVT U1122 ( .A1(mul_frac_in2[43]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[40]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[41]) );
  AO22X1_RVT U1123 ( .A1(mul_frac_in2[42]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[39]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[40]) );
  AO22X1_RVT U1124 ( .A1(mul_frac_in2[41]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[38]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[39]) );
  AO22X1_RVT U1125 ( .A1(mul_frac_in2[40]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[37]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[38]) );
  AO22X1_RVT U1126 ( .A1(mul_frac_in2[39]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[36]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[37]) );
  AO22X1_RVT U1127 ( .A1(mul_frac_in2[38]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[35]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[36]) );
  AO22X1_RVT U1128 ( .A1(mul_frac_in2[37]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[34]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[35]) );
  AO22X1_RVT U1129 ( .A1(mul_frac_in2[36]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[33]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[34]) );
  AO22X1_RVT U1130 ( .A1(mul_frac_in2[35]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[32]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[33]) );
  AO22X1_RVT U1131 ( .A1(mul_frac_in2[34]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[31]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[32]) );
  AO22X1_RVT U1132 ( .A1(mul_frac_in2[33]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[30]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[31]) );
  AO22X1_RVT U1133 ( .A1(mul_frac_in2[32]), .A2(m1stg_dblop_inv), .A3(
        mul_frac_in2[29]), .A4(m1stg_dblop), .Y(m1stg_ld0_2_din[30]) );
  AND2X1_RVT U1134 ( .A1(mul_frac_in2[28]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[29]) );
  AND2X1_RVT U1135 ( .A1(mul_frac_in2[27]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[28]) );
  AND2X1_RVT U1136 ( .A1(mul_frac_in2[26]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[27]) );
  AND2X1_RVT U1137 ( .A1(mul_frac_in2[25]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[26]) );
  AND2X1_RVT U1138 ( .A1(mul_frac_in2[24]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[25]) );
  AND2X1_RVT U1139 ( .A1(mul_frac_in2[23]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[24]) );
  AND2X1_RVT U1140 ( .A1(mul_frac_in2[22]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[23]) );
  AND2X1_RVT U1141 ( .A1(mul_frac_in2[21]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[22]) );
  AND2X1_RVT U1142 ( .A1(mul_frac_in2[20]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[21]) );
  AND2X1_RVT U1143 ( .A1(mul_frac_in2[19]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[20]) );
  AND2X1_RVT U1144 ( .A1(mul_frac_in2[18]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[19]) );
  AND2X1_RVT U1145 ( .A1(mul_frac_in2[17]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[18]) );
  AND2X1_RVT U1146 ( .A1(mul_frac_in2[16]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[17]) );
  AND2X1_RVT U1147 ( .A1(mul_frac_in2[15]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[16]) );
  AND2X1_RVT U1148 ( .A1(mul_frac_in2[14]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[15]) );
  AND2X1_RVT U1149 ( .A1(mul_frac_in2[13]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[14]) );
  AND2X1_RVT U1150 ( .A1(mul_frac_in2[12]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[13]) );
  AND2X1_RVT U1151 ( .A1(mul_frac_in2[11]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[12]) );
  AND2X1_RVT U1152 ( .A1(mul_frac_in2[10]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[11]) );
  AND2X1_RVT U1153 ( .A1(mul_frac_in2[9]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[10]) );
  AND2X1_RVT U1154 ( .A1(mul_frac_in2[8]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[9]) );
  AND2X1_RVT U1155 ( .A1(mul_frac_in2[7]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[8]) );
  AND2X1_RVT U1156 ( .A1(mul_frac_in2[6]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[7]) );
  AND2X1_RVT U1157 ( .A1(mul_frac_in2[5]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[6]) );
  AND2X1_RVT U1158 ( .A1(mul_frac_in2[4]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[5]) );
  AND2X1_RVT U1159 ( .A1(mul_frac_in2[3]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[4]) );
  AND2X1_RVT U1160 ( .A1(mul_frac_in2[2]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[3]) );
  AND2X1_RVT U1161 ( .A1(mul_frac_in2[1]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[2]) );
  AND2X1_RVT U1162 ( .A1(mul_frac_in2[0]), .A2(m1stg_dblop), .Y(
        m1stg_ld0_2_din[1]) );
  INVX1_RVT U1163 ( .A(\add_x_3/A[1] ), .Y(n1638) );
  INVX1_RVT U1164 ( .A(\add_x_3/A[2] ), .Y(n1631) );
  INVX1_RVT U1165 ( .A(\add_x_3/A[3] ), .Y(n1628) );
  INVX1_RVT U1166 ( .A(\add_x_3/A[4] ), .Y(n1620) );
  INVX1_RVT U1167 ( .A(\add_x_3/A[5] ), .Y(n1614) );
  AND4X1_RVT U1168 ( .A1(n1631), .A2(n1628), .A3(n1620), .A4(n1614), .Y(n535)
         );
  AND4X1_RVT U1169 ( .A1(n1361), .A2(n1638), .A3(n1644), .A4(n535), .Y(n543)
         );
  NAND4X0_RVT U1170 ( .A1(n1405), .A2(n1392), .A3(n1383), .A4(n1370), .Y(n536)
         );
  NOR4X1_RVT U1171 ( .A1(\add_x_3/A[22] ), .A2(\add_x_3/A[23] ), .A3(
        m5stg_frac_dbl_nx), .A4(n536), .Y(n542) );
  INVX1_RVT U1172 ( .A(\add_x_3/A[10] ), .Y(n1570) );
  INVX1_RVT U1173 ( .A(\add_x_3/A[11] ), .Y(n1557) );
  NAND4X0_RVT U1174 ( .A1(n1570), .A2(n1557), .A3(n1548), .A4(n1536), .Y(n540)
         );
  INVX1_RVT U1175 ( .A(\add_x_3/A[6] ), .Y(n1605) );
  INVX1_RVT U1176 ( .A(\add_x_3/A[7] ), .Y(n1599) );
  INVX1_RVT U1177 ( .A(\add_x_3/A[8] ), .Y(n1589) );
  INVX1_RVT U1178 ( .A(\add_x_3/A[9] ), .Y(n1576) );
  NAND4X0_RVT U1179 ( .A1(n1605), .A2(n1599), .A3(n1589), .A4(n1576), .Y(n539)
         );
  NAND4X0_RVT U1180 ( .A1(n1484), .A2(n1467), .A3(n1456), .A4(n1440), .Y(n538)
         );
  NAND4X0_RVT U1181 ( .A1(n1526), .A2(n1515), .A3(n1504), .A4(n1492), .Y(n537)
         );
  NOR4X1_RVT U1182 ( .A1(n540), .A2(n539), .A3(n538), .A4(n537), .Y(n541) );
  NAND3X0_RVT U1183 ( .A1(n543), .A2(n542), .A3(n541), .Y(m5stg_frac_sng_nx)
         );
  AND4X1_RVT U1184 ( .A1(n1108), .A2(n1153), .A3(n1124), .A4(n1183), .Y(n550)
         );
  AND4X1_RVT U1185 ( .A1(n1212), .A2(n1261), .A3(n1246), .A4(n1276), .Y(n549)
         );
  AND4X1_RVT U1186 ( .A1(n1312), .A2(n1336), .A3(n1321), .A4(n1346), .Y(n544)
         );
  NAND4X0_RVT U1187 ( .A1(n553), .A2(n1290), .A3(n1298), .A4(n544), .Y(n547)
         );
  NAND4X0_RVT U1188 ( .A1(n913), .A2(n996), .A3(n982), .A4(n1013), .Y(n546) );
  NAND4X0_RVT U1189 ( .A1(n1028), .A2(n1064), .A3(n1044), .A4(n1086), .Y(n545)
         );
  NOR4X1_RVT U1190 ( .A1(m5stg_frac_sng_nx), .A2(n547), .A3(n546), .A4(n545), 
        .Y(n548) );
  NAND3X0_RVT U1191 ( .A1(n550), .A2(n549), .A3(n548), .Y(m5stg_frac_neq_0) );
  INVX1_RVT U1192 ( .A(mul_frac_out_fracadd), .Y(n762) );
  INVX1_RVT U1193 ( .A(mul_frac_out_frac), .Y(n761) );
  OA21X1_RVT U1194 ( .A1(n551), .A2(n762), .A3(n761), .Y(n556) );
  AO221X1_RVT U1195 ( .A1(n913), .A2(n553), .A3(n836), .A4(n555), .A5(n557), 
        .Y(n552) );
  OA22X1_RVT U1196 ( .A1(n553), .A2(n556), .A3(n762), .A4(n552), .Y(n554) );
  NAND2X0_RVT U1197 ( .A1(n554), .A2(n5), .Y(mul_frac_out_in[51]) );
  AO222X1_RVT U1198 ( .A1(n913), .A2(n762), .A3(n913), .A4(n557), .A5(n556), 
        .A6(n555), .Y(n558) );
  NAND2X0_RVT U1199 ( .A1(n558), .A2(n5), .Y(mul_frac_out_in[50]) );
  NAND2X0_RVT U1200 ( .A1(n566), .A2(n564), .Y(n559) );
  AO221X1_RVT U1201 ( .A1(n982), .A2(n559), .A3(n566), .A4(n561), .A5(n762), 
        .Y(n563) );
  AO21X1_RVT U1202 ( .A1(mul_frac_out_fracadd), .A2(n560), .A3(
        mul_frac_out_frac), .Y(n565) );
  NAND2X0_RVT U1203 ( .A1(n561), .A2(n565), .Y(n562) );
  NAND3X0_RVT U1204 ( .A1(n563), .A2(n562), .A3(n5), .Y(mul_frac_out_in[49])
         );
  NAND3X0_RVT U1205 ( .A1(mul_frac_out_fracadd), .A2(n996), .A3(n564), .Y(n568) );
  NAND2X0_RVT U1206 ( .A1(n566), .A2(n565), .Y(n567) );
  NAND3X0_RVT U1207 ( .A1(n568), .A2(n567), .A3(n5), .Y(mul_frac_out_in[48])
         );
  NAND2X0_RVT U1208 ( .A1(n576), .A2(n574), .Y(n569) );
  AO221X1_RVT U1209 ( .A1(n1013), .A2(n569), .A3(n576), .A4(n571), .A5(n762), 
        .Y(n573) );
  AO21X1_RVT U1210 ( .A1(mul_frac_out_fracadd), .A2(n570), .A3(
        mul_frac_out_frac), .Y(n575) );
  NAND2X0_RVT U1211 ( .A1(n571), .A2(n575), .Y(n572) );
  NAND3X0_RVT U1212 ( .A1(n573), .A2(n572), .A3(n5), .Y(mul_frac_out_in[47])
         );
  NAND3X0_RVT U1213 ( .A1(mul_frac_out_fracadd), .A2(n1028), .A3(n574), .Y(
        n578) );
  NAND2X0_RVT U1214 ( .A1(n576), .A2(n575), .Y(n577) );
  NAND3X0_RVT U1215 ( .A1(n578), .A2(n577), .A3(n5), .Y(mul_frac_out_in[46])
         );
  NAND2X0_RVT U1216 ( .A1(n586), .A2(n584), .Y(n579) );
  AO221X1_RVT U1217 ( .A1(n1044), .A2(n579), .A3(n586), .A4(n581), .A5(n762), 
        .Y(n583) );
  AO21X1_RVT U1218 ( .A1(mul_frac_out_fracadd), .A2(n580), .A3(
        mul_frac_out_frac), .Y(n585) );
  NAND2X0_RVT U1219 ( .A1(n581), .A2(n585), .Y(n582) );
  NAND3X0_RVT U1220 ( .A1(n583), .A2(n582), .A3(n5), .Y(mul_frac_out_in[45])
         );
  NAND3X0_RVT U1221 ( .A1(mul_frac_out_fracadd), .A2(n1064), .A3(n584), .Y(
        n588) );
  NAND2X0_RVT U1222 ( .A1(n586), .A2(n585), .Y(n587) );
  NAND3X0_RVT U1223 ( .A1(n588), .A2(n587), .A3(n5), .Y(mul_frac_out_in[44])
         );
  NAND2X0_RVT U1224 ( .A1(n596), .A2(n594), .Y(n589) );
  AO221X1_RVT U1225 ( .A1(n1086), .A2(n589), .A3(n596), .A4(n591), .A5(n762), 
        .Y(n593) );
  AO21X1_RVT U1226 ( .A1(mul_frac_out_fracadd), .A2(n590), .A3(
        mul_frac_out_frac), .Y(n595) );
  NAND2X0_RVT U1227 ( .A1(n591), .A2(n595), .Y(n592) );
  NAND3X0_RVT U1228 ( .A1(n593), .A2(n592), .A3(n5), .Y(mul_frac_out_in[43])
         );
  NAND3X0_RVT U1229 ( .A1(mul_frac_out_fracadd), .A2(n1108), .A3(n594), .Y(
        n598) );
  NAND2X0_RVT U1230 ( .A1(n596), .A2(n595), .Y(n597) );
  NAND3X0_RVT U1231 ( .A1(n598), .A2(n597), .A3(n5), .Y(mul_frac_out_in[42])
         );
  NAND2X0_RVT U1232 ( .A1(n606), .A2(n604), .Y(n599) );
  AO221X1_RVT U1233 ( .A1(n1124), .A2(n599), .A3(n606), .A4(n601), .A5(n762), 
        .Y(n603) );
  AO21X1_RVT U1234 ( .A1(mul_frac_out_fracadd), .A2(n600), .A3(
        mul_frac_out_frac), .Y(n605) );
  NAND2X0_RVT U1235 ( .A1(n601), .A2(n605), .Y(n602) );
  NAND3X0_RVT U1236 ( .A1(n603), .A2(n602), .A3(n5), .Y(mul_frac_out_in[41])
         );
  NAND3X0_RVT U1237 ( .A1(mul_frac_out_fracadd), .A2(n1153), .A3(n604), .Y(
        n608) );
  NAND2X0_RVT U1238 ( .A1(n606), .A2(n605), .Y(n607) );
  NAND3X0_RVT U1239 ( .A1(n608), .A2(n607), .A3(n5), .Y(mul_frac_out_in[40])
         );
  NAND2X0_RVT U1240 ( .A1(n616), .A2(n614), .Y(n609) );
  AO221X1_RVT U1241 ( .A1(n1183), .A2(n609), .A3(n616), .A4(n611), .A5(n762), 
        .Y(n613) );
  AO21X1_RVT U1242 ( .A1(mul_frac_out_fracadd), .A2(n610), .A3(
        mul_frac_out_frac), .Y(n615) );
  NAND2X0_RVT U1243 ( .A1(n611), .A2(n615), .Y(n612) );
  NAND3X0_RVT U1244 ( .A1(n613), .A2(n612), .A3(n5), .Y(mul_frac_out_in[39])
         );
  NAND3X0_RVT U1245 ( .A1(mul_frac_out_fracadd), .A2(n1212), .A3(n614), .Y(
        n618) );
  NAND2X0_RVT U1246 ( .A1(n616), .A2(n615), .Y(n617) );
  NAND3X0_RVT U1247 ( .A1(n618), .A2(n617), .A3(n5), .Y(mul_frac_out_in[38])
         );
  NAND2X0_RVT U1248 ( .A1(n626), .A2(n624), .Y(n619) );
  AO221X1_RVT U1249 ( .A1(n1246), .A2(n619), .A3(n626), .A4(n621), .A5(n762), 
        .Y(n623) );
  AO21X1_RVT U1250 ( .A1(mul_frac_out_fracadd), .A2(n620), .A3(
        mul_frac_out_frac), .Y(n625) );
  NAND2X0_RVT U1251 ( .A1(n621), .A2(n625), .Y(n622) );
  NAND3X0_RVT U1252 ( .A1(n623), .A2(n622), .A3(n5), .Y(mul_frac_out_in[37])
         );
  NAND3X0_RVT U1253 ( .A1(mul_frac_out_fracadd), .A2(n1261), .A3(n624), .Y(
        n628) );
  NAND2X0_RVT U1254 ( .A1(n626), .A2(n625), .Y(n627) );
  NAND3X0_RVT U1255 ( .A1(n628), .A2(n627), .A3(n5), .Y(mul_frac_out_in[36])
         );
  NAND2X0_RVT U1256 ( .A1(n636), .A2(n634), .Y(n629) );
  AO221X1_RVT U1257 ( .A1(n1276), .A2(n629), .A3(n636), .A4(n631), .A5(n762), 
        .Y(n633) );
  AO21X1_RVT U1258 ( .A1(mul_frac_out_fracadd), .A2(n630), .A3(
        mul_frac_out_frac), .Y(n635) );
  NAND2X0_RVT U1259 ( .A1(n631), .A2(n635), .Y(n632) );
  NAND3X0_RVT U1260 ( .A1(n633), .A2(n632), .A3(n5), .Y(mul_frac_out_in[35])
         );
  NAND3X0_RVT U1261 ( .A1(mul_frac_out_fracadd), .A2(n1290), .A3(n634), .Y(
        n638) );
  NAND2X0_RVT U1262 ( .A1(n636), .A2(n635), .Y(n637) );
  NAND3X0_RVT U1263 ( .A1(n638), .A2(n637), .A3(n5), .Y(mul_frac_out_in[34])
         );
  NAND2X0_RVT U1264 ( .A1(n646), .A2(n644), .Y(n639) );
  AO221X1_RVT U1265 ( .A1(n1298), .A2(n639), .A3(n646), .A4(n641), .A5(n762), 
        .Y(n643) );
  AO21X1_RVT U1266 ( .A1(mul_frac_out_fracadd), .A2(n640), .A3(
        mul_frac_out_frac), .Y(n645) );
  NAND2X0_RVT U1267 ( .A1(n641), .A2(n645), .Y(n642) );
  NAND3X0_RVT U1268 ( .A1(n643), .A2(n642), .A3(n5), .Y(mul_frac_out_in[33])
         );
  NAND3X0_RVT U1269 ( .A1(mul_frac_out_fracadd), .A2(n1312), .A3(n644), .Y(
        n648) );
  NAND2X0_RVT U1270 ( .A1(n646), .A2(n645), .Y(n647) );
  NAND3X0_RVT U1271 ( .A1(n648), .A2(n647), .A3(n5), .Y(mul_frac_out_in[32])
         );
  NAND2X0_RVT U1272 ( .A1(n655), .A2(n653), .Y(n649) );
  AO221X1_RVT U1273 ( .A1(n1321), .A2(n649), .A3(n655), .A4(n650), .A5(n762), 
        .Y(n652) );
  OAI21X1_RVT U1274 ( .A1(n762), .A2(n653), .A3(n761), .Y(n654) );
  NAND2X0_RVT U1275 ( .A1(n650), .A2(n654), .Y(n651) );
  NAND3X0_RVT U1276 ( .A1(n652), .A2(n651), .A3(n5), .Y(mul_frac_out_in[31])
         );
  NAND3X0_RVT U1277 ( .A1(mul_frac_out_fracadd), .A2(n1336), .A3(n653), .Y(
        n657) );
  NAND2X0_RVT U1278 ( .A1(n655), .A2(n654), .Y(n656) );
  NAND3X0_RVT U1279 ( .A1(n657), .A2(n656), .A3(n5), .Y(mul_frac_out_in[30])
         );
  HADDX1_RVT U1280 ( .A0(n661), .B0(m5stg_fmuls), .SO(n658) );
  HADDX1_RVT U1281 ( .A0(n1346), .B0(n658), .SO(n659) );
  OA22X1_RVT U1282 ( .A1(n761), .A2(n1346), .A3(n762), .A4(n659), .Y(n660) );
  NAND2X0_RVT U1283 ( .A1(n660), .A2(n5), .Y(mul_frac_out_in[29]) );
  NAND3X0_RVT U1284 ( .A1(n671), .A2(\add_x_3/A[26] ), .A3(\add_x_3/A[27] ), 
        .Y(n662) );
  NAND2X0_RVT U1285 ( .A1(n1361), .A2(n662), .Y(n663) );
  NAND3X0_RVT U1286 ( .A1(mul_frac_out_fracadd), .A2(n664), .A3(n663), .Y(n666) );
  NAND2X0_RVT U1287 ( .A1(mul_frac_out_frac), .A2(\add_x_3/A[28] ), .Y(n665)
         );
  NAND3X0_RVT U1288 ( .A1(n5), .A2(n666), .A3(n665), .Y(mul_frac_out_in[28])
         );
  NAND2X0_RVT U1289 ( .A1(\add_x_3/A[26] ), .A2(n671), .Y(n667) );
  AO221X1_RVT U1290 ( .A1(n1370), .A2(n667), .A3(\add_x_3/A[26] ), .A4(
        \add_x_3/A[27] ), .A5(n762), .Y(n670) );
  NAND3X0_RVT U1291 ( .A1(n679), .A2(\add_x_3/A[24] ), .A3(\add_x_3/A[25] ), 
        .Y(n668) );
  AO21X1_RVT U1292 ( .A1(mul_frac_out_fracadd), .A2(n668), .A3(
        mul_frac_out_frac), .Y(n672) );
  NAND2X0_RVT U1293 ( .A1(\add_x_3/A[27] ), .A2(n672), .Y(n669) );
  NAND3X0_RVT U1294 ( .A1(n670), .A2(n669), .A3(n5), .Y(mul_frac_out_in[27])
         );
  NAND3X0_RVT U1295 ( .A1(mul_frac_out_fracadd), .A2(n671), .A3(n1383), .Y(
        n674) );
  NAND2X0_RVT U1296 ( .A1(\add_x_3/A[26] ), .A2(n672), .Y(n673) );
  NAND3X0_RVT U1297 ( .A1(n674), .A2(n673), .A3(n5), .Y(mul_frac_out_in[26])
         );
  NAND2X0_RVT U1298 ( .A1(\add_x_3/A[24] ), .A2(n679), .Y(n675) );
  AO221X1_RVT U1299 ( .A1(n1392), .A2(n675), .A3(\add_x_3/A[24] ), .A4(
        \add_x_3/A[25] ), .A5(n762), .Y(n678) );
  AO21X1_RVT U1300 ( .A1(mul_frac_out_fracadd), .A2(n676), .A3(
        mul_frac_out_frac), .Y(n680) );
  NAND2X0_RVT U1301 ( .A1(\add_x_3/A[25] ), .A2(n680), .Y(n677) );
  NAND3X0_RVT U1302 ( .A1(n678), .A2(n677), .A3(n5), .Y(mul_frac_out_in[25])
         );
  NAND3X0_RVT U1303 ( .A1(mul_frac_out_fracadd), .A2(n679), .A3(n1405), .Y(
        n682) );
  NAND2X0_RVT U1304 ( .A1(\add_x_3/A[24] ), .A2(n680), .Y(n681) );
  NAND3X0_RVT U1305 ( .A1(n682), .A2(n681), .A3(n5), .Y(mul_frac_out_in[24])
         );
  NAND2X0_RVT U1306 ( .A1(\add_x_3/A[22] ), .A2(n687), .Y(n683) );
  AO221X1_RVT U1307 ( .A1(n1420), .A2(n683), .A3(\add_x_3/A[22] ), .A4(
        \add_x_3/A[23] ), .A5(n762), .Y(n686) );
  AO21X1_RVT U1308 ( .A1(mul_frac_out_fracadd), .A2(n684), .A3(
        mul_frac_out_frac), .Y(n688) );
  NAND2X0_RVT U1309 ( .A1(\add_x_3/A[23] ), .A2(n688), .Y(n685) );
  NAND3X0_RVT U1310 ( .A1(n686), .A2(n685), .A3(n5), .Y(mul_frac_out_in[23])
         );
  NAND3X0_RVT U1311 ( .A1(mul_frac_out_fracadd), .A2(n687), .A3(n1431), .Y(
        n690) );
  NAND2X0_RVT U1312 ( .A1(\add_x_3/A[22] ), .A2(n688), .Y(n689) );
  NAND3X0_RVT U1313 ( .A1(n690), .A2(n689), .A3(n5), .Y(mul_frac_out_in[22])
         );
  NAND2X0_RVT U1314 ( .A1(\add_x_3/A[20] ), .A2(n695), .Y(n691) );
  AO221X1_RVT U1315 ( .A1(n1440), .A2(n691), .A3(\add_x_3/A[20] ), .A4(
        \add_x_3/A[21] ), .A5(n762), .Y(n694) );
  AO21X1_RVT U1316 ( .A1(mul_frac_out_fracadd), .A2(n692), .A3(
        mul_frac_out_frac), .Y(n696) );
  NAND2X0_RVT U1317 ( .A1(\add_x_3/A[21] ), .A2(n696), .Y(n693) );
  NAND3X0_RVT U1318 ( .A1(n694), .A2(n693), .A3(n5), .Y(mul_frac_out_in[21])
         );
  NAND3X0_RVT U1319 ( .A1(mul_frac_out_fracadd), .A2(n695), .A3(n1456), .Y(
        n698) );
  NAND2X0_RVT U1320 ( .A1(\add_x_3/A[20] ), .A2(n696), .Y(n697) );
  NAND3X0_RVT U1321 ( .A1(n698), .A2(n697), .A3(n5), .Y(mul_frac_out_in[20])
         );
  NAND2X0_RVT U1322 ( .A1(\add_x_3/A[18] ), .A2(n703), .Y(n699) );
  AO221X1_RVT U1323 ( .A1(n1467), .A2(n699), .A3(\add_x_3/A[18] ), .A4(
        \add_x_3/A[19] ), .A5(n762), .Y(n702) );
  AO21X1_RVT U1324 ( .A1(mul_frac_out_fracadd), .A2(n700), .A3(
        mul_frac_out_frac), .Y(n704) );
  NAND2X0_RVT U1325 ( .A1(\add_x_3/A[19] ), .A2(n704), .Y(n701) );
  NAND3X0_RVT U1326 ( .A1(n702), .A2(n701), .A3(n5), .Y(mul_frac_out_in[19])
         );
  NAND3X0_RVT U1327 ( .A1(mul_frac_out_fracadd), .A2(n703), .A3(n1484), .Y(
        n706) );
  NAND2X0_RVT U1328 ( .A1(\add_x_3/A[18] ), .A2(n704), .Y(n705) );
  NAND3X0_RVT U1329 ( .A1(n706), .A2(n705), .A3(n5), .Y(mul_frac_out_in[18])
         );
  NAND2X0_RVT U1330 ( .A1(m5stg_frac_32_0[19]), .A2(n711), .Y(n707) );
  AO221X1_RVT U1331 ( .A1(n1492), .A2(n707), .A3(m5stg_frac_32_0[19]), .A4(
        m5stg_frac_32_0[20]), .A5(n762), .Y(n710) );
  AO21X1_RVT U1332 ( .A1(mul_frac_out_fracadd), .A2(n708), .A3(
        mul_frac_out_frac), .Y(n712) );
  NAND2X0_RVT U1333 ( .A1(m5stg_frac_32_0[20]), .A2(n712), .Y(n709) );
  NAND3X0_RVT U1334 ( .A1(n710), .A2(n709), .A3(n5), .Y(mul_frac_out_in[17])
         );
  NAND3X0_RVT U1335 ( .A1(mul_frac_out_fracadd), .A2(n711), .A3(n1504), .Y(
        n714) );
  NAND2X0_RVT U1336 ( .A1(m5stg_frac_32_0[19]), .A2(n712), .Y(n713) );
  NAND3X0_RVT U1337 ( .A1(n714), .A2(n713), .A3(n5), .Y(mul_frac_out_in[16])
         );
  NAND2X0_RVT U1338 ( .A1(\add_x_3/A[14] ), .A2(n499), .Y(n715) );
  AO221X1_RVT U1339 ( .A1(n1515), .A2(n715), .A3(\add_x_3/A[14] ), .A4(
        \add_x_3/A[15] ), .A5(n762), .Y(n718) );
  AO21X1_RVT U1340 ( .A1(mul_frac_out_fracadd), .A2(n716), .A3(
        mul_frac_out_frac), .Y(n719) );
  NAND2X0_RVT U1341 ( .A1(\add_x_3/A[15] ), .A2(n719), .Y(n717) );
  NAND3X0_RVT U1342 ( .A1(n718), .A2(n717), .A3(n5), .Y(mul_frac_out_in[15])
         );
  NAND3X0_RVT U1343 ( .A1(mul_frac_out_fracadd), .A2(n499), .A3(n1526), .Y(
        n721) );
  NAND2X0_RVT U1344 ( .A1(\add_x_3/A[14] ), .A2(n719), .Y(n720) );
  NAND3X0_RVT U1345 ( .A1(n721), .A2(n720), .A3(n5), .Y(mul_frac_out_in[14])
         );
  NAND2X0_RVT U1346 ( .A1(\add_x_3/A[12] ), .A2(n726), .Y(n722) );
  AO221X1_RVT U1347 ( .A1(n1536), .A2(n722), .A3(\add_x_3/A[12] ), .A4(
        \add_x_3/A[13] ), .A5(n762), .Y(n725) );
  AO21X1_RVT U1348 ( .A1(mul_frac_out_fracadd), .A2(n723), .A3(
        mul_frac_out_frac), .Y(n727) );
  NAND2X0_RVT U1349 ( .A1(\add_x_3/A[13] ), .A2(n727), .Y(n724) );
  NAND3X0_RVT U1350 ( .A1(n725), .A2(n724), .A3(n5), .Y(mul_frac_out_in[13])
         );
  NAND3X0_RVT U1351 ( .A1(mul_frac_out_fracadd), .A2(n726), .A3(n1548), .Y(
        n729) );
  NAND2X0_RVT U1352 ( .A1(\add_x_3/A[12] ), .A2(n727), .Y(n728) );
  NAND3X0_RVT U1353 ( .A1(n729), .A2(n728), .A3(n5), .Y(mul_frac_out_in[12])
         );
  OA21X1_RVT U1354 ( .A1(n730), .A2(n762), .A3(n761), .Y(n733) );
  AO221X1_RVT U1355 ( .A1(n1570), .A2(n1557), .A3(\add_x_3/A[11] ), .A4(
        \add_x_3/A[10] ), .A5(n734), .Y(n731) );
  OA22X1_RVT U1356 ( .A1(n1557), .A2(n733), .A3(n762), .A4(n731), .Y(n732) );
  NAND2X0_RVT U1357 ( .A1(n732), .A2(n5), .Y(mul_frac_out_in[11]) );
  AO222X1_RVT U1358 ( .A1(n1570), .A2(n762), .A3(n1570), .A4(n734), .A5(n733), 
        .A6(\add_x_3/A[10] ), .Y(n735) );
  NAND2X0_RVT U1359 ( .A1(n735), .A2(n5), .Y(mul_frac_out_in[10]) );
  OA21X1_RVT U1360 ( .A1(n736), .A2(n762), .A3(n761), .Y(n739) );
  AO221X1_RVT U1361 ( .A1(n1589), .A2(n1576), .A3(\add_x_3/A[9] ), .A4(
        \add_x_3/A[8] ), .A5(n740), .Y(n737) );
  OA22X1_RVT U1362 ( .A1(n1576), .A2(n739), .A3(n762), .A4(n737), .Y(n738) );
  NAND2X0_RVT U1363 ( .A1(n738), .A2(n5), .Y(mul_frac_out_in[9]) );
  AO222X1_RVT U1364 ( .A1(n1589), .A2(n762), .A3(n1589), .A4(n740), .A5(n739), 
        .A6(\add_x_3/A[8] ), .Y(n741) );
  NAND2X0_RVT U1365 ( .A1(n5), .A2(n741), .Y(mul_frac_out_in[8]) );
  OA21X1_RVT U1366 ( .A1(n742), .A2(n762), .A3(n761), .Y(n745) );
  AO221X1_RVT U1367 ( .A1(n1605), .A2(n1599), .A3(\add_x_3/A[7] ), .A4(
        \add_x_3/A[6] ), .A5(n746), .Y(n743) );
  OA22X1_RVT U1368 ( .A1(n1599), .A2(n745), .A3(n762), .A4(n743), .Y(n744) );
  NAND2X0_RVT U1369 ( .A1(n744), .A2(n5), .Y(mul_frac_out_in[7]) );
  AO222X1_RVT U1370 ( .A1(n1605), .A2(n762), .A3(n1605), .A4(n746), .A5(n745), 
        .A6(\add_x_3/A[6] ), .Y(n747) );
  NAND2X0_RVT U1371 ( .A1(n747), .A2(n5), .Y(mul_frac_out_in[6]) );
  OA21X1_RVT U1372 ( .A1(n748), .A2(n762), .A3(n761), .Y(n751) );
  AO221X1_RVT U1373 ( .A1(n1620), .A2(n1614), .A3(\add_x_3/A[5] ), .A4(
        \add_x_3/A[4] ), .A5(n752), .Y(n749) );
  OA22X1_RVT U1374 ( .A1(n1614), .A2(n751), .A3(n762), .A4(n749), .Y(n750) );
  NAND2X0_RVT U1375 ( .A1(n750), .A2(n5), .Y(mul_frac_out_in[5]) );
  AO222X1_RVT U1376 ( .A1(n1620), .A2(n762), .A3(n1620), .A4(n752), .A5(n751), 
        .A6(\add_x_3/A[4] ), .Y(n753) );
  NAND2X0_RVT U1377 ( .A1(n753), .A2(n5), .Y(mul_frac_out_in[4]) );
  OA21X1_RVT U1378 ( .A1(n754), .A2(n762), .A3(n761), .Y(n757) );
  AO221X1_RVT U1379 ( .A1(n1631), .A2(n1628), .A3(\add_x_3/A[3] ), .A4(
        \add_x_3/A[2] ), .A5(n758), .Y(n755) );
  OA22X1_RVT U1380 ( .A1(n1628), .A2(n757), .A3(n762), .A4(n755), .Y(n756) );
  NAND2X0_RVT U1381 ( .A1(n756), .A2(n5), .Y(mul_frac_out_in[3]) );
  AO222X1_RVT U1382 ( .A1(n1631), .A2(n762), .A3(n1631), .A4(n758), .A5(n757), 
        .A6(\add_x_3/A[2] ), .Y(n759) );
  NAND2X0_RVT U1383 ( .A1(n759), .A2(n5), .Y(mul_frac_out_in[2]) );
  NAND2X0_RVT U1384 ( .A1(m5stg_fmulda), .A2(\add_x_3/A[0] ), .Y(n760) );
  AO221X1_RVT U1385 ( .A1(n1638), .A2(n760), .A3(\add_x_3/A[1] ), .A4(
        \add_x_3/A[0] ), .A5(n762), .Y(n764) );
  OAI21X1_RVT U1386 ( .A1(n762), .A2(m5stg_fmulda), .A3(n761), .Y(n765) );
  NAND2X0_RVT U1387 ( .A1(\add_x_3/A[1] ), .A2(n765), .Y(n763) );
  NAND3X0_RVT U1388 ( .A1(n764), .A2(n763), .A3(n5), .Y(mul_frac_out_in[1]) );
  NAND3X0_RVT U1389 ( .A1(mul_frac_out_fracadd), .A2(n1644), .A3(m5stg_fmulda), 
        .Y(n767) );
  NAND2X0_RVT U1390 ( .A1(\add_x_3/A[0] ), .A2(n765), .Y(n766) );
  NAND3X0_RVT U1391 ( .A1(n767), .A2(n766), .A3(n5), .Y(mul_frac_out_in[0]) );
  AND4X1_RVT U1392 ( .A1(n771), .A2(n770), .A3(n769), .A4(n768), .Y(n1154) );
  NAND2X0_RVT U1393 ( .A1(n2069), .A2(n1879), .Y(n1632) );
  INVX1_RVT U1394 ( .A(n1632), .Y(n1891) );
  NAND2X0_RVT U1395 ( .A1(n6), .A2(n1891), .Y(n1219) );
  NAND2X0_RVT U1396 ( .A1(n1268), .A2(n1891), .Y(n1221) );
  OA22X1_RVT U1397 ( .A1(m4stg_frac[96]), .A2(n772), .A3(m4stg_frac[95]), .A4(
        n842), .Y(n774) );
  OA22X1_RVT U1398 ( .A1(m4stg_frac[94]), .A2(n844), .A3(m4stg_frac[93]), .A4(
        n779), .Y(n773) );
  NAND2X0_RVT U1399 ( .A1(n774), .A2(n773), .Y(n1065) );
  OA22X1_RVT U1400 ( .A1(n1154), .A2(n1219), .A3(n1221), .A4(n1065), .Y(n835)
         );
  NAND2X0_RVT U1401 ( .A1(n1894), .A2(n2069), .Y(n1213) );
  INVX1_RVT U1402 ( .A(n1213), .Y(n1090) );
  NAND2X0_RVT U1403 ( .A1(n1593), .A2(m4stg_frac[104]), .Y(n776) );
  AO22X1_RVT U1404 ( .A1(m4stg_sh_cnt[0]), .A2(m4stg_frac[101]), .A3(n778), 
        .A4(m4stg_frac[102]), .Y(n974) );
  NAND2X0_RVT U1405 ( .A1(m4stg_sh_cnt[1]), .A2(n974), .Y(n775) );
  NAND3X0_RVT U1406 ( .A1(n777), .A2(n776), .A3(n775), .Y(n780) );
  NAND3X0_RVT U1407 ( .A1(m4stg_sh_cnt[2]), .A2(n2101), .A3(n2069), .Y(n1215)
         );
  INVX1_RVT U1408 ( .A(n1215), .Y(n1088) );
  AO22X1_RVT U1409 ( .A1(m4stg_sh_cnt[0]), .A2(m4stg_frac[99]), .A3(n778), 
        .A4(m4stg_frac[100]), .Y(n976) );
  OA222X1_RVT U1410 ( .A1(n779), .A2(m4stg_frac[97]), .A3(n844), .A4(
        m4stg_frac[98]), .A5(n976), .A6(m4stg_sh_cnt[1]), .Y(n1004) );
  AOI22X1_RVT U1411 ( .A1(n1090), .A2(n780), .A3(n1088), .A4(n1004), .Y(n834)
         );
  NAND4X0_RVT U1412 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .Y(n1165) );
  NAND2X0_RVT U1413 ( .A1(n1539), .A2(n1165), .Y(n794) );
  AND4X1_RVT U1414 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .Y(n1166) );
  NAND4X0_RVT U1415 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .Y(n1175) );
  OA22X1_RVT U1416 ( .A1(n1166), .A2(n1616), .A3(n1075), .A4(n1095), .Y(n793)
         );
  AND2X1_RVT U1417 ( .A1(n794), .A2(n793), .Y(n800) );
  NAND4X0_RVT U1418 ( .A1(n798), .A2(n797), .A3(n796), .A4(n795), .Y(n1068) );
  NAND2X0_RVT U1419 ( .A1(n1068), .A2(n1582), .Y(n799) );
  AND2X1_RVT U1420 ( .A1(n800), .A2(n799), .Y(n1457) );
  AO22X1_RVT U1421 ( .A1(n1579), .A2(m4stg_frac[47]), .A3(n1593), .A4(
        m4stg_frac[48]), .Y(n802) );
  AO22X1_RVT U1422 ( .A1(n1573), .A2(m4stg_frac[46]), .A3(n1422), .A4(
        m4stg_frac[45]), .Y(n801) );
  OR2X1_RVT U1423 ( .A1(n802), .A2(n801), .Y(n1173) );
  AO22X1_RVT U1424 ( .A1(n1579), .A2(m4stg_frac[43]), .A3(n1593), .A4(
        m4stg_frac[44]), .Y(n804) );
  AO22X1_RVT U1425 ( .A1(n1573), .A2(m4stg_frac[42]), .A3(n1422), .A4(
        m4stg_frac[41]), .Y(n803) );
  OR2X1_RVT U1426 ( .A1(n804), .A2(n803), .Y(n1158) );
  AO22X1_RVT U1427 ( .A1(n1268), .A2(n1173), .A3(n6), .A4(n1158), .Y(n813) );
  AOI22X1_RVT U1428 ( .A1(n1573), .A2(m4stg_frac[50]), .A3(n1422), .A4(
        m4stg_frac[49]), .Y(n807) );
  NAND2X0_RVT U1429 ( .A1(n1579), .A2(m4stg_frac[51]), .Y(n805) );
  NAND3X0_RVT U1430 ( .A1(n807), .A2(n806), .A3(n805), .Y(n1174) );
  NAND2X0_RVT U1431 ( .A1(n1422), .A2(m4stg_frac[53]), .Y(n808) );
  NAND4X0_RVT U1432 ( .A1(n811), .A2(n810), .A3(n809), .A4(n808), .Y(n1176) );
  AO22X1_RVT U1433 ( .A1(n1582), .A2(n1174), .A3(n1539), .A4(n1176), .Y(n812)
         );
  NOR2X0_RVT U1434 ( .A1(n813), .A2(n812), .Y(n1621) );
  OA22X1_RVT U1435 ( .A1(n1457), .A2(n257), .A3(n1621), .A4(n1625), .Y(n833)
         );
  AND2X1_RVT U1436 ( .A1(m4stg_sh_cnt[4]), .A2(n2069), .Y(n1651) );
  AND4X1_RVT U1437 ( .A1(n817), .A2(n816), .A3(n815), .A4(n814), .Y(n1157) );
  NAND4X0_RVT U1438 ( .A1(n821), .A2(n820), .A3(n819), .A4(n818), .Y(n997) );
  INVX1_RVT U1439 ( .A(n997), .Y(n1170) );
  OA22X1_RVT U1440 ( .A1(n1157), .A2(n1616), .A3(n1170), .A4(n1095), .Y(n831)
         );
  NAND4X0_RVT U1441 ( .A1(n825), .A2(n824), .A3(n823), .A4(n822), .Y(n1067) );
  INVX1_RVT U1442 ( .A(n1067), .Y(n1156) );
  NAND4X0_RVT U1443 ( .A1(n829), .A2(n828), .A3(n827), .A4(n826), .Y(n1066) );
  INVX1_RVT U1444 ( .A(n1066), .Y(n1155) );
  OA22X1_RVT U1445 ( .A1(n1156), .A2(n35), .A3(n1155), .A4(n1623), .Y(n830) );
  NAND2X0_RVT U1446 ( .A1(n831), .A2(n830), .Y(n1262) );
  NAND2X0_RVT U1447 ( .A1(n1651), .A2(n1262), .Y(n832) );
  NAND4X0_RVT U1448 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .Y(
        m4stg_shl_54) );
  AND2X1_RVT U1449 ( .A1(m4stg_left_shift_step), .A2(m4stg_shl_55), .Y(n1973)
         );
  AOI22X1_RVT U1450 ( .A1(n1973), .A2(m4stg_shl_54), .A3(n836), .A4(n1972), 
        .Y(n1878) );
  NAND4X0_RVT U1451 ( .A1(n840), .A2(n839), .A3(n838), .A4(n837), .Y(n848) );
  OA22X1_RVT U1452 ( .A1(n844), .A2(n843), .A3(n842), .A4(n841), .Y(n847) );
  NAND3X0_RVT U1453 ( .A1(n847), .A2(n846), .A3(n845), .Y(n1014) );
  OAI221X1_RVT U1454 ( .A1(m4stg_sh_cnt[2]), .A2(n848), .A3(n1908), .A4(n1014), 
        .A5(n2101), .Y(n879) );
  NAND4X0_RVT U1455 ( .A1(n852), .A2(n851), .A3(n850), .A4(n849), .Y(n1089) );
  NAND4X0_RVT U1456 ( .A1(n856), .A2(n855), .A3(n854), .A4(n853), .Y(n1087) );
  AOI22X1_RVT U1457 ( .A1(n858), .A2(n1089), .A3(n857), .A4(n1087), .Y(n878)
         );
  AND4X1_RVT U1458 ( .A1(n862), .A2(n861), .A3(n860), .A4(n859), .Y(n1186) );
  AND4X1_RVT U1459 ( .A1(n866), .A2(n865), .A3(n864), .A4(n863), .Y(n1205) );
  OA22X1_RVT U1460 ( .A1(n1186), .A2(n1616), .A3(n1205), .A4(n1095), .Y(n876)
         );
  AND4X1_RVT U1461 ( .A1(n870), .A2(n869), .A3(n868), .A4(n867), .Y(n1187) );
  AND4X1_RVT U1462 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .Y(n1185) );
  OA22X1_RVT U1463 ( .A1(n1187), .A2(n35), .A3(n1185), .A4(n1623), .Y(n875) );
  NAND2X0_RVT U1464 ( .A1(n876), .A2(n875), .Y(n1277) );
  NAND2X0_RVT U1465 ( .A1(m4stg_sh_cnt[4]), .A2(n1277), .Y(n877) );
  NAND3X0_RVT U1466 ( .A1(n879), .A2(n878), .A3(n877), .Y(n912) );
  AO22X1_RVT U1467 ( .A1(n1579), .A2(m4stg_frac[42]), .A3(n1593), .A4(
        m4stg_frac[43]), .Y(n881) );
  AO22X1_RVT U1468 ( .A1(n1573), .A2(m4stg_frac[41]), .A3(n1422), .A4(
        m4stg_frac[40]), .Y(n880) );
  OR2X1_RVT U1469 ( .A1(n881), .A2(n880), .Y(n1188) );
  INVX1_RVT U1470 ( .A(n1188), .Y(n1017) );
  AO22X1_RVT U1471 ( .A1(n1579), .A2(m4stg_frac[46]), .A3(n1593), .A4(
        m4stg_frac[47]), .Y(n883) );
  AO22X1_RVT U1472 ( .A1(n1573), .A2(m4stg_frac[45]), .A3(n1422), .A4(
        m4stg_frac[44]), .Y(n882) );
  OR2X1_RVT U1473 ( .A1(n883), .A2(n882), .Y(n1091) );
  INVX1_RVT U1474 ( .A(n1091), .Y(n1197) );
  OA22X1_RVT U1475 ( .A1(n1017), .A2(n1095), .A3(n1197), .A4(n1616), .Y(n893)
         );
  AOI22X1_RVT U1476 ( .A1(n1422), .A2(m4stg_frac[48]), .A3(n1579), .A4(
        m4stg_frac[50]), .Y(n884) );
  AND2X1_RVT U1477 ( .A1(n885), .A2(n884), .Y(n887) );
  NAND2X0_RVT U1478 ( .A1(m4stg_frac[49]), .A2(n1573), .Y(n886) );
  AND2X1_RVT U1479 ( .A1(n887), .A2(n886), .Y(n1196) );
  AND4X1_RVT U1480 ( .A1(n891), .A2(n890), .A3(n889), .A4(n888), .Y(n1199) );
  OA22X1_RVT U1481 ( .A1(n1196), .A2(n35), .A3(n1199), .A4(n1623), .Y(n892) );
  NAND2X0_RVT U1482 ( .A1(n893), .A2(n892), .Y(n1469) );
  AND4X1_RVT U1483 ( .A1(n897), .A2(n896), .A3(n895), .A4(n894), .Y(n1202) );
  AND4X1_RVT U1484 ( .A1(n901), .A2(n900), .A3(n899), .A4(n898), .Y(n1198) );
  OA22X1_RVT U1485 ( .A1(n1202), .A2(n1616), .A3(n1198), .A4(n1095), .Y(n911)
         );
  AND4X1_RVT U1486 ( .A1(n905), .A2(n904), .A3(n903), .A4(n902), .Y(n1203) );
  AND4X1_RVT U1487 ( .A1(n909), .A2(n908), .A3(n907), .A4(n906), .Y(n1204) );
  OA22X1_RVT U1488 ( .A1(n1203), .A2(n35), .A3(n1204), .A4(n1623), .Y(n910) );
  NAND2X0_RVT U1489 ( .A1(n911), .A2(n910), .Y(n1468) );
  AOI222X1_RVT U1490 ( .A1(n912), .A2(n2069), .A3(n1469), .A4(n1647), .A5(
        n1468), .A6(n1916), .Y(n2035) );
  INVX1_RVT U1491 ( .A(n1973), .Y(n1652) );
  OA22X1_RVT U1492 ( .A1(n913), .A2(m6stg_step), .A3(n2035), .A4(n1652), .Y(
        n1877) );
  NAND4X0_RVT U1493 ( .A1(n917), .A2(n916), .A3(n915), .A4(n914), .Y(n1110) );
  NAND4X0_RVT U1494 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .Y(n1109) );
  OA22X1_RVT U1495 ( .A1(n1221), .A2(n1110), .A3(n1219), .A4(n1109), .Y(n981)
         );
  NAND4X0_RVT U1496 ( .A1(n925), .A2(n924), .A3(n923), .A4(n922), .Y(n1236) );
  NAND4X0_RVT U1497 ( .A1(n929), .A2(n928), .A3(n927), .A4(n926), .Y(n1232) );
  OA22X1_RVT U1498 ( .A1(n1616), .A2(n1236), .A3(n1095), .A4(n1232), .Y(n939)
         );
  NAND4X0_RVT U1499 ( .A1(n933), .A2(n932), .A3(n931), .A4(n930), .Y(n1237) );
  NAND4X0_RVT U1500 ( .A1(n937), .A2(n936), .A3(n935), .A4(n934), .Y(n1239) );
  OA22X1_RVT U1501 ( .A1(n35), .A2(n1237), .A3(n1623), .A4(n1239), .Y(n938) );
  AND2X1_RVT U1502 ( .A1(n939), .A2(n938), .Y(n1485) );
  AO22X1_RVT U1503 ( .A1(n1579), .A2(m4stg_frac[45]), .A3(n1593), .A4(
        m4stg_frac[46]), .Y(n941) );
  AO22X1_RVT U1504 ( .A1(n1573), .A2(m4stg_frac[44]), .A3(n1422), .A4(
        m4stg_frac[43]), .Y(n940) );
  OR2X1_RVT U1505 ( .A1(n941), .A2(n940), .Y(n1230) );
  AO22X1_RVT U1506 ( .A1(n1579), .A2(m4stg_frac[41]), .A3(n1593), .A4(
        m4stg_frac[42]), .Y(n943) );
  AO22X1_RVT U1507 ( .A1(n1573), .A2(m4stg_frac[40]), .A3(n1422), .A4(
        m4stg_frac[39]), .Y(n942) );
  OR2X1_RVT U1508 ( .A1(n943), .A2(n942), .Y(n1223) );
  OA22X1_RVT U1509 ( .A1(n1616), .A2(n1230), .A3(n1095), .A4(n1223), .Y(n950)
         );
  AO22X1_RVT U1510 ( .A1(n1579), .A2(m4stg_frac[49]), .A3(n1593), .A4(
        m4stg_frac[50]), .Y(n945) );
  AO22X1_RVT U1511 ( .A1(n1573), .A2(m4stg_frac[48]), .A3(n1422), .A4(
        m4stg_frac[47]), .Y(n944) );
  OR2X1_RVT U1512 ( .A1(n945), .A2(n944), .Y(n1231) );
  NAND3X0_RVT U1513 ( .A1(n948), .A2(n947), .A3(n946), .Y(n1233) );
  OA22X1_RVT U1514 ( .A1(n35), .A2(n1231), .A3(n1623), .A4(n1233), .Y(n949) );
  AND2X1_RVT U1515 ( .A1(n950), .A2(n949), .Y(n1633) );
  OA22X1_RVT U1516 ( .A1(n1485), .A2(n257), .A3(n1633), .A4(n1625), .Y(n980)
         );
  NAND4X0_RVT U1517 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .Y(n1218) );
  NAND4X0_RVT U1518 ( .A1(n958), .A2(n957), .A3(n956), .A4(n955), .Y(n1238) );
  OA22X1_RVT U1519 ( .A1(n1616), .A2(n1218), .A3(n1095), .A4(n1238), .Y(n968)
         );
  NAND4X0_RVT U1520 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .Y(n1217) );
  NAND4X0_RVT U1521 ( .A1(n966), .A2(n965), .A3(n964), .A4(n963), .Y(n1111) );
  OA22X1_RVT U1522 ( .A1(n35), .A2(n1217), .A3(n1623), .A4(n1111), .Y(n967) );
  NAND2X0_RVT U1523 ( .A1(n968), .A2(n967), .Y(n1296) );
  NAND2X0_RVT U1524 ( .A1(n1651), .A2(n1296), .Y(n979) );
  NAND2X0_RVT U1525 ( .A1(n1593), .A2(m4stg_frac[98]), .Y(n971) );
  NAND4X0_RVT U1526 ( .A1(n972), .A2(n971), .A3(n970), .A4(n969), .Y(n1029) );
  NAND2X0_RVT U1527 ( .A1(n2101), .A2(n2069), .Y(n973) );
  AO221X1_RVT U1528 ( .A1(m4stg_sh_cnt[1]), .A2(n976), .A3(n975), .A4(n974), 
        .A5(n973), .Y(n977) );
  AO22X1_RVT U1529 ( .A1(m4stg_sh_cnt[2]), .A2(n1029), .A3(n1215), .A4(n977), 
        .Y(n978) );
  NAND4X0_RVT U1530 ( .A1(n981), .A2(n980), .A3(n979), .A4(n978), .Y(n2034) );
  OA22X1_RVT U1531 ( .A1(n982), .A2(m6stg_step), .A3(n2034), .A4(n1652), .Y(
        n1876) );
  AOI22X1_RVT U1532 ( .A1(n1088), .A2(n1045), .A3(n1090), .A4(n983), .Y(n995)
         );
  OA22X1_RVT U1533 ( .A1(n1126), .A2(n1221), .A3(n1125), .A4(n1219), .Y(n994)
         );
  OA22X1_RVT U1534 ( .A1(n1140), .A2(n1095), .A3(n1139), .A4(n1616), .Y(n985)
         );
  OA22X1_RVT U1535 ( .A1(n1144), .A2(n1623), .A3(n1143), .A4(n35), .Y(n984) );
  AND2X1_RVT U1536 ( .A1(n985), .A2(n984), .Y(n1493) );
  AO22X1_RVT U1537 ( .A1(n1579), .A2(m4stg_frac[40]), .A3(n1593), .A4(
        m4stg_frac[41]), .Y(n987) );
  AO22X1_RVT U1538 ( .A1(n1573), .A2(m4stg_frac[39]), .A3(n1422), .A4(
        m4stg_frac[38]), .Y(n986) );
  OR2X1_RVT U1539 ( .A1(n987), .A2(n986), .Y(n1250) );
  INVX1_RVT U1540 ( .A(n1250), .Y(n1050) );
  OA22X1_RVT U1541 ( .A1(n1050), .A2(n1095), .A3(n1053), .A4(n1616), .Y(n989)
         );
  OA22X1_RVT U1542 ( .A1(n1138), .A2(n35), .A3(n1137), .A4(n1623), .Y(n988) );
  AND2X1_RVT U1543 ( .A1(n989), .A2(n988), .Y(n1639) );
  OA22X1_RVT U1544 ( .A1(n1493), .A2(n257), .A3(n1639), .A4(n1625), .Y(n993)
         );
  OA22X1_RVT U1545 ( .A1(n1146), .A2(n1616), .A3(n1145), .A4(n1095), .Y(n991)
         );
  OA22X1_RVT U1546 ( .A1(n1127), .A2(n1623), .A3(n1128), .A4(n35), .Y(n990) );
  NAND2X0_RVT U1547 ( .A1(n991), .A2(n990), .Y(n1299) );
  NAND2X0_RVT U1548 ( .A1(n1651), .A2(n1299), .Y(n992) );
  AND4X1_RVT U1549 ( .A1(n995), .A2(n994), .A3(n993), .A4(n992), .Y(n2033) );
  OA22X1_RVT U1550 ( .A1(n996), .A2(m6stg_step), .A3(n2033), .A4(n1652), .Y(
        n1875) );
  OA22X1_RVT U1551 ( .A1(n1616), .A2(n997), .A3(n1095), .A4(n1165), .Y(n999)
         );
  AOI22X1_RVT U1552 ( .A1(n1582), .A2(n1157), .A3(n1539), .A4(n1156), .Y(n998)
         );
  NAND2X0_RVT U1553 ( .A1(n999), .A2(n998), .Y(n1313) );
  AO22X1_RVT U1554 ( .A1(n1579), .A2(m4stg_frac[39]), .A3(n1593), .A4(
        m4stg_frac[40]), .Y(n1001) );
  AO22X1_RVT U1555 ( .A1(n1573), .A2(m4stg_frac[38]), .A3(n1422), .A4(
        m4stg_frac[37]), .Y(n1000) );
  OR2X1_RVT U1556 ( .A1(n1001), .A2(n1000), .Y(n1265) );
  OA22X1_RVT U1557 ( .A1(n1616), .A2(n1158), .A3(n1095), .A4(n1265), .Y(n1003)
         );
  OA22X1_RVT U1558 ( .A1(n35), .A2(n1173), .A3(n1623), .A4(n1174), .Y(n1002)
         );
  NAND2X0_RVT U1559 ( .A1(n1003), .A2(n1002), .Y(n1645) );
  AOI22X1_RVT U1560 ( .A1(n1651), .A2(n1313), .A3(n1647), .A4(n1645), .Y(n1012) );
  AO22X1_RVT U1561 ( .A1(m4stg_sh_cnt[2]), .A2(n1065), .A3(n1908), .A4(n1005), 
        .Y(n1007) );
  AO22X1_RVT U1562 ( .A1(m4stg_sh_cnt[2]), .A2(n1155), .A3(n1908), .A4(n1154), 
        .Y(n1006) );
  OAI221X1_RVT U1563 ( .A1(m4stg_sh_cnt[3]), .A2(n1007), .A3(n1636), .A4(n1006), .A5(n1891), .Y(n1011) );
  OA22X1_RVT U1564 ( .A1(n1616), .A2(n1175), .A3(n1095), .A4(n1176), .Y(n1009)
         );
  AOI22X1_RVT U1565 ( .A1(n1582), .A2(n1166), .A3(n1539), .A4(n1167), .Y(n1008) );
  NAND2X0_RVT U1566 ( .A1(n1009), .A2(n1008), .Y(n1505) );
  NAND2X0_RVT U1567 ( .A1(n1916), .A2(n1505), .Y(n1010) );
  NAND3X0_RVT U1568 ( .A1(n1012), .A2(n1011), .A3(n1010), .Y(n2031) );
  OA22X1_RVT U1569 ( .A1(n1013), .A2(m6stg_step), .A3(n2031), .A4(n1652), .Y(
        n1874) );
  AOI22X1_RVT U1570 ( .A1(n1090), .A2(n1014), .A3(n1088), .A4(n1089), .Y(n1027) );
  INVX1_RVT U1571 ( .A(n1087), .Y(n1184) );
  OA22X1_RVT U1572 ( .A1(n1185), .A2(n1219), .A3(n1184), .A4(n1221), .Y(n1026)
         );
  AO22X1_RVT U1573 ( .A1(n1579), .A2(m4stg_frac[38]), .A3(n1593), .A4(
        m4stg_frac[39]), .Y(n1016) );
  AO22X1_RVT U1574 ( .A1(n1573), .A2(m4stg_frac[37]), .A3(n1422), .A4(
        m4stg_frac[36]), .Y(n1015) );
  OR2X1_RVT U1575 ( .A1(n1016), .A2(n1015), .Y(n1280) );
  INVX1_RVT U1576 ( .A(n1280), .Y(n1094) );
  OA22X1_RVT U1577 ( .A1(n1094), .A2(n1095), .A3(n1017), .A4(n1616), .Y(n1019)
         );
  OA22X1_RVT U1578 ( .A1(n1197), .A2(n35), .A3(n1196), .A4(n1623), .Y(n1018)
         );
  AND2X1_RVT U1579 ( .A1(n1019), .A2(n1018), .Y(n1650) );
  OA22X1_RVT U1580 ( .A1(n1199), .A2(n1095), .A3(n1198), .A4(n1616), .Y(n1021)
         );
  OA22X1_RVT U1581 ( .A1(n1203), .A2(n1623), .A3(n1202), .A4(n35), .Y(n1020)
         );
  AND2X1_RVT U1582 ( .A1(n1021), .A2(n1020), .Y(n1516) );
  OA22X1_RVT U1583 ( .A1(n1650), .A2(n1625), .A3(n1516), .A4(n257), .Y(n1025)
         );
  OA22X1_RVT U1584 ( .A1(n1205), .A2(n1616), .A3(n1204), .A4(n1095), .Y(n1023)
         );
  OA22X1_RVT U1585 ( .A1(n1187), .A2(n1623), .A3(n1186), .A4(n35), .Y(n1022)
         );
  NAND2X0_RVT U1586 ( .A1(n1023), .A2(n1022), .Y(n1322) );
  NAND2X0_RVT U1587 ( .A1(n1651), .A2(n1322), .Y(n1024) );
  AND4X1_RVT U1588 ( .A1(n1027), .A2(n1026), .A3(n1025), .A4(n1024), .Y(n2030)
         );
  OA22X1_RVT U1589 ( .A1(n1028), .A2(m6stg_step), .A3(n2030), .A4(n1652), .Y(
        n1873) );
  AOI22X1_RVT U1590 ( .A1(n1090), .A2(n1029), .A3(n1088), .A4(n1110), .Y(n1043) );
  OA22X1_RVT U1591 ( .A1(n1216), .A2(n1219), .A3(n1214), .A4(n1221), .Y(n1042)
         );
  NAND2X0_RVT U1592 ( .A1(n1539), .A2(n1231), .Y(n1033) );
  AO22X1_RVT U1593 ( .A1(n1579), .A2(m4stg_frac[37]), .A3(n1593), .A4(
        m4stg_frac[38]), .Y(n1031) );
  AO22X1_RVT U1594 ( .A1(n1573), .A2(m4stg_frac[36]), .A3(n1422), .A4(
        m4stg_frac[35]), .Y(n1030) );
  OR2X1_RVT U1595 ( .A1(n1031), .A2(n1030), .Y(n1293) );
  AOI22X1_RVT U1596 ( .A1(n1223), .A2(n1268), .A3(n1293), .A4(n6), .Y(n1032)
         );
  AND2X1_RVT U1597 ( .A1(n1033), .A2(n1032), .Y(n1035) );
  NAND2X0_RVT U1598 ( .A1(n1230), .A2(n1582), .Y(n1034) );
  AND2X1_RVT U1599 ( .A1(n1035), .A2(n1034), .Y(n1528) );
  AO22X1_RVT U1600 ( .A1(n1268), .A2(n1232), .A3(n6), .A4(n1233), .Y(n1037) );
  AO22X1_RVT U1601 ( .A1(n1582), .A2(n1236), .A3(n1539), .A4(n1237), .Y(n1036)
         );
  NOR2X0_RVT U1602 ( .A1(n1037), .A2(n1036), .Y(n1527) );
  OA22X1_RVT U1603 ( .A1(n1528), .A2(n1625), .A3(n1527), .A4(n257), .Y(n1041)
         );
  AO22X1_RVT U1604 ( .A1(n1268), .A2(n1238), .A3(n6), .A4(n1239), .Y(n1039) );
  AO22X1_RVT U1605 ( .A1(n1582), .A2(n1218), .A3(n1539), .A4(n1217), .Y(n1038)
         );
  OR2X1_RVT U1606 ( .A1(n1039), .A2(n1038), .Y(n1344) );
  NAND2X0_RVT U1607 ( .A1(n1651), .A2(n1344), .Y(n1040) );
  AND4X1_RVT U1608 ( .A1(n1043), .A2(n1042), .A3(n1041), .A4(n1040), .Y(n2029)
         );
  OA22X1_RVT U1609 ( .A1(n1044), .A2(m6stg_step), .A3(n2029), .A4(n1652), .Y(
        n1872) );
  AOI22X1_RVT U1610 ( .A1(n1088), .A2(n1046), .A3(n1090), .A4(n1045), .Y(n1063) );
  OA22X1_RVT U1611 ( .A1(n1125), .A2(n1221), .A3(n1127), .A4(n1219), .Y(n1062)
         );
  NAND2X0_RVT U1612 ( .A1(n1539), .A2(n1047), .Y(n1052) );
  AO22X1_RVT U1613 ( .A1(n1579), .A2(m4stg_frac[36]), .A3(n1593), .A4(
        m4stg_frac[37]), .Y(n1049) );
  AO22X1_RVT U1614 ( .A1(n1573), .A2(m4stg_frac[35]), .A3(n1422), .A4(
        m4stg_frac[34]), .Y(n1048) );
  OR2X1_RVT U1615 ( .A1(n1049), .A2(n1048), .Y(n1302) );
  OA22X1_RVT U1616 ( .A1(n1132), .A2(n1095), .A3(n1050), .A4(n1616), .Y(n1051)
         );
  AND2X1_RVT U1617 ( .A1(n1052), .A2(n1051), .Y(n1055) );
  NAND2X0_RVT U1618 ( .A1(n1129), .A2(n1582), .Y(n1054) );
  AND2X1_RVT U1619 ( .A1(n1055), .A2(n1054), .Y(n1888) );
  OA22X1_RVT U1620 ( .A1(n1137), .A2(n1095), .A3(n1140), .A4(n1616), .Y(n1057)
         );
  OA22X1_RVT U1621 ( .A1(n1143), .A2(n1623), .A3(n1139), .A4(n35), .Y(n1056)
         );
  AND2X1_RVT U1622 ( .A1(n1057), .A2(n1056), .Y(n1537) );
  OA22X1_RVT U1623 ( .A1(n1888), .A2(n1625), .A3(n1537), .A4(n257), .Y(n1061)
         );
  OA22X1_RVT U1624 ( .A1(n1144), .A2(n1095), .A3(n1145), .A4(n1616), .Y(n1059)
         );
  OA22X1_RVT U1625 ( .A1(n1128), .A2(n1623), .A3(n1146), .A4(n35), .Y(n1058)
         );
  NAND2X0_RVT U1626 ( .A1(n1059), .A2(n1058), .Y(n1347) );
  NAND2X0_RVT U1627 ( .A1(n1651), .A2(n1347), .Y(n1060) );
  AND4X1_RVT U1628 ( .A1(n1063), .A2(n1062), .A3(n1061), .A4(n1060), .Y(n2028)
         );
  OA22X1_RVT U1629 ( .A1(n1064), .A2(m6stg_step), .A3(n2028), .A4(n1652), .Y(
        n1871) );
  AOI22X1_RVT U1630 ( .A1(n1090), .A2(n1065), .A3(n1154), .A4(n1088), .Y(n1085) );
  OA22X1_RVT U1631 ( .A1(n1067), .A2(n1219), .A3(n1066), .A4(n1221), .Y(n1084)
         );
  NAND2X0_RVT U1632 ( .A1(n1539), .A2(n1157), .Y(n1070) );
  OA22X1_RVT U1633 ( .A1(n1616), .A2(n1165), .A3(n1095), .A4(n1068), .Y(n1069)
         );
  AND2X1_RVT U1634 ( .A1(n1070), .A2(n1069), .Y(n1072) );
  NAND2X0_RVT U1635 ( .A1(n1170), .A2(n1582), .Y(n1071) );
  AND2X1_RVT U1636 ( .A1(n1072), .A2(n1071), .Y(n1363) );
  NAND2X0_RVT U1637 ( .A1(n1539), .A2(n1166), .Y(n1074) );
  OA22X1_RVT U1638 ( .A1(n1616), .A2(n1176), .A3(n1095), .A4(n1174), .Y(n1073)
         );
  AND2X1_RVT U1639 ( .A1(n1074), .A2(n1073), .Y(n1077) );
  NAND2X0_RVT U1640 ( .A1(n1075), .A2(n1582), .Y(n1076) );
  AND2X1_RVT U1641 ( .A1(n1077), .A2(n1076), .Y(n1362) );
  OA22X1_RVT U1642 ( .A1(n1363), .A2(n397), .A3(n1362), .A4(n257), .Y(n1083)
         );
  AO22X1_RVT U1643 ( .A1(n1579), .A2(m4stg_frac[35]), .A3(n1593), .A4(
        m4stg_frac[36]), .Y(n1079) );
  AO22X1_RVT U1644 ( .A1(n1573), .A2(m4stg_frac[34]), .A3(n1422), .A4(
        m4stg_frac[33]), .Y(n1078) );
  OR2X1_RVT U1645 ( .A1(n1079), .A2(n1078), .Y(n1316) );
  OA22X1_RVT U1646 ( .A1(n1316), .A2(n1095), .A3(n1616), .A4(n1265), .Y(n1081)
         );
  OA22X1_RVT U1647 ( .A1(n35), .A2(n1158), .A3(n1623), .A4(n1173), .Y(n1080)
         );
  NAND2X0_RVT U1648 ( .A1(n1081), .A2(n1080), .Y(n1549) );
  NAND2X0_RVT U1649 ( .A1(n1647), .A2(n1549), .Y(n1082) );
  NAND4X0_RVT U1650 ( .A1(n1085), .A2(n1084), .A3(n1083), .A4(n1082), .Y(n2027) );
  OA22X1_RVT U1651 ( .A1(n1086), .A2(m6stg_step), .A3(n2027), .A4(n1652), .Y(
        n1870) );
  AOI22X1_RVT U1652 ( .A1(n1090), .A2(n1089), .A3(n1088), .A4(n1087), .Y(n1107) );
  OA22X1_RVT U1653 ( .A1(n1187), .A2(n1219), .A3(n1185), .A4(n1221), .Y(n1106)
         );
  NAND2X0_RVT U1654 ( .A1(n1539), .A2(n1091), .Y(n1097) );
  AO22X1_RVT U1655 ( .A1(n1579), .A2(m4stg_frac[34]), .A3(n1593), .A4(
        m4stg_frac[35]), .Y(n1093) );
  AO22X1_RVT U1656 ( .A1(n1573), .A2(m4stg_frac[33]), .A3(n1422), .A4(
        m4stg_frac[32]), .Y(n1092) );
  OR2X1_RVT U1657 ( .A1(n1093), .A2(n1092), .Y(n1325) );
  OA22X1_RVT U1658 ( .A1(n1191), .A2(n1095), .A3(n1094), .A4(n1616), .Y(n1096)
         );
  AND2X1_RVT U1659 ( .A1(n1097), .A2(n1096), .Y(n1099) );
  NAND2X0_RVT U1660 ( .A1(n1188), .A2(n1582), .Y(n1098) );
  AND2X1_RVT U1661 ( .A1(n1099), .A2(n1098), .Y(n1904) );
  OA22X1_RVT U1662 ( .A1(n1196), .A2(n1095), .A3(n1199), .A4(n1616), .Y(n1101)
         );
  OA22X1_RVT U1663 ( .A1(n1202), .A2(n1623), .A3(n1198), .A4(n35), .Y(n1100)
         );
  AND2X1_RVT U1664 ( .A1(n1101), .A2(n1100), .Y(n1558) );
  OA22X1_RVT U1665 ( .A1(n1904), .A2(n1625), .A3(n1558), .A4(n257), .Y(n1105)
         );
  OA22X1_RVT U1666 ( .A1(n1203), .A2(n1095), .A3(n1204), .A4(n1616), .Y(n1103)
         );
  OA22X1_RVT U1667 ( .A1(n1186), .A2(n1623), .A3(n1205), .A4(n35), .Y(n1102)
         );
  NAND2X0_RVT U1668 ( .A1(n1103), .A2(n1102), .Y(n1371) );
  NAND2X0_RVT U1669 ( .A1(n1651), .A2(n1371), .Y(n1104) );
  AND4X1_RVT U1670 ( .A1(n1107), .A2(n1106), .A3(n1105), .A4(n1104), .Y(n2026)
         );
  OA22X1_RVT U1671 ( .A1(n1108), .A2(m6stg_step), .A3(n2026), .A4(n1652), .Y(
        n1869) );
  OA22X1_RVT U1672 ( .A1(n1213), .A2(n1110), .A3(n1215), .A4(n1109), .Y(n1123)
         );
  OA22X1_RVT U1673 ( .A1(n1221), .A2(n1111), .A3(n1219), .A4(n1217), .Y(n1122)
         );
  OA22X1_RVT U1674 ( .A1(n1616), .A2(n1239), .A3(n1095), .A4(n1237), .Y(n1113)
         );
  OA22X1_RVT U1675 ( .A1(n35), .A2(n1238), .A3(n1623), .A4(n1218), .Y(n1112)
         );
  AND2X1_RVT U1676 ( .A1(n1113), .A2(n1112), .Y(n1384) );
  OA22X1_RVT U1677 ( .A1(n1616), .A2(n1233), .A3(n1095), .A4(n1231), .Y(n1115)
         );
  OA22X1_RVT U1678 ( .A1(n35), .A2(n1232), .A3(n1623), .A4(n1236), .Y(n1114)
         );
  AND2X1_RVT U1679 ( .A1(n1115), .A2(n1114), .Y(n1571) );
  OA22X1_RVT U1680 ( .A1(n1384), .A2(n397), .A3(n1571), .A4(n257), .Y(n1121)
         );
  AO22X1_RVT U1681 ( .A1(n1579), .A2(m4stg_frac[33]), .A3(n1593), .A4(
        m4stg_frac[34]), .Y(n1117) );
  AO22X1_RVT U1682 ( .A1(n1573), .A2(m4stg_frac[32]), .A3(n1422), .A4(
        m4stg_frac[31]), .Y(n1116) );
  OR2X1_RVT U1683 ( .A1(n1117), .A2(n1116), .Y(n1337) );
  OA22X1_RVT U1684 ( .A1(n1616), .A2(n1293), .A3(n1095), .A4(n1337), .Y(n1119)
         );
  OA22X1_RVT U1685 ( .A1(n35), .A2(n1223), .A3(n1623), .A4(n1230), .Y(n1118)
         );
  NAND2X0_RVT U1686 ( .A1(n1119), .A2(n1118), .Y(n1901) );
  NAND2X0_RVT U1687 ( .A1(n1647), .A2(n1901), .Y(n1120) );
  NAND4X0_RVT U1688 ( .A1(n1123), .A2(n1122), .A3(n1121), .A4(n1120), .Y(n2025) );
  OA22X1_RVT U1689 ( .A1(n1124), .A2(m6stg_step), .A3(n2025), .A4(n1652), .Y(
        n1868) );
  OA22X1_RVT U1690 ( .A1(n1126), .A2(n1213), .A3(n1125), .A4(n1215), .Y(n1152)
         );
  OA22X1_RVT U1691 ( .A1(n1128), .A2(n1219), .A3(n1127), .A4(n1221), .Y(n1151)
         );
  NAND2X0_RVT U1692 ( .A1(n1539), .A2(n1129), .Y(n1134) );
  AO22X1_RVT U1693 ( .A1(n1579), .A2(m4stg_frac[32]), .A3(n1593), .A4(
        m4stg_frac[33]), .Y(n1131) );
  AO22X1_RVT U1694 ( .A1(n1573), .A2(m4stg_frac[31]), .A3(m4stg_frac[30]), 
        .A4(n1422), .Y(n1130) );
  OR2X1_RVT U1695 ( .A1(n1131), .A2(n1130), .Y(n1350) );
  INVX1_RVT U1696 ( .A(n1350), .Y(n1253) );
  OA22X1_RVT U1697 ( .A1(n1253), .A2(n1095), .A3(n1132), .A4(n1616), .Y(n1133)
         );
  AND2X1_RVT U1698 ( .A1(n1134), .A2(n1133), .Y(n1136) );
  NAND2X0_RVT U1699 ( .A1(n1250), .A2(n1582), .Y(n1135) );
  AND2X1_RVT U1700 ( .A1(n1136), .A2(n1135), .Y(n1903) );
  OA22X1_RVT U1701 ( .A1(n1138), .A2(n1095), .A3(n1137), .A4(n1616), .Y(n1142)
         );
  OA22X1_RVT U1702 ( .A1(n1140), .A2(n35), .A3(n1139), .A4(n1623), .Y(n1141)
         );
  AND2X1_RVT U1703 ( .A1(n1142), .A2(n1141), .Y(n1577) );
  OA22X1_RVT U1704 ( .A1(n1903), .A2(n1625), .A3(n1577), .A4(n257), .Y(n1150)
         );
  OA22X1_RVT U1705 ( .A1(n1144), .A2(n1616), .A3(n1143), .A4(n1095), .Y(n1148)
         );
  OA22X1_RVT U1706 ( .A1(n1146), .A2(n1623), .A3(n1145), .A4(n35), .Y(n1147)
         );
  NAND2X0_RVT U1707 ( .A1(n1148), .A2(n1147), .Y(n1393) );
  NAND2X0_RVT U1708 ( .A1(n1651), .A2(n1393), .Y(n1149) );
  AND4X1_RVT U1709 ( .A1(n1152), .A2(n1151), .A3(n1150), .A4(n1149), .Y(n2024)
         );
  OA22X1_RVT U1710 ( .A1(n1153), .A2(m6stg_step), .A3(n2024), .A4(n1652), .Y(
        n1867) );
  OA22X1_RVT U1711 ( .A1(n1155), .A2(n1215), .A3(n1154), .A4(n1213), .Y(n1182)
         );
  OA22X1_RVT U1712 ( .A1(n1157), .A2(n1219), .A3(n1156), .A4(n1221), .Y(n1181)
         );
  NAND2X0_RVT U1713 ( .A1(n1539), .A2(n1158), .Y(n1162) );
  AO22X1_RVT U1714 ( .A1(n1579), .A2(m4stg_frac[31]), .A3(n1593), .A4(
        m4stg_frac[32]), .Y(n1160) );
  AO22X1_RVT U1715 ( .A1(n1573), .A2(m4stg_frac[30]), .A3(n1422), .A4(
        m4stg_frac[29]), .Y(n1159) );
  OR2X1_RVT U1716 ( .A1(n1160), .A2(n1159), .Y(n1366) );
  AOI22X1_RVT U1717 ( .A1(n1316), .A2(n1268), .A3(n1366), .A4(n6), .Y(n1161)
         );
  AND2X1_RVT U1718 ( .A1(n1162), .A2(n1161), .Y(n1164) );
  NAND2X0_RVT U1719 ( .A1(n1265), .A2(n1582), .Y(n1163) );
  AND2X1_RVT U1720 ( .A1(n1164), .A2(n1163), .Y(n1902) );
  NAND2X0_RVT U1721 ( .A1(n1582), .A2(n1165), .Y(n1169) );
  OA22X1_RVT U1722 ( .A1(n1167), .A2(n1616), .A3(n1166), .A4(n1095), .Y(n1168)
         );
  AND2X1_RVT U1723 ( .A1(n1169), .A2(n1168), .Y(n1172) );
  NAND2X0_RVT U1724 ( .A1(n997), .A2(n1539), .Y(n1171) );
  AND2X1_RVT U1725 ( .A1(n1172), .A2(n1171), .Y(n1406) );
  OA22X1_RVT U1726 ( .A1(n1902), .A2(n1625), .A3(n1406), .A4(n397), .Y(n1180)
         );
  AO22X1_RVT U1727 ( .A1(n1268), .A2(n1174), .A3(n6), .A4(n1173), .Y(n1178) );
  AO22X1_RVT U1728 ( .A1(n1582), .A2(n1176), .A3(n1539), .A4(n1175), .Y(n1177)
         );
  OR2X1_RVT U1729 ( .A1(n1178), .A2(n1177), .Y(n1590) );
  NAND2X0_RVT U1730 ( .A1(n1916), .A2(n1590), .Y(n1179) );
  AND4X1_RVT U1731 ( .A1(n1182), .A2(n1181), .A3(n1180), .A4(n1179), .Y(n2023)
         );
  OA22X1_RVT U1732 ( .A1(n1183), .A2(m6stg_step), .A3(n2023), .A4(n1652), .Y(
        n1866) );
  OA22X1_RVT U1733 ( .A1(n1185), .A2(n1215), .A3(n1184), .A4(n1213), .Y(n1211)
         );
  OA22X1_RVT U1734 ( .A1(n1187), .A2(n1221), .A3(n1186), .A4(n1219), .Y(n1210)
         );
  NAND2X0_RVT U1735 ( .A1(n1539), .A2(n1188), .Y(n1193) );
  AO22X1_RVT U1736 ( .A1(m4stg_frac[30]), .A2(n1579), .A3(m4stg_frac[31]), 
        .A4(n1593), .Y(n1190) );
  AO22X1_RVT U1737 ( .A1(n1573), .A2(m4stg_frac[29]), .A3(n1422), .A4(
        m4stg_frac[28]), .Y(n1189) );
  NOR2X0_RVT U1738 ( .A1(n1190), .A2(n1189), .Y(n1378) );
  OA22X1_RVT U1739 ( .A1(n1378), .A2(n1095), .A3(n1191), .A4(n1616), .Y(n1192)
         );
  AND2X1_RVT U1740 ( .A1(n1193), .A2(n1192), .Y(n1195) );
  NAND2X0_RVT U1741 ( .A1(n1280), .A2(n1582), .Y(n1194) );
  AND2X1_RVT U1742 ( .A1(n1195), .A2(n1194), .Y(n1601) );
  OA22X1_RVT U1743 ( .A1(n1197), .A2(n1095), .A3(n1196), .A4(n1616), .Y(n1201)
         );
  OA22X1_RVT U1744 ( .A1(n1199), .A2(n35), .A3(n1198), .A4(n1623), .Y(n1200)
         );
  AND2X1_RVT U1745 ( .A1(n1201), .A2(n1200), .Y(n1600) );
  OA22X1_RVT U1746 ( .A1(n1601), .A2(n1625), .A3(n1600), .A4(n257), .Y(n1209)
         );
  OA22X1_RVT U1747 ( .A1(n1203), .A2(n1616), .A3(n1202), .A4(n1095), .Y(n1207)
         );
  OA22X1_RVT U1748 ( .A1(n1205), .A2(n1623), .A3(n1204), .A4(n35), .Y(n1206)
         );
  NAND2X0_RVT U1749 ( .A1(n1207), .A2(n1206), .Y(n1429) );
  NAND2X0_RVT U1750 ( .A1(n1651), .A2(n1429), .Y(n1208) );
  AND4X1_RVT U1751 ( .A1(n1211), .A2(n1210), .A3(n1209), .A4(n1208), .Y(n2022)
         );
  OA22X1_RVT U1752 ( .A1(n1212), .A2(m6stg_step), .A3(n2022), .A4(n1652), .Y(
        n1865) );
  OA22X1_RVT U1753 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), .Y(n1245)
         );
  OA22X1_RVT U1754 ( .A1(n1222), .A2(n1221), .A3(n1220), .A4(n1219), .Y(n1244)
         );
  NAND2X0_RVT U1755 ( .A1(n1539), .A2(n1223), .Y(n1227) );
  AO22X1_RVT U1756 ( .A1(m4stg_frac[30]), .A2(n1593), .A3(m4stg_frac[29]), 
        .A4(n1579), .Y(n1225) );
  AO22X1_RVT U1757 ( .A1(n1573), .A2(m4stg_frac[28]), .A3(n1422), .A4(
        m4stg_frac[27]), .Y(n1224) );
  OR2X1_RVT U1758 ( .A1(n1225), .A2(n1224), .Y(n1387) );
  AOI22X1_RVT U1759 ( .A1(n1387), .A2(n6), .A3(n1337), .A4(n1268), .Y(n1226)
         );
  AND2X1_RVT U1760 ( .A1(n1227), .A2(n1226), .Y(n1229) );
  NAND2X0_RVT U1761 ( .A1(n1293), .A2(n1582), .Y(n1228) );
  AND2X1_RVT U1762 ( .A1(n1229), .A2(n1228), .Y(n1607) );
  AO22X1_RVT U1763 ( .A1(n1268), .A2(n1231), .A3(n6), .A4(n1230), .Y(n1235) );
  AO22X1_RVT U1764 ( .A1(n1582), .A2(n1233), .A3(n1539), .A4(n1232), .Y(n1234)
         );
  NOR2X0_RVT U1765 ( .A1(n1235), .A2(n1234), .Y(n1606) );
  OA22X1_RVT U1766 ( .A1(n1607), .A2(n1625), .A3(n1606), .A4(n257), .Y(n1243)
         );
  AO22X1_RVT U1767 ( .A1(n1268), .A2(n1237), .A3(n6), .A4(n1236), .Y(n1241) );
  AO22X1_RVT U1768 ( .A1(n1582), .A2(n1239), .A3(n1539), .A4(n1238), .Y(n1240)
         );
  OR2X1_RVT U1769 ( .A1(n1241), .A2(n1240), .Y(n1438) );
  NAND2X0_RVT U1770 ( .A1(n1651), .A2(n1438), .Y(n1242) );
  AND4X1_RVT U1771 ( .A1(n1245), .A2(n1244), .A3(n1243), .A4(n1242), .Y(n2021)
         );
  OA22X1_RVT U1772 ( .A1(n1246), .A2(m6stg_step), .A3(n2021), .A4(n1652), .Y(
        n1864) );
  NAND2X0_RVT U1773 ( .A1(n1916), .A2(n1442), .Y(n1249) );
  AOI22X1_RVT U1774 ( .A1(n1651), .A2(n1441), .A3(n1891), .A4(n1247), .Y(n1248) );
  AND2X1_RVT U1775 ( .A1(n1249), .A2(n1248), .Y(n1260) );
  NAND2X0_RVT U1776 ( .A1(n1539), .A2(n1250), .Y(n1255) );
  AO22X1_RVT U1777 ( .A1(m4stg_frac[29]), .A2(n1593), .A3(n1579), .A4(
        m4stg_frac[28]), .Y(n1252) );
  AO22X1_RVT U1778 ( .A1(n1573), .A2(m4stg_frac[27]), .A3(n1422), .A4(
        m4stg_frac[26]), .Y(n1251) );
  NOR2X0_RVT U1779 ( .A1(n1252), .A2(n1251), .Y(n1400) );
  OA22X1_RVT U1780 ( .A1(n1400), .A2(n1095), .A3(n1253), .A4(n1616), .Y(n1254)
         );
  AND2X1_RVT U1781 ( .A1(n1255), .A2(n1254), .Y(n1257) );
  NAND2X0_RVT U1782 ( .A1(n1302), .A2(n1582), .Y(n1256) );
  AND2X1_RVT U1783 ( .A1(n1257), .A2(n1256), .Y(n1957) );
  INVX1_RVT U1784 ( .A(n1957), .Y(n1258) );
  NAND2X0_RVT U1785 ( .A1(n1258), .A2(n1647), .Y(n1259) );
  AND2X1_RVT U1786 ( .A1(n1260), .A2(n1259), .Y(n2020) );
  OA22X1_RVT U1787 ( .A1(n1261), .A2(m6stg_step), .A3(n2020), .A4(n1652), .Y(
        n1863) );
  NAND2X0_RVT U1788 ( .A1(n1891), .A2(n1262), .Y(n1264) );
  OA22X1_RVT U1789 ( .A1(n1457), .A2(n397), .A3(n1621), .A4(n257), .Y(n1263)
         );
  AND2X1_RVT U1790 ( .A1(n1264), .A2(n1263), .Y(n1275) );
  NAND2X0_RVT U1791 ( .A1(n1539), .A2(n1265), .Y(n1270) );
  AO22X1_RVT U1792 ( .A1(n1579), .A2(m4stg_frac[27]), .A3(n1593), .A4(
        m4stg_frac[28]), .Y(n1267) );
  AO22X1_RVT U1793 ( .A1(n1573), .A2(m4stg_frac[26]), .A3(n1422), .A4(
        m4stg_frac[25]), .Y(n1266) );
  OR2X1_RVT U1794 ( .A1(n1267), .A2(n1266), .Y(n1409) );
  AOI22X1_RVT U1795 ( .A1(n1409), .A2(n6), .A3(n1366), .A4(n1268), .Y(n1269)
         );
  AND2X1_RVT U1796 ( .A1(n1270), .A2(n1269), .Y(n1272) );
  NAND2X0_RVT U1797 ( .A1(n1316), .A2(n1582), .Y(n1271) );
  AND2X1_RVT U1798 ( .A1(n1272), .A2(n1271), .Y(n1956) );
  INVX1_RVT U1799 ( .A(n1956), .Y(n1273) );
  NAND2X0_RVT U1800 ( .A1(n1273), .A2(n1647), .Y(n1274) );
  AND2X1_RVT U1801 ( .A1(n1275), .A2(n1274), .Y(n2019) );
  OA22X1_RVT U1802 ( .A1(n1276), .A2(m6stg_step), .A3(n2019), .A4(n1652), .Y(
        n1862) );
  NAND2X0_RVT U1803 ( .A1(n1916), .A2(n1469), .Y(n1279) );
  AOI22X1_RVT U1804 ( .A1(n1651), .A2(n1468), .A3(n1891), .A4(n1277), .Y(n1278) );
  AND2X1_RVT U1805 ( .A1(n1279), .A2(n1278), .Y(n1289) );
  NAND2X0_RVT U1806 ( .A1(n1539), .A2(n1280), .Y(n1284) );
  AO22X1_RVT U1807 ( .A1(n1579), .A2(m4stg_frac[26]), .A3(n1593), .A4(
        m4stg_frac[27]), .Y(n1282) );
  AO22X1_RVT U1808 ( .A1(n1573), .A2(m4stg_frac[25]), .A3(n1422), .A4(
        m4stg_frac[24]), .Y(n1281) );
  OR2X1_RVT U1809 ( .A1(n1282), .A2(n1281), .Y(n1421) );
  INVX1_RVT U1810 ( .A(n1421), .Y(n1377) );
  OA22X1_RVT U1811 ( .A1(n1378), .A2(n1616), .A3(n1377), .A4(n1095), .Y(n1283)
         );
  AND2X1_RVT U1812 ( .A1(n1284), .A2(n1283), .Y(n1286) );
  NAND2X0_RVT U1813 ( .A1(n1325), .A2(n1582), .Y(n1285) );
  AND2X1_RVT U1814 ( .A1(n1286), .A2(n1285), .Y(n1955) );
  NAND2X0_RVT U1815 ( .A1(n1287), .A2(n1647), .Y(n1288) );
  AND2X1_RVT U1816 ( .A1(n1289), .A2(n1288), .Y(n2018) );
  OA22X1_RVT U1817 ( .A1(n1290), .A2(m6stg_step), .A3(n2018), .A4(n1652), .Y(
        n1861) );
  OA22X1_RVT U1818 ( .A1(n1485), .A2(n397), .A3(n1633), .A4(n257), .Y(n2016)
         );
  AO22X1_RVT U1819 ( .A1(n1579), .A2(m4stg_frac[25]), .A3(n1593), .A4(
        m4stg_frac[26]), .Y(n1292) );
  AO22X1_RVT U1820 ( .A1(n1573), .A2(m4stg_frac[24]), .A3(n1422), .A4(
        m4stg_frac[23]), .Y(n1291) );
  OR2X1_RVT U1821 ( .A1(n1292), .A2(n1291), .Y(n1388) );
  OA22X1_RVT U1822 ( .A1(n1616), .A2(n1387), .A3(n1095), .A4(n1388), .Y(n1295)
         );
  OA22X1_RVT U1823 ( .A1(n35), .A2(n1337), .A3(n1623), .A4(n1293), .Y(n1294)
         );
  NAND2X0_RVT U1824 ( .A1(n1295), .A2(n1294), .Y(n1887) );
  AOI22X1_RVT U1825 ( .A1(n1891), .A2(n1296), .A3(n1647), .A4(n1887), .Y(n2015) );
  NAND2X0_RVT U1826 ( .A1(n2016), .A2(n2015), .Y(n1297) );
  OA22X1_RVT U1827 ( .A1(n1298), .A2(m6stg_step), .A3(n1297), .A4(n1652), .Y(
        n1860) );
  NAND2X0_RVT U1828 ( .A1(n1891), .A2(n1299), .Y(n1301) );
  OA22X1_RVT U1829 ( .A1(n1493), .A2(n397), .A3(n1639), .A4(n257), .Y(n1300)
         );
  AND2X1_RVT U1830 ( .A1(n1301), .A2(n1300), .Y(n1311) );
  NAND2X0_RVT U1831 ( .A1(n1539), .A2(n1302), .Y(n1306) );
  AO22X1_RVT U1832 ( .A1(n1579), .A2(m4stg_frac[24]), .A3(n1593), .A4(
        m4stg_frac[25]), .Y(n1304) );
  AO22X1_RVT U1833 ( .A1(n1573), .A2(m4stg_frac[23]), .A3(n1422), .A4(
        m4stg_frac[22]), .Y(n1303) );
  OR2X1_RVT U1834 ( .A1(n1304), .A2(n1303), .Y(n1445) );
  INVX1_RVT U1835 ( .A(n1445), .Y(n1399) );
  OA22X1_RVT U1836 ( .A1(n1400), .A2(n1616), .A3(n1399), .A4(n1095), .Y(n1305)
         );
  AND2X1_RVT U1837 ( .A1(n1306), .A2(n1305), .Y(n1308) );
  NAND2X0_RVT U1838 ( .A1(n1350), .A2(n1582), .Y(n1307) );
  AND2X1_RVT U1839 ( .A1(n1308), .A2(n1307), .Y(n1954) );
  NAND2X0_RVT U1840 ( .A1(n1309), .A2(n1647), .Y(n1310) );
  AND2X1_RVT U1841 ( .A1(n1311), .A2(n1310), .Y(n2014) );
  OA22X1_RVT U1842 ( .A1(n1312), .A2(m6stg_step), .A3(n2014), .A4(n1652), .Y(
        n1859) );
  AO22X1_RVT U1843 ( .A1(n1651), .A2(n1505), .A3(n1891), .A4(n1313), .Y(n1320)
         );
  AO22X1_RVT U1844 ( .A1(n1579), .A2(m4stg_frac[23]), .A3(n1593), .A4(
        m4stg_frac[24]), .Y(n1315) );
  AO22X1_RVT U1845 ( .A1(n1573), .A2(m4stg_frac[22]), .A3(n1422), .A4(
        m4stg_frac[21]), .Y(n1314) );
  OR2X1_RVT U1846 ( .A1(n1315), .A2(n1314), .Y(n1458) );
  OA22X1_RVT U1847 ( .A1(n1616), .A2(n1409), .A3(n1095), .A4(n1458), .Y(n1318)
         );
  OA22X1_RVT U1848 ( .A1(n35), .A2(n1366), .A3(n1623), .A4(n1316), .Y(n1317)
         );
  NAND2X0_RVT U1849 ( .A1(n1318), .A2(n1317), .Y(n1960) );
  AO22X1_RVT U1850 ( .A1(n1916), .A2(n1645), .A3(n1647), .A4(n1960), .Y(n1319)
         );
  OR2X1_RVT U1851 ( .A1(n1320), .A2(n1319), .Y(n2013) );
  OA22X1_RVT U1852 ( .A1(n1321), .A2(m6stg_step), .A3(n2013), .A4(n1652), .Y(
        n1858) );
  NAND2X0_RVT U1853 ( .A1(n1891), .A2(n1322), .Y(n1324) );
  OA22X1_RVT U1854 ( .A1(n1650), .A2(n257), .A3(n1516), .A4(n397), .Y(n1323)
         );
  AND2X1_RVT U1855 ( .A1(n1324), .A2(n1323), .Y(n1335) );
  NAND2X0_RVT U1856 ( .A1(n1539), .A2(n1325), .Y(n1329) );
  AO22X1_RVT U1857 ( .A1(n1579), .A2(m4stg_frac[22]), .A3(n1593), .A4(
        m4stg_frac[23]), .Y(n1327) );
  AO22X1_RVT U1858 ( .A1(n1573), .A2(m4stg_frac[21]), .A3(n1422), .A4(
        m4stg_frac[20]), .Y(n1326) );
  OR2X1_RVT U1859 ( .A1(n1327), .A2(n1326), .Y(n1472) );
  INVX1_RVT U1860 ( .A(n1472), .Y(n1376) );
  OA22X1_RVT U1861 ( .A1(n1377), .A2(n1616), .A3(n1376), .A4(n1095), .Y(n1328)
         );
  AND2X1_RVT U1862 ( .A1(n1329), .A2(n1328), .Y(n1332) );
  NAND2X0_RVT U1863 ( .A1(n1330), .A2(n1582), .Y(n1331) );
  AND2X1_RVT U1864 ( .A1(n1332), .A2(n1331), .Y(n1961) );
  NAND2X0_RVT U1865 ( .A1(n1333), .A2(n1647), .Y(n1334) );
  AND2X1_RVT U1866 ( .A1(n1335), .A2(n1334), .Y(n2012) );
  OA22X1_RVT U1867 ( .A1(n1336), .A2(m6stg_step), .A3(n2012), .A4(n1652), .Y(
        n1857) );
  NAND2X0_RVT U1868 ( .A1(n1539), .A2(n1337), .Y(n1341) );
  AO22X1_RVT U1869 ( .A1(n1579), .A2(m4stg_frac[21]), .A3(n1593), .A4(
        m4stg_frac[22]), .Y(n1339) );
  AO22X1_RVT U1870 ( .A1(n1573), .A2(m4stg_frac[20]), .A3(n1422), .A4(
        m4stg_frac[19]), .Y(n1338) );
  OR2X1_RVT U1871 ( .A1(n1339), .A2(n1338), .Y(n1488) );
  INVX1_RVT U1872 ( .A(n1488), .Y(n1434) );
  OA22X1_RVT U1873 ( .A1(n1435), .A2(n1616), .A3(n1434), .A4(n1095), .Y(n1340)
         );
  AND2X1_RVT U1874 ( .A1(n1341), .A2(n1340), .Y(n1343) );
  NAND2X0_RVT U1875 ( .A1(n1387), .A2(n1582), .Y(n1342) );
  AND2X1_RVT U1876 ( .A1(n1343), .A2(n1342), .Y(n1965) );
  AO22X1_RVT U1877 ( .A1(m4stg_sh_cnt[4]), .A2(n1965), .A3(n1879), .A4(n1528), 
        .Y(n1951) );
  INVX1_RVT U1878 ( .A(n1344), .Y(n1345) );
  OA222X1_RVT U1879 ( .A1(n2069), .A2(n1951), .A3(n397), .A4(n1527), .A5(n1632), .A6(n1345), .Y(n2011) );
  OA22X1_RVT U1880 ( .A1(n1346), .A2(m6stg_step), .A3(n2011), .A4(n1652), .Y(
        n1856) );
  NAND2X0_RVT U1881 ( .A1(n1891), .A2(n1347), .Y(n1349) );
  OA22X1_RVT U1882 ( .A1(n1888), .A2(n257), .A3(n1537), .A4(n397), .Y(n1348)
         );
  AND2X1_RVT U1883 ( .A1(n1349), .A2(n1348), .Y(n1360) );
  NAND2X0_RVT U1884 ( .A1(n1539), .A2(n1350), .Y(n1354) );
  AO22X1_RVT U1885 ( .A1(n1579), .A2(m4stg_frac[20]), .A3(n1593), .A4(
        m4stg_frac[21]), .Y(n1352) );
  AO22X1_RVT U1886 ( .A1(n1573), .A2(m4stg_frac[19]), .A3(n1422), .A4(
        m4stg_frac[18]), .Y(n1351) );
  OR2X1_RVT U1887 ( .A1(n1352), .A2(n1351), .Y(n1494) );
  INVX1_RVT U1888 ( .A(n1494), .Y(n1398) );
  OA22X1_RVT U1889 ( .A1(n1399), .A2(n1616), .A3(n1398), .A4(n1095), .Y(n1353)
         );
  AND2X1_RVT U1890 ( .A1(n1354), .A2(n1353), .Y(n1357) );
  NAND2X0_RVT U1891 ( .A1(n1355), .A2(n1582), .Y(n1356) );
  AND2X1_RVT U1892 ( .A1(n1357), .A2(n1356), .Y(n1964) );
  INVX1_RVT U1893 ( .A(n1964), .Y(n1358) );
  NAND2X0_RVT U1894 ( .A1(n1358), .A2(n1647), .Y(n1359) );
  AND2X1_RVT U1895 ( .A1(n1360), .A2(n1359), .Y(n2010) );
  OA22X1_RVT U1896 ( .A1(n1361), .A2(m6stg_step), .A3(n2010), .A4(n1652), .Y(
        n1855) );
  INVX1_RVT U1897 ( .A(n1362), .Y(n1550) );
  INVX1_RVT U1898 ( .A(n1363), .Y(n1369) );
  AO22X1_RVT U1899 ( .A1(n1579), .A2(m4stg_frac[19]), .A3(n1593), .A4(
        m4stg_frac[20]), .Y(n1365) );
  AO22X1_RVT U1900 ( .A1(n1573), .A2(m4stg_frac[18]), .A3(n1422), .A4(
        m4stg_frac[17]), .Y(n1364) );
  OR2X1_RVT U1901 ( .A1(n1365), .A2(n1364), .Y(n1509) );
  OA22X1_RVT U1902 ( .A1(n1616), .A2(n1458), .A3(n1095), .A4(n1509), .Y(n1368)
         );
  OA22X1_RVT U1903 ( .A1(n35), .A2(n1409), .A3(n1366), .A4(n1623), .Y(n1367)
         );
  NAND2X0_RVT U1904 ( .A1(n1368), .A2(n1367), .Y(n1959) );
  AO22X1_RVT U1905 ( .A1(m4stg_sh_cnt[4]), .A2(n1959), .A3(n1879), .A4(n1549), 
        .Y(n1882) );
  AO222X1_RVT U1906 ( .A1(n1550), .A2(n1651), .A3(n1369), .A4(n1891), .A5(
        n1882), .A6(\m4stg_sh_cnt_5[0] ), .Y(n2009) );
  OA22X1_RVT U1907 ( .A1(n1370), .A2(m6stg_step), .A3(n2009), .A4(n1652), .Y(
        n1854) );
  NAND2X0_RVT U1908 ( .A1(n1891), .A2(n1371), .Y(n1373) );
  OA22X1_RVT U1909 ( .A1(n1904), .A2(n257), .A3(n1558), .A4(n397), .Y(n1372)
         );
  AND2X1_RVT U1910 ( .A1(n1373), .A2(n1372), .Y(n1382) );
  AO22X1_RVT U1911 ( .A1(n1579), .A2(m4stg_frac[18]), .A3(n1593), .A4(
        m4stg_frac[19]), .Y(n1375) );
  AO22X1_RVT U1912 ( .A1(n1573), .A2(m4stg_frac[17]), .A3(n1422), .A4(
        m4stg_frac[16]), .Y(n1374) );
  OR2X1_RVT U1913 ( .A1(n1375), .A2(n1374), .Y(n1517) );
  INVX1_RVT U1914 ( .A(n1517), .Y(n1478) );
  OA22X1_RVT U1915 ( .A1(n1376), .A2(n1616), .A3(n1478), .A4(n1095), .Y(n1380)
         );
  OA22X1_RVT U1916 ( .A1(n1378), .A2(n1623), .A3(n1377), .A4(n35), .Y(n1379)
         );
  NAND2X0_RVT U1917 ( .A1(n1380), .A2(n1379), .Y(n1941) );
  NAND2X0_RVT U1918 ( .A1(n1941), .A2(n1647), .Y(n1381) );
  AND2X1_RVT U1919 ( .A1(n1382), .A2(n1381), .Y(n2008) );
  OA22X1_RVT U1920 ( .A1(n1383), .A2(m6stg_step), .A3(n2008), .A4(n1652), .Y(
        n1853) );
  OA22X1_RVT U1921 ( .A1(n1384), .A2(n1632), .A3(n1571), .A4(n397), .Y(n2007)
         );
  AO22X1_RVT U1922 ( .A1(n1579), .A2(m4stg_frac[17]), .A3(n1593), .A4(
        m4stg_frac[18]), .Y(n1386) );
  AO22X1_RVT U1923 ( .A1(n1573), .A2(m4stg_frac[16]), .A3(n1422), .A4(
        m4stg_frac[15]), .Y(n1385) );
  OR2X1_RVT U1924 ( .A1(n1386), .A2(n1385), .Y(n1531) );
  OA22X1_RVT U1925 ( .A1(n1616), .A2(n1488), .A3(n1095), .A4(n1531), .Y(n1390)
         );
  OA22X1_RVT U1926 ( .A1(n35), .A2(n1388), .A3(n1623), .A4(n1387), .Y(n1389)
         );
  NAND2X0_RVT U1927 ( .A1(n1390), .A2(n1389), .Y(n1958) );
  AOI22X1_RVT U1928 ( .A1(n1916), .A2(n1901), .A3(n1647), .A4(n1958), .Y(n2006) );
  NAND2X0_RVT U1929 ( .A1(n2007), .A2(n2006), .Y(n1391) );
  OA22X1_RVT U1930 ( .A1(n1392), .A2(m6stg_step), .A3(n1391), .A4(n1652), .Y(
        n1852) );
  NAND2X0_RVT U1931 ( .A1(n1891), .A2(n1393), .Y(n1395) );
  OA22X1_RVT U1932 ( .A1(n1903), .A2(n257), .A3(n1577), .A4(n397), .Y(n1394)
         );
  AND2X1_RVT U1933 ( .A1(n1395), .A2(n1394), .Y(n1404) );
  AO22X1_RVT U1934 ( .A1(n1579), .A2(m4stg_frac[16]), .A3(n1593), .A4(
        m4stg_frac[17]), .Y(n1397) );
  AO22X1_RVT U1935 ( .A1(n1573), .A2(m4stg_frac[15]), .A3(n1422), .A4(
        m4stg_frac[14]), .Y(n1396) );
  OR2X1_RVT U1936 ( .A1(n1397), .A2(n1396), .Y(n1538) );
  INVX1_RVT U1937 ( .A(n1538), .Y(n1448) );
  OA22X1_RVT U1938 ( .A1(n1398), .A2(n1616), .A3(n1448), .A4(n1095), .Y(n1402)
         );
  OA22X1_RVT U1939 ( .A1(n1400), .A2(n1623), .A3(n1399), .A4(n35), .Y(n1401)
         );
  NAND2X0_RVT U1940 ( .A1(n1402), .A2(n1401), .Y(n1940) );
  NAND2X0_RVT U1941 ( .A1(n1940), .A2(n1647), .Y(n1403) );
  AND2X1_RVT U1942 ( .A1(n1404), .A2(n1403), .Y(n2005) );
  OA22X1_RVT U1943 ( .A1(n1405), .A2(m6stg_step), .A3(n2005), .A4(n1652), .Y(
        n1851) );
  NAND2X0_RVT U1944 ( .A1(n1651), .A2(n1590), .Y(n1408) );
  OA22X1_RVT U1945 ( .A1(n1902), .A2(n257), .A3(n1406), .A4(n1632), .Y(n1407)
         );
  AND2X1_RVT U1946 ( .A1(n1408), .A2(n1407), .Y(n1419) );
  NAND2X0_RVT U1947 ( .A1(n1539), .A2(n1409), .Y(n1414) );
  AO22X1_RVT U1948 ( .A1(n1579), .A2(m4stg_frac[15]), .A3(n1593), .A4(
        m4stg_frac[16]), .Y(n1411) );
  AO22X1_RVT U1949 ( .A1(n1573), .A2(m4stg_frac[14]), .A3(n1422), .A4(
        m4stg_frac[13]), .Y(n1410) );
  OR2X1_RVT U1950 ( .A1(n1411), .A2(n1410), .Y(n1510) );
  INVX1_RVT U1951 ( .A(n1510), .Y(n1554) );
  OA22X1_RVT U1952 ( .A1(n1412), .A2(n1616), .A3(n1554), .A4(n1095), .Y(n1413)
         );
  AND2X1_RVT U1953 ( .A1(n1414), .A2(n1413), .Y(n1416) );
  NAND2X0_RVT U1954 ( .A1(n1458), .A2(n1582), .Y(n1415) );
  AND2X1_RVT U1955 ( .A1(n1416), .A2(n1415), .Y(n1936) );
  INVX1_RVT U1956 ( .A(n1936), .Y(n1417) );
  NAND2X0_RVT U1957 ( .A1(n1417), .A2(n1647), .Y(n1418) );
  AND2X1_RVT U1958 ( .A1(n1419), .A2(n1418), .Y(n2004) );
  OA22X1_RVT U1959 ( .A1(n1420), .A2(m6stg_step), .A3(n2004), .A4(n1652), .Y(
        n1850) );
  NAND2X0_RVT U1960 ( .A1(n1539), .A2(n1421), .Y(n1426) );
  AO22X1_RVT U1961 ( .A1(n1579), .A2(m4stg_frac[14]), .A3(n1593), .A4(
        m4stg_frac[15]), .Y(n1424) );
  AO22X1_RVT U1962 ( .A1(n1573), .A2(m4stg_frac[13]), .A3(n1422), .A4(
        m4stg_frac[12]), .Y(n1423) );
  OR2X1_RVT U1963 ( .A1(n1424), .A2(n1423), .Y(n1559) );
  INVX1_RVT U1964 ( .A(n1559), .Y(n1475) );
  OA22X1_RVT U1965 ( .A1(n1478), .A2(n1616), .A3(n1475), .A4(n1095), .Y(n1425)
         );
  AND2X1_RVT U1966 ( .A1(n1426), .A2(n1425), .Y(n1428) );
  NAND2X0_RVT U1967 ( .A1(n1472), .A2(n1582), .Y(n1427) );
  AND2X1_RVT U1968 ( .A1(n1428), .A2(n1427), .Y(n1937) );
  AO22X1_RVT U1969 ( .A1(m4stg_sh_cnt[4]), .A2(n1937), .A3(n1879), .A4(n1601), 
        .Y(n1950) );
  OA222X1_RVT U1970 ( .A1(n2069), .A2(n1950), .A3(n397), .A4(n1600), .A5(n1632), .A6(n1430), .Y(n2003) );
  OA22X1_RVT U1971 ( .A1(n1431), .A2(m6stg_step), .A3(n2003), .A4(n1652), .Y(
        n1849) );
  AO22X1_RVT U1972 ( .A1(n1579), .A2(m4stg_frac[13]), .A3(n1593), .A4(
        m4stg_frac[14]), .Y(n1433) );
  AO22X1_RVT U1973 ( .A1(n1573), .A2(m4stg_frac[12]), .A3(n1422), .A4(
        m4stg_frac[11]), .Y(n1432) );
  OR2X1_RVT U1974 ( .A1(n1433), .A2(n1432), .Y(n1574) );
  AOI22X1_RVT U1975 ( .A1(n1531), .A2(n1268), .A3(n1574), .A4(n6), .Y(n1437)
         );
  OA22X1_RVT U1976 ( .A1(n1435), .A2(n1623), .A3(n1434), .A4(n35), .Y(n1436)
         );
  NAND2X0_RVT U1977 ( .A1(n1437), .A2(n1436), .Y(n1889) );
  INVX1_RVT U1978 ( .A(n1889), .Y(n1611) );
  AO22X1_RVT U1979 ( .A1(m4stg_sh_cnt[4]), .A2(n1611), .A3(n1879), .A4(n1607), 
        .Y(n1924) );
  INVX1_RVT U1980 ( .A(n1438), .Y(n1439) );
  OA222X1_RVT U1981 ( .A1(n2069), .A2(n1924), .A3(n397), .A4(n1606), .A5(n1632), .A6(n1439), .Y(n2002) );
  OA22X1_RVT U1982 ( .A1(n1440), .A2(m6stg_step), .A3(n2002), .A4(n1652), .Y(
        n1848) );
  NAND2X0_RVT U1983 ( .A1(n1891), .A2(n1441), .Y(n1444) );
  OA22X1_RVT U1984 ( .A1(n1957), .A2(n257), .A3(n1615), .A4(n397), .Y(n1443)
         );
  AND2X1_RVT U1985 ( .A1(n1444), .A2(n1443), .Y(n1455) );
  NAND2X0_RVT U1986 ( .A1(n1539), .A2(n1445), .Y(n1450) );
  AO22X1_RVT U1987 ( .A1(n1579), .A2(m4stg_frac[12]), .A3(n1593), .A4(
        m4stg_frac[13]), .Y(n1447) );
  AO22X1_RVT U1988 ( .A1(n1573), .A2(m4stg_frac[11]), .A3(n1422), .A4(
        m4stg_frac[10]), .Y(n1446) );
  OR2X1_RVT U1989 ( .A1(n1447), .A2(n1446), .Y(n1578) );
  INVX1_RVT U1990 ( .A(n1578), .Y(n1497) );
  OA22X1_RVT U1991 ( .A1(n1497), .A2(n1095), .A3(n1448), .A4(n1616), .Y(n1449)
         );
  AND2X1_RVT U1992 ( .A1(n1450), .A2(n1449), .Y(n1452) );
  NAND2X0_RVT U1993 ( .A1(n1494), .A2(n1582), .Y(n1451) );
  AND2X1_RVT U1994 ( .A1(n1452), .A2(n1451), .Y(n1935) );
  INVX1_RVT U1995 ( .A(n1935), .Y(n1453) );
  NAND2X0_RVT U1996 ( .A1(n1453), .A2(n1647), .Y(n1454) );
  AND2X1_RVT U1997 ( .A1(n1455), .A2(n1454), .Y(n2001) );
  OA22X1_RVT U1998 ( .A1(n1456), .A2(m6stg_step), .A3(n2001), .A4(n1652), .Y(
        n1847) );
  OA22X1_RVT U1999 ( .A1(n1457), .A2(n1632), .A3(n1621), .A4(n397), .Y(n1466)
         );
  NAND2X0_RVT U2000 ( .A1(n1539), .A2(n1458), .Y(n1462) );
  AO22X1_RVT U2001 ( .A1(n1579), .A2(m4stg_frac[11]), .A3(n1593), .A4(
        m4stg_frac[12]), .Y(n1460) );
  AO22X1_RVT U2002 ( .A1(n1573), .A2(m4stg_frac[10]), .A3(n1422), .A4(
        m4stg_frac[9]), .Y(n1459) );
  OR2X1_RVT U2003 ( .A1(n1460), .A2(n1459), .Y(n1508) );
  INVX1_RVT U2004 ( .A(n1508), .Y(n1595) );
  OA22X1_RVT U2005 ( .A1(n1595), .A2(n1095), .A3(n1554), .A4(n1616), .Y(n1461)
         );
  AND2X1_RVT U2006 ( .A1(n1462), .A2(n1461), .Y(n1464) );
  NAND2X0_RVT U2007 ( .A1(n1509), .A2(n1582), .Y(n1463) );
  AND2X1_RVT U2008 ( .A1(n1464), .A2(n1463), .Y(n1934) );
  OA22X1_RVT U2009 ( .A1(n1934), .A2(n1625), .A3(n1956), .A4(n257), .Y(n1465)
         );
  AND2X1_RVT U2010 ( .A1(n1466), .A2(n1465), .Y(n2000) );
  OA22X1_RVT U2011 ( .A1(n1467), .A2(m6stg_step), .A3(n2000), .A4(n1652), .Y(
        n1846) );
  NAND2X0_RVT U2012 ( .A1(n1891), .A2(n1468), .Y(n1471) );
  OA22X1_RVT U2013 ( .A1(n1955), .A2(n257), .A3(n1630), .A4(n397), .Y(n1470)
         );
  AND2X1_RVT U2014 ( .A1(n1471), .A2(n1470), .Y(n1483) );
  NAND2X0_RVT U2015 ( .A1(n1539), .A2(n1472), .Y(n1477) );
  AO22X1_RVT U2016 ( .A1(n1579), .A2(m4stg_frac[10]), .A3(n1593), .A4(
        m4stg_frac[11]), .Y(n1474) );
  AO22X1_RVT U2017 ( .A1(n1573), .A2(m4stg_frac[9]), .A3(n1422), .A4(
        m4stg_frac[8]), .Y(n1473) );
  NOR2X0_RVT U2018 ( .A1(n1474), .A2(n1473), .Y(n1602) );
  OA22X1_RVT U2019 ( .A1(n1475), .A2(n1616), .A3(n1602), .A4(n1095), .Y(n1476)
         );
  AND2X1_RVT U2020 ( .A1(n1477), .A2(n1476), .Y(n1480) );
  NAND2X0_RVT U2021 ( .A1(n1517), .A2(n1582), .Y(n1479) );
  AND2X1_RVT U2022 ( .A1(n1480), .A2(n1479), .Y(n1931) );
  INVX1_RVT U2023 ( .A(n1931), .Y(n1481) );
  NAND2X0_RVT U2024 ( .A1(n1481), .A2(n1647), .Y(n1482) );
  AND2X1_RVT U2025 ( .A1(n1483), .A2(n1482), .Y(n1999) );
  OA22X1_RVT U2026 ( .A1(n1484), .A2(m6stg_step), .A3(n1999), .A4(n1652), .Y(
        n1845) );
  OA22X1_RVT U2027 ( .A1(n1485), .A2(n1632), .A3(n1633), .A4(n397), .Y(n1998)
         );
  AO22X1_RVT U2028 ( .A1(n1579), .A2(m4stg_frac[9]), .A3(n1593), .A4(
        m4stg_frac[10]), .Y(n1487) );
  AO22X1_RVT U2029 ( .A1(n1573), .A2(m4stg_frac[8]), .A3(n1422), .A4(
        m4stg_frac[7]), .Y(n1486) );
  OR2X1_RVT U2030 ( .A1(n1487), .A2(n1486), .Y(n1608) );
  OA22X1_RVT U2031 ( .A1(n1616), .A2(n1574), .A3(n1095), .A4(n1608), .Y(n1490)
         );
  OA22X1_RVT U2032 ( .A1(n35), .A2(n1531), .A3(n1623), .A4(n1488), .Y(n1489)
         );
  NAND2X0_RVT U2033 ( .A1(n1490), .A2(n1489), .Y(n1881) );
  AOI22X1_RVT U2034 ( .A1(n1916), .A2(n1887), .A3(n1647), .A4(n1881), .Y(n1997) );
  NAND2X0_RVT U2035 ( .A1(n1998), .A2(n1997), .Y(n1491) );
  OA22X1_RVT U2036 ( .A1(n1492), .A2(m6stg_step), .A3(n1491), .A4(n1652), .Y(
        n1844) );
  OA22X1_RVT U2037 ( .A1(n1493), .A2(n1632), .A3(n1639), .A4(n397), .Y(n1503)
         );
  NAND2X0_RVT U2038 ( .A1(n1539), .A2(n1494), .Y(n1499) );
  AO22X1_RVT U2039 ( .A1(n1579), .A2(m4stg_frac[8]), .A3(n1593), .A4(
        m4stg_frac[9]), .Y(n1496) );
  AO22X1_RVT U2040 ( .A1(n1573), .A2(m4stg_frac[7]), .A3(n1422), .A4(
        m4stg_frac[6]), .Y(n1495) );
  NOR2X0_RVT U2041 ( .A1(n1496), .A2(n1495), .Y(n1617) );
  OA22X1_RVT U2042 ( .A1(n1617), .A2(n1095), .A3(n1497), .A4(n1616), .Y(n1498)
         );
  AND2X1_RVT U2043 ( .A1(n1499), .A2(n1498), .Y(n1501) );
  NAND2X0_RVT U2044 ( .A1(n1538), .A2(n1582), .Y(n1500) );
  AND2X1_RVT U2045 ( .A1(n1501), .A2(n1500), .Y(n1930) );
  OA22X1_RVT U2046 ( .A1(n1930), .A2(n1625), .A3(n1954), .A4(n257), .Y(n1502)
         );
  AND2X1_RVT U2047 ( .A1(n1503), .A2(n1502), .Y(n1996) );
  OA22X1_RVT U2048 ( .A1(n1504), .A2(m6stg_step), .A3(n1996), .A4(n1652), .Y(
        n1843) );
  AO22X1_RVT U2049 ( .A1(n1651), .A2(n1645), .A3(n1891), .A4(n1505), .Y(n1514)
         );
  AO22X1_RVT U2050 ( .A1(n1579), .A2(m4stg_frac[7]), .A3(n1593), .A4(
        m4stg_frac[8]), .Y(n1507) );
  AO22X1_RVT U2051 ( .A1(n1573), .A2(m4stg_frac[6]), .A3(n1422), .A4(
        m4stg_frac[5]), .Y(n1506) );
  OR2X1_RVT U2052 ( .A1(n1507), .A2(n1506), .Y(n1551) );
  OA22X1_RVT U2053 ( .A1(n1616), .A2(n1508), .A3(n1095), .A4(n1551), .Y(n1512)
         );
  OA22X1_RVT U2054 ( .A1(n35), .A2(n1510), .A3(n1623), .A4(n1509), .Y(n1511)
         );
  NAND2X0_RVT U2055 ( .A1(n1512), .A2(n1511), .Y(n1929) );
  AO22X1_RVT U2056 ( .A1(n1647), .A2(n1929), .A3(n1916), .A4(n1960), .Y(n1513)
         );
  OR2X1_RVT U2057 ( .A1(n1514), .A2(n1513), .Y(n1995) );
  OA22X1_RVT U2058 ( .A1(n1515), .A2(m6stg_step), .A3(n1995), .A4(n1652), .Y(
        n1842) );
  OA22X1_RVT U2059 ( .A1(n1650), .A2(n397), .A3(n1516), .A4(n1632), .Y(n1525)
         );
  NAND2X0_RVT U2060 ( .A1(n1539), .A2(n1517), .Y(n1521) );
  AO22X1_RVT U2061 ( .A1(n1579), .A2(m4stg_frac[6]), .A3(n1593), .A4(
        m4stg_frac[7]), .Y(n1519) );
  AO22X1_RVT U2062 ( .A1(n1573), .A2(m4stg_frac[5]), .A3(n1422), .A4(
        m4stg_frac[4]), .Y(n1518) );
  NOR2X0_RVT U2063 ( .A1(n1519), .A2(n1518), .Y(n1907) );
  OA22X1_RVT U2064 ( .A1(n1602), .A2(n1616), .A3(n1907), .A4(n1095), .Y(n1520)
         );
  AND2X1_RVT U2065 ( .A1(n1521), .A2(n1520), .Y(n1523) );
  NAND2X0_RVT U2066 ( .A1(n1559), .A2(n1582), .Y(n1522) );
  AND2X1_RVT U2067 ( .A1(n1523), .A2(n1522), .Y(n1932) );
  OA22X1_RVT U2068 ( .A1(n1932), .A2(n1625), .A3(n1961), .A4(n257), .Y(n1524)
         );
  AND2X1_RVT U2069 ( .A1(n1525), .A2(n1524), .Y(n1994) );
  OA22X1_RVT U2070 ( .A1(n1526), .A2(m6stg_step), .A3(n1994), .A4(n1652), .Y(
        n1841) );
  OA22X1_RVT U2071 ( .A1(n1528), .A2(n397), .A3(n1527), .A4(n1632), .Y(n1535)
         );
  AO22X1_RVT U2072 ( .A1(n1579), .A2(m4stg_frac[5]), .A3(n1593), .A4(
        m4stg_frac[6]), .Y(n1530) );
  AO22X1_RVT U2073 ( .A1(n1573), .A2(m4stg_frac[4]), .A3(n1422), .A4(
        m4stg_frac[3]), .Y(n1529) );
  OR2X1_RVT U2074 ( .A1(n1530), .A2(n1529), .Y(n1609) );
  AO22X1_RVT U2075 ( .A1(n1268), .A2(n1608), .A3(n6), .A4(n1609), .Y(n1533) );
  AO22X1_RVT U2076 ( .A1(n1582), .A2(n1574), .A3(n1539), .A4(n1531), .Y(n1532)
         );
  OR2X1_RVT U2077 ( .A1(n1533), .A2(n1532), .Y(n1654) );
  INVX1_RVT U2078 ( .A(n1654), .Y(n1945) );
  OA22X1_RVT U2079 ( .A1(n1945), .A2(n1625), .A3(n1965), .A4(n257), .Y(n1534)
         );
  AND2X1_RVT U2080 ( .A1(n1535), .A2(n1534), .Y(n1993) );
  OA22X1_RVT U2081 ( .A1(n1536), .A2(m6stg_step), .A3(n1993), .A4(n1652), .Y(
        n1840) );
  OA22X1_RVT U2082 ( .A1(n1888), .A2(n397), .A3(n1537), .A4(n1632), .Y(n1547)
         );
  NAND2X0_RVT U2083 ( .A1(n1539), .A2(n1538), .Y(n1543) );
  AO22X1_RVT U2084 ( .A1(n1579), .A2(m4stg_frac[4]), .A3(n1593), .A4(
        m4stg_frac[5]), .Y(n1541) );
  AO22X1_RVT U2085 ( .A1(n1573), .A2(m4stg_frac[3]), .A3(n1422), .A4(
        m4stg_frac[2]), .Y(n1540) );
  NOR2X0_RVT U2086 ( .A1(n1541), .A2(n1540), .Y(n1640) );
  OA22X1_RVT U2087 ( .A1(n1640), .A2(n1095), .A3(n1617), .A4(n1616), .Y(n1542)
         );
  AND2X1_RVT U2088 ( .A1(n1543), .A2(n1542), .Y(n1545) );
  NAND2X0_RVT U2089 ( .A1(n1578), .A2(n1582), .Y(n1544) );
  AND2X1_RVT U2090 ( .A1(n1545), .A2(n1544), .Y(n1944) );
  OA22X1_RVT U2091 ( .A1(n1944), .A2(n1625), .A3(n1964), .A4(n257), .Y(n1546)
         );
  AND2X1_RVT U2092 ( .A1(n1547), .A2(n1546), .Y(n1992) );
  OA22X1_RVT U2093 ( .A1(n1548), .A2(m6stg_step), .A3(n1992), .A4(n1652), .Y(
        n1839) );
  AO22X1_RVT U2094 ( .A1(n1891), .A2(n1550), .A3(n1651), .A4(n1549), .Y(n1556)
         );
  INVX1_RVT U2095 ( .A(n1551), .Y(n1622) );
  AO22X1_RVT U2096 ( .A1(n1579), .A2(m4stg_frac[3]), .A3(n1593), .A4(
        m4stg_frac[4]), .Y(n1553) );
  AO22X1_RVT U2097 ( .A1(n1573), .A2(m4stg_frac[2]), .A3(n1422), .A4(
        m4stg_frac[1]), .Y(n1552) );
  NOR2X0_RVT U2098 ( .A1(n1553), .A2(n1552), .Y(n1624) );
  MUX41X1_RVT U2099 ( .A1(n1554), .A3(n1595), .A2(n1622), .A4(n1624), .S0(
        m4stg_sh_cnt[2]), .S1(m4stg_sh_cnt[3]), .Y(n1926) );
  AO22X1_RVT U2100 ( .A1(n1647), .A2(n1926), .A3(n1916), .A4(n1959), .Y(n1555)
         );
  OR2X1_RVT U2101 ( .A1(n1556), .A2(n1555), .Y(n1991) );
  OA22X1_RVT U2102 ( .A1(n1557), .A2(m6stg_step), .A3(n1991), .A4(n1652), .Y(
        n1838) );
  OA22X1_RVT U2103 ( .A1(n1904), .A2(n397), .A3(n1558), .A4(n1632), .Y(n1569)
         );
  NAND2X0_RVT U2104 ( .A1(n1539), .A2(n1559), .Y(n1563) );
  AO22X1_RVT U2105 ( .A1(n1422), .A2(m4stg_frac[0]), .A3(n1593), .A4(
        m4stg_frac[3]), .Y(n1561) );
  AO22X1_RVT U2106 ( .A1(n1573), .A2(m4stg_frac[1]), .A3(n1579), .A4(
        m4stg_frac[2]), .Y(n1560) );
  OR2X1_RVT U2107 ( .A1(n1561), .A2(n1560), .Y(n1886) );
  INVX1_RVT U2108 ( .A(n1886), .Y(n1909) );
  OA22X1_RVT U2109 ( .A1(n1909), .A2(n1095), .A3(n1907), .A4(n1616), .Y(n1562)
         );
  AND2X1_RVT U2110 ( .A1(n1563), .A2(n1562), .Y(n1566) );
  NAND2X0_RVT U2111 ( .A1(n1564), .A2(n1582), .Y(n1565) );
  AND2X1_RVT U2112 ( .A1(n1566), .A2(n1565), .Y(n1896) );
  OA22X1_RVT U2113 ( .A1(n1896), .A2(n1625), .A3(n1567), .A4(n257), .Y(n1568)
         );
  AND2X1_RVT U2114 ( .A1(n1569), .A2(n1568), .Y(n1990) );
  OA22X1_RVT U2115 ( .A1(n1570), .A2(m6stg_step), .A3(n1990), .A4(n1652), .Y(
        n1837) );
  OA22X1_RVT U2116 ( .A1(n1572), .A2(n397), .A3(n1571), .A4(n1632), .Y(n1989)
         );
  AO222X1_RVT U2117 ( .A1(n1573), .A2(m4stg_frac[0]), .A3(n1593), .A4(
        m4stg_frac[2]), .A5(n1579), .A6(m4stg_frac[1]), .Y(n1897) );
  AO22X1_RVT U2118 ( .A1(m4stg_sh_cnt[2]), .A2(n1897), .A3(n1908), .A4(n1609), 
        .Y(n1635) );
  OAI222X1_RVT U2119 ( .A1(n1636), .A2(n1635), .A3(n1623), .A4(n1574), .A5(n35), .A6(n1608), .Y(n1880) );
  AOI22X1_RVT U2120 ( .A1(n1647), .A2(n1880), .A3(n1916), .A4(n1958), .Y(n1988) );
  NAND2X0_RVT U2121 ( .A1(n1989), .A2(n1988), .Y(n1575) );
  OA22X1_RVT U2122 ( .A1(n1576), .A2(m6stg_step), .A3(n1575), .A4(n1652), .Y(
        n1836) );
  OA22X1_RVT U2123 ( .A1(n1903), .A2(n397), .A3(n1577), .A4(n1632), .Y(n1588)
         );
  NAND2X0_RVT U2124 ( .A1(n1539), .A2(n1578), .Y(n1581) );
  AO22X1_RVT U2125 ( .A1(n1579), .A2(m4stg_frac[0]), .A3(n1593), .A4(
        m4stg_frac[1]), .Y(n1893) );
  INVX1_RVT U2126 ( .A(n1893), .Y(n1641) );
  OA22X1_RVT U2127 ( .A1(n1641), .A2(n1095), .A3(n1640), .A4(n1616), .Y(n1580)
         );
  AND2X1_RVT U2128 ( .A1(n1581), .A2(n1580), .Y(n1585) );
  NAND2X0_RVT U2129 ( .A1(n1583), .A2(n1582), .Y(n1584) );
  AND2X1_RVT U2130 ( .A1(n1585), .A2(n1584), .Y(n1659) );
  OA22X1_RVT U2131 ( .A1(n1586), .A2(n257), .A3(n1659), .A4(n1625), .Y(n1587)
         );
  AND2X1_RVT U2132 ( .A1(n1588), .A2(n1587), .Y(n1987) );
  OA22X1_RVT U2133 ( .A1(n1589), .A2(m6stg_step), .A3(n1987), .A4(n1652), .Y(
        n1835) );
  NAND2X0_RVT U2134 ( .A1(n1891), .A2(n1590), .Y(n1592) );
  OA22X1_RVT U2135 ( .A1(n1936), .A2(n257), .A3(n1902), .A4(n397), .Y(n1591)
         );
  AND2X1_RVT U2136 ( .A1(n1592), .A2(n1591), .Y(n1598) );
  NAND2X0_RVT U2137 ( .A1(n1593), .A2(m4stg_frac[0]), .Y(n1594) );
  AO22X1_RVT U2138 ( .A1(m4stg_sh_cnt[2]), .A2(n1594), .A3(n1908), .A4(n1624), 
        .Y(n1923) );
  OA222X1_RVT U2139 ( .A1(n1636), .A2(n1923), .A3(n35), .A4(n1622), .A5(n1623), 
        .A6(n1595), .Y(n1658) );
  INVX1_RVT U2140 ( .A(n1658), .Y(n1596) );
  NAND2X0_RVT U2141 ( .A1(n1596), .A2(n1647), .Y(n1597) );
  AND2X1_RVT U2142 ( .A1(n1598), .A2(n1597), .Y(n1986) );
  OA22X1_RVT U2143 ( .A1(n1599), .A2(m6stg_step), .A3(n1986), .A4(n1652), .Y(
        n1834) );
  OA22X1_RVT U2144 ( .A1(n1601), .A2(n397), .A3(n1600), .A4(n1632), .Y(n1604)
         );
  OA222X1_RVT U2145 ( .A1(n35), .A2(n1907), .A3(n1623), .A4(n1602), .A5(n1616), 
        .A6(n1909), .Y(n1895) );
  OA22X1_RVT U2146 ( .A1(n1895), .A2(n1625), .A3(n1937), .A4(n257), .Y(n1603)
         );
  AND2X1_RVT U2147 ( .A1(n1604), .A2(n1603), .Y(n1985) );
  OA22X1_RVT U2148 ( .A1(n1605), .A2(m6stg_step), .A3(n1985), .A4(n1652), .Y(
        n1833) );
  OA22X1_RVT U2149 ( .A1(n1607), .A2(n397), .A3(n1606), .A4(n1632), .Y(n1613)
         );
  AO22X1_RVT U2150 ( .A1(m4stg_sh_cnt[2]), .A2(n1609), .A3(n1908), .A4(n1608), 
        .Y(n1610) );
  AO22X1_RVT U2151 ( .A1(n1268), .A2(n1897), .A3(n1610), .A4(n1636), .Y(n1915)
         );
  INVX1_RVT U2152 ( .A(n1915), .Y(n1925) );
  OA22X1_RVT U2153 ( .A1(n1925), .A2(n1625), .A3(n1611), .A4(n257), .Y(n1612)
         );
  AND2X1_RVT U2154 ( .A1(n1613), .A2(n1612), .Y(n1984) );
  OA22X1_RVT U2155 ( .A1(n1614), .A2(m6stg_step), .A3(n1984), .A4(n1652), .Y(
        n1832) );
  OA22X1_RVT U2156 ( .A1(n1957), .A2(n397), .A3(n1615), .A4(n1632), .Y(n1619)
         );
  OA222X1_RVT U2157 ( .A1(n35), .A2(n1640), .A3(n1623), .A4(n1617), .A5(n1616), 
        .A6(n1641), .Y(n1657) );
  OA22X1_RVT U2158 ( .A1(n1935), .A2(n257), .A3(n1657), .A4(n1625), .Y(n1618)
         );
  AND2X1_RVT U2159 ( .A1(n1619), .A2(n1618), .Y(n1983) );
  OA22X1_RVT U2160 ( .A1(n1620), .A2(m6stg_step), .A3(n1983), .A4(n1652), .Y(
        n1831) );
  OA22X1_RVT U2161 ( .A1(n1956), .A2(n397), .A3(n1621), .A4(n1632), .Y(n1627)
         );
  NAND3X0_RVT U2162 ( .A1(n1593), .A2(m4stg_frac[0]), .A3(n1908), .Y(n1898) );
  OA222X1_RVT U2163 ( .A1(n1636), .A2(n1898), .A3(n35), .A4(n1624), .A5(n1623), 
        .A6(n1622), .Y(n1656) );
  OA22X1_RVT U2164 ( .A1(n1934), .A2(n257), .A3(n1656), .A4(n1625), .Y(n1626)
         );
  AND2X1_RVT U2165 ( .A1(n1627), .A2(n1626), .Y(n1982) );
  OA22X1_RVT U2166 ( .A1(n1628), .A2(m6stg_step), .A3(n1982), .A4(n1652), .Y(
        n1830) );
  AO222X1_RVT U2167 ( .A1(m4stg_sh_cnt[4]), .A2(n1909), .A3(m4stg_sh_cnt[4]), 
        .A4(n35), .A5(n1931), .A6(n1879), .Y(n1629) );
  OA21X1_RVT U2168 ( .A1(n1907), .A2(n1899), .A3(n1629), .Y(n1928) );
  OA222X1_RVT U2169 ( .A1(n2069), .A2(n1928), .A3(n1632), .A4(n1630), .A5(n397), .A6(n1955), .Y(n1981) );
  OA22X1_RVT U2170 ( .A1(n1631), .A2(m6stg_step), .A3(n1981), .A4(n1652), .Y(
        n1829) );
  OA22X1_RVT U2171 ( .A1(n1634), .A2(n397), .A3(n1633), .A4(n1632), .Y(n1980)
         );
  NAND2X0_RVT U2172 ( .A1(n1636), .A2(n1635), .Y(n1922) );
  AOI22X1_RVT U2173 ( .A1(n1916), .A2(n1881), .A3(n1647), .A4(n1922), .Y(n1979) );
  NAND2X0_RVT U2174 ( .A1(n1980), .A2(n1979), .Y(n1637) );
  OA22X1_RVT U2175 ( .A1(n1638), .A2(m6stg_step), .A3(n1637), .A4(n1652), .Y(
        n1828) );
  AO22X1_RVT U2176 ( .A1(n1954), .A2(n1651), .A3(n1891), .A4(n1639), .Y(n1643)
         );
  AO221X1_RVT U2177 ( .A1(m4stg_sh_cnt[2]), .A2(n1641), .A3(n1908), .A4(n1640), 
        .A5(m4stg_sh_cnt[3]), .Y(n1921) );
  AO22X1_RVT U2178 ( .A1(n1916), .A2(n1930), .A3(n1647), .A4(n1921), .Y(n1642)
         );
  OR2X1_RVT U2179 ( .A1(n1643), .A2(n1642), .Y(n1978) );
  OA22X1_RVT U2180 ( .A1(n1644), .A2(m6stg_step), .A3(n1978), .A4(n1652), .Y(
        n1827) );
  AO22X1_RVT U2181 ( .A1(n1891), .A2(n1645), .A3(n1651), .A4(n1960), .Y(n1646)
         );
  AO221X1_RVT U2182 ( .A1(n1647), .A2(m4stg_sh_cnt[3]), .A3(n1647), .A4(n1923), 
        .A5(n1646), .Y(n1648) );
  AO21X1_RVT U2183 ( .A1(n1916), .A2(n1929), .A3(n1648), .Y(n1977) );
  OA22X1_RVT U2184 ( .A1(m6stg_step), .A2(n1649), .A3(n1652), .A4(n1977), .Y(
        n1826) );
  OA22X1_RVT U2185 ( .A1(n1909), .A2(n1899), .A3(m4stg_sh_cnt[4]), .A4(n1932), 
        .Y(n1927) );
  AO222X1_RVT U2186 ( .A1(\m4stg_sh_cnt_5[0] ), .A2(n1927), .A3(n1961), .A4(
        n1651), .A5(n1891), .A6(n1650), .Y(n1976) );
  OA22X1_RVT U2187 ( .A1(m6stg_step), .A2(n1653), .A3(n1652), .A4(n1976), .Y(
        n1825) );
  NAND2X0_RVT U2188 ( .A1(n1879), .A2(n1654), .Y(n1655) );
  OA221X1_RVT U2189 ( .A1(n397), .A2(n1964), .A3(n397), .A4(n1958), .A5(n1655), 
        .Y(n1971) );
  NAND2X0_RVT U2190 ( .A1(n1657), .A2(n1656), .Y(n1939) );
  NAND2X0_RVT U2191 ( .A1(n1659), .A2(n1658), .Y(n1949) );
  AOI222X1_RVT U2192 ( .A1(n1879), .A2(n1939), .A3(n1879), .A4(n1949), .A5(
        n1879), .A6(n1660), .Y(n1970) );
  NAND3X0_RVT U2193 ( .A1(n1926), .A2(n1922), .A3(n1880), .Y(n1884) );
  NAND3X0_RVT U2194 ( .A1(n1882), .A2(n1881), .A3(n1880), .Y(n1883) );
  AO22X1_RVT U2195 ( .A1(n1916), .A2(n1884), .A3(n2069), .A4(n1883), .Y(n1920)
         );
  AO22X1_RVT U2196 ( .A1(n1894), .A2(n1886), .A3(n1885), .A4(n1893), .Y(n1919)
         );
  NAND2X0_RVT U2197 ( .A1(n1888), .A2(n1887), .Y(n1890) );
  AO22X1_RVT U2198 ( .A1(n1891), .A2(n1890), .A3(n2069), .A4(n1889), .Y(n1892)
         );
  AO221X1_RVT U2199 ( .A1(n1894), .A2(n1893), .A3(n1894), .A4(n1897), .A5(
        n1892), .Y(n1918) );
  NAND2X0_RVT U2200 ( .A1(n1896), .A2(n1895), .Y(n1933) );
  OA22X1_RVT U2201 ( .A1(n1900), .A2(n1899), .A3(m4stg_sh_cnt[3]), .A4(n1898), 
        .Y(n1913) );
  OA22X1_RVT U2202 ( .A1(m4stg_sh_cnt[4]), .A2(n1921), .A3(n1906), .A4(n1923), 
        .Y(n1912) );
  NAND4X0_RVT U2203 ( .A1(n1904), .A2(n1903), .A3(n1902), .A4(n1901), .Y(n1905) );
  NAND2X0_RVT U2204 ( .A1(n1891), .A2(n1905), .Y(n1911) );
  AO221X1_RVT U2205 ( .A1(m4stg_sh_cnt[2]), .A2(n1909), .A3(n1908), .A4(n1907), 
        .A5(n1906), .Y(n1910) );
  NAND4X0_RVT U2206 ( .A1(n1913), .A2(n1912), .A3(n1911), .A4(n1910), .Y(n1914) );
  AO221X1_RVT U2207 ( .A1(n1916), .A2(n1933), .A3(n1916), .A4(n1915), .A5(
        n1914), .Y(n1917) );
  NOR4X1_RVT U2208 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), .Y(n1969)
         );
  AND4X1_RVT U2209 ( .A1(n1924), .A2(n1923), .A3(n1922), .A4(n1921), .Y(n1953)
         );
  NAND4X0_RVT U2210 ( .A1(n1928), .A2(n1927), .A3(n1926), .A4(n1925), .Y(n1948) );
  NAND4X0_RVT U2211 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .Y(n1947) );
  NAND4X0_RVT U2212 ( .A1(n1937), .A2(n1936), .A3(n1935), .A4(n1934), .Y(n1938) );
  NOR4X1_RVT U2213 ( .A1(n1941), .A2(n1940), .A3(n1939), .A4(n1938), .Y(n1942)
         );
  NAND4X0_RVT U2214 ( .A1(n1945), .A2(n1944), .A3(n1943), .A4(n1942), .Y(n1946) );
  NOR4X1_RVT U2215 ( .A1(n1949), .A2(n1948), .A3(n1947), .A4(n1946), .Y(n1952)
         );
  AND4X1_RVT U2216 ( .A1(n1953), .A2(n1952), .A3(n1951), .A4(n1950), .Y(n1967)
         );
  AND4X1_RVT U2217 ( .A1(n1957), .A2(n1956), .A3(n1955), .A4(n1954), .Y(n1963)
         );
  AND4X1_RVT U2218 ( .A1(n1961), .A2(n1960), .A3(n1959), .A4(n1958), .Y(n1962)
         );
  AND4X1_RVT U2219 ( .A1(n1965), .A2(n1964), .A3(n1963), .A4(n1962), .Y(n1966)
         );
  AO221X1_RVT U2220 ( .A1(n1967), .A2(m4stg_sh_cnt[4]), .A3(n1967), .A4(n1966), 
        .A5(\m4stg_sh_cnt_5[0] ), .Y(n1968) );
  NAND4X0_RVT U2221 ( .A1(n1971), .A2(n1970), .A3(n1969), .A4(n1968), .Y(n1975) );
  AOI22X1_RVT U2222 ( .A1(n1973), .A2(n1975), .A3(m5stg_frac_32_0[0]), .A4(
        n1972), .Y(n1824) );
  NAND2X0_RVT U2223 ( .A1(n1974), .A2(m4stg_left_shift_step), .Y(n2032) );
  INVX1_RVT U2224 ( .A(n2032), .Y(n2017) );
  NAND2X0_RVT U2225 ( .A1(n2017), .A2(n1975), .Y(n1823) );
  OR2X1_RVT U2226 ( .A1(n2032), .A2(n1976), .Y(n1822) );
  OR2X1_RVT U2227 ( .A1(n2032), .A2(n1977), .Y(n1821) );
  OR2X1_RVT U2228 ( .A1(n2032), .A2(n1978), .Y(n1820) );
  NAND3X0_RVT U2229 ( .A1(n2017), .A2(n1980), .A3(n1979), .Y(n1819) );
  OR2X1_RVT U2230 ( .A1(n1981), .A2(n2032), .Y(n1818) );
  OR2X1_RVT U2231 ( .A1(n1982), .A2(n2032), .Y(n1817) );
  OR2X1_RVT U2232 ( .A1(n1983), .A2(n2032), .Y(n1816) );
  OR2X1_RVT U2233 ( .A1(n1984), .A2(n2032), .Y(n1815) );
  OR2X1_RVT U2234 ( .A1(n1985), .A2(n2032), .Y(n1814) );
  OR2X1_RVT U2235 ( .A1(n1986), .A2(n2032), .Y(n1813) );
  OR2X1_RVT U2236 ( .A1(n1987), .A2(n2032), .Y(n1812) );
  NAND3X0_RVT U2237 ( .A1(n2017), .A2(n1989), .A3(n1988), .Y(n1811) );
  OR2X1_RVT U2238 ( .A1(n1990), .A2(n2032), .Y(n1810) );
  OR2X1_RVT U2239 ( .A1(n2032), .A2(n1991), .Y(n1809) );
  OR2X1_RVT U2240 ( .A1(n1992), .A2(n2032), .Y(n1808) );
  OR2X1_RVT U2241 ( .A1(n1993), .A2(n2032), .Y(n1807) );
  OR2X1_RVT U2242 ( .A1(n1994), .A2(n2032), .Y(n1806) );
  OR2X1_RVT U2243 ( .A1(n2032), .A2(n1995), .Y(n1805) );
  OR2X1_RVT U2244 ( .A1(n1996), .A2(n2032), .Y(n1804) );
  NAND3X0_RVT U2245 ( .A1(n2017), .A2(n1998), .A3(n1997), .Y(n1803) );
  OR2X1_RVT U2246 ( .A1(n1999), .A2(n2032), .Y(n1802) );
  OR2X1_RVT U2247 ( .A1(n2000), .A2(n2032), .Y(n1801) );
  OR2X1_RVT U2248 ( .A1(n2001), .A2(n2032), .Y(n1800) );
  OR2X1_RVT U2249 ( .A1(n2002), .A2(n2032), .Y(n1799) );
  OR2X1_RVT U2250 ( .A1(n2003), .A2(n2032), .Y(n1798) );
  OR2X1_RVT U2251 ( .A1(n2004), .A2(n2032), .Y(n1797) );
  OR2X1_RVT U2252 ( .A1(n2005), .A2(n2032), .Y(n1796) );
  NAND3X0_RVT U2253 ( .A1(n2017), .A2(n2007), .A3(n2006), .Y(n1795) );
  OR2X1_RVT U2254 ( .A1(n2008), .A2(n2032), .Y(n1794) );
  OR2X1_RVT U2255 ( .A1(n2032), .A2(n2009), .Y(n1793) );
  OR2X1_RVT U2256 ( .A1(n2010), .A2(n2032), .Y(n1792) );
  OR2X1_RVT U2257 ( .A1(n2011), .A2(n2032), .Y(n1791) );
  OR2X1_RVT U2258 ( .A1(n2012), .A2(n2032), .Y(n1790) );
  OR2X1_RVT U2259 ( .A1(n2032), .A2(n2013), .Y(n1789) );
  OR2X1_RVT U2260 ( .A1(n2014), .A2(n2032), .Y(n1788) );
  NAND3X0_RVT U2261 ( .A1(n2017), .A2(n2016), .A3(n2015), .Y(n1787) );
  OR2X1_RVT U2262 ( .A1(n2018), .A2(n2032), .Y(n1786) );
  OR2X1_RVT U2263 ( .A1(n2019), .A2(n2032), .Y(n1785) );
  OR2X1_RVT U2264 ( .A1(n2020), .A2(n2032), .Y(n1784) );
  OR2X1_RVT U2265 ( .A1(n2021), .A2(n2032), .Y(n1783) );
  OR2X1_RVT U2266 ( .A1(n2022), .A2(n2032), .Y(n1782) );
  OR2X1_RVT U2267 ( .A1(n2023), .A2(n2032), .Y(n1781) );
  OR2X1_RVT U2268 ( .A1(n2024), .A2(n2032), .Y(n1780) );
  OR2X1_RVT U2269 ( .A1(n2032), .A2(n2025), .Y(n1779) );
  OR2X1_RVT U2270 ( .A1(n2026), .A2(n2032), .Y(n1778) );
  OR2X1_RVT U2271 ( .A1(n2032), .A2(n2027), .Y(n1777) );
  OR2X1_RVT U2272 ( .A1(n2028), .A2(n2032), .Y(n1776) );
  OR2X1_RVT U2273 ( .A1(n2029), .A2(n2032), .Y(n1775) );
  OR2X1_RVT U2274 ( .A1(n2030), .A2(n2032), .Y(n1774) );
  OR2X1_RVT U2275 ( .A1(n2032), .A2(n2031), .Y(n1773) );
  OR2X1_RVT U2276 ( .A1(n2033), .A2(n2032), .Y(n1772) );
  OR2X1_RVT U2277 ( .A1(n2032), .A2(n2034), .Y(n1771) );
  OR2X1_RVT U2278 ( .A1(n2035), .A2(n2032), .Y(n1770) );
  NAND2X0_RVT U2279 ( .A1(n2103), .A2(n2043), .Y(n1768) );
  NAND2X0_RVT U2280 ( .A1(n2102), .A2(n2043), .Y(n1767) );
  INVX1_RVT U2281 ( .A(n2036), .Y(n2100) );
  NAND2X0_RVT U2282 ( .A1(n2100), .A2(n2043), .Y(n1766) );
  INVX1_RVT U2283 ( .A(n2037), .Y(n2097) );
  NAND2X0_RVT U2284 ( .A1(n2097), .A2(n2043), .Y(n1764) );
  NAND2X0_RVT U2285 ( .A1(n2096), .A2(n2043), .Y(n1763) );
  INVX1_RVT U2286 ( .A(n2038), .Y(n2077) );
  NAND2X0_RVT U2287 ( .A1(n2077), .A2(n2043), .Y(n1746) );
  NAND2X0_RVT U2288 ( .A1(n2076), .A2(n2043), .Y(n1745) );
  INVX1_RVT U2289 ( .A(n2039), .Y(n2075) );
  NAND2X0_RVT U2290 ( .A1(n2075), .A2(n2043), .Y(n1744) );
  INVX1_RVT U2291 ( .A(n2040), .Y(n2074) );
  NAND2X0_RVT U2292 ( .A1(n2074), .A2(n2043), .Y(n1743) );
  NAND2X0_RVT U2293 ( .A1(n2073), .A2(n2043), .Y(n1742) );
  INVX1_RVT U2294 ( .A(n2041), .Y(n2072) );
  NAND2X0_RVT U2295 ( .A1(n2072), .A2(n2043), .Y(n1741) );
  INVX1_RVT U2296 ( .A(n2042), .Y(n2071) );
  NAND2X0_RVT U2297 ( .A1(n2071), .A2(n2043), .Y(n1740) );
  NAND2X0_RVT U2298 ( .A1(n2070), .A2(n2043), .Y(n1739) );
  NAND4X0_RVT U2299 ( .A1(n1593), .A2(n1539), .A3(m4stg_frac[105]), .A4(n2087), 
        .Y(n2044) );
  AND2X1_RVT U2300 ( .A1(m4stg_right_shift_step), .A2(n2044), .Y(n2086) );
  NAND2X0_RVT U2301 ( .A1(n2086), .A2(n2045), .Y(n1714) );
  NAND2X0_RVT U2302 ( .A1(n2086), .A2(n2046), .Y(n1713) );
  NAND2X0_RVT U2303 ( .A1(n2086), .A2(n2047), .Y(n1712) );
  NAND2X0_RVT U2304 ( .A1(n2086), .A2(n2048), .Y(n1711) );
  NAND2X0_RVT U2305 ( .A1(n2086), .A2(n2049), .Y(n1710) );
  NAND2X0_RVT U2306 ( .A1(n2086), .A2(n2050), .Y(n1709) );
  NAND2X0_RVT U2307 ( .A1(n2086), .A2(n2051), .Y(n1708) );
  NAND2X0_RVT U2308 ( .A1(n2086), .A2(n2052), .Y(n1707) );
  NAND2X0_RVT U2309 ( .A1(n2086), .A2(n2053), .Y(n1706) );
  NAND2X0_RVT U2310 ( .A1(n2086), .A2(n2054), .Y(n1705) );
  NAND2X0_RVT U2311 ( .A1(n2086), .A2(n2055), .Y(n1704) );
  NAND2X0_RVT U2312 ( .A1(n2086), .A2(n2056), .Y(n1703) );
  NAND2X0_RVT U2313 ( .A1(n2086), .A2(n2057), .Y(n1702) );
  NAND2X0_RVT U2314 ( .A1(n2086), .A2(n2058), .Y(n1701) );
  NAND2X0_RVT U2315 ( .A1(n2086), .A2(n2059), .Y(n1700) );
  NAND2X0_RVT U2316 ( .A1(n2086), .A2(n2060), .Y(n1699) );
  NAND2X0_RVT U2317 ( .A1(n2086), .A2(n2061), .Y(n1698) );
  NAND2X0_RVT U2318 ( .A1(n2086), .A2(n2062), .Y(n1697) );
  NAND2X0_RVT U2319 ( .A1(n2086), .A2(n2063), .Y(n1696) );
  NAND2X0_RVT U2320 ( .A1(n2086), .A2(n2064), .Y(n1695) );
  NAND2X0_RVT U2321 ( .A1(n2086), .A2(n2065), .Y(n1694) );
  NAND2X0_RVT U2322 ( .A1(n2086), .A2(n2066), .Y(n1693) );
  NAND2X0_RVT U2323 ( .A1(n2086), .A2(n2067), .Y(n1692) );
  NAND2X0_RVT U2324 ( .A1(n2086), .A2(n2068), .Y(n1691) );
  AND2X1_RVT U2325 ( .A1(n2086), .A2(n2069), .Y(n2099) );
  NAND2X0_RVT U2326 ( .A1(n2070), .A2(n2099), .Y(n1690) );
  NAND2X0_RVT U2327 ( .A1(n2071), .A2(n2099), .Y(n1689) );
  NAND2X0_RVT U2328 ( .A1(n2072), .A2(n2099), .Y(n1688) );
  NAND2X0_RVT U2329 ( .A1(n2073), .A2(n2099), .Y(n1687) );
  NAND2X0_RVT U2330 ( .A1(n2074), .A2(n2099), .Y(n1686) );
  NAND2X0_RVT U2331 ( .A1(n2075), .A2(n2099), .Y(n1685) );
  NAND2X0_RVT U2332 ( .A1(n2076), .A2(n2099), .Y(n1684) );
  NAND2X0_RVT U2333 ( .A1(n2077), .A2(n2099), .Y(n1683) );
  NAND2X0_RVT U2334 ( .A1(n2099), .A2(n2078), .Y(n1682) );
  NAND2X0_RVT U2335 ( .A1(n2099), .A2(n2079), .Y(n1681) );
  NAND2X0_RVT U2336 ( .A1(n2099), .A2(n2080), .Y(n1680) );
  NAND2X0_RVT U2337 ( .A1(n2099), .A2(n2081), .Y(n1679) );
  NAND2X0_RVT U2338 ( .A1(n2082), .A2(n2099), .Y(n1678) );
  NAND2X0_RVT U2339 ( .A1(n2083), .A2(n2099), .Y(n1677) );
  NAND2X0_RVT U2340 ( .A1(n2099), .A2(n2084), .Y(n1676) );
  NAND2X0_RVT U2341 ( .A1(n2085), .A2(n2099), .Y(n1675) );
  AND2X1_RVT U2342 ( .A1(n2087), .A2(n2086), .Y(n2104) );
  NAND2X0_RVT U2343 ( .A1(n2104), .A2(n2088), .Y(n1674) );
  NAND2X0_RVT U2344 ( .A1(n2104), .A2(n2089), .Y(n1673) );
  NAND2X0_RVT U2345 ( .A1(n2104), .A2(n2090), .Y(n1672) );
  NAND2X0_RVT U2346 ( .A1(n2104), .A2(n2091), .Y(n1671) );
  NAND2X0_RVT U2347 ( .A1(n2104), .A2(n2092), .Y(n1670) );
  NAND2X0_RVT U2348 ( .A1(n2104), .A2(n2093), .Y(n1669) );
  NAND2X0_RVT U2349 ( .A1(n2104), .A2(n2094), .Y(n1668) );
  NAND2X0_RVT U2350 ( .A1(n2104), .A2(n2095), .Y(n1667) );
  NAND3X0_RVT U2351 ( .A1(n2101), .A2(n2096), .A3(n2099), .Y(n1666) );
  NAND3X0_RVT U2352 ( .A1(n2101), .A2(n2097), .A3(n2099), .Y(n1665) );
  NAND3X0_RVT U2353 ( .A1(n2101), .A2(n2099), .A3(n2098), .Y(n1664) );
  NAND3X0_RVT U2354 ( .A1(n2101), .A2(n2100), .A3(n2099), .Y(n1663) );
  NAND3X0_RVT U2355 ( .A1(n1539), .A2(n2104), .A3(n2102), .Y(n1662) );
  NAND3X0_RVT U2356 ( .A1(n1539), .A2(n2104), .A3(n2103), .Y(n1661) );
  AO22X1_RVT U2357 ( .A1(mul_frac_in1[51]), .A2(m2stg_frac1_dbl_dnrm), .A3(
        m2stg_frac1_sng_dnrm), .A4(mul_frac_in1[54]), .Y(n2105) );
  NOR4X1_RVT U2358 ( .A1(m2stg_frac1_dbl_norm), .A2(m2stg_frac1_sng_norm), 
        .A3(m2stg_frac1_inf), .A4(n2105), .Y(m2stg_frac1_array_in[52]) );
  AO22X1_RVT U2359 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[50]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[49]), .Y(n2107) );
  AO22X1_RVT U2360 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[52]), .A3(
        mul_frac_in1[53]), .A4(m2stg_frac1_sng_norm), .Y(n2106) );
  NOR2X0_RVT U2361 ( .A1(n2107), .A2(n2106), .Y(m2stg_frac1_array_in[50]) );
  AO22X1_RVT U2362 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[49]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[48]), .Y(n2109) );
  AO22X1_RVT U2363 ( .A1(mul_frac_in1[51]), .A2(m2stg_frac1_sng_dnrm), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[52]), .Y(n2108) );
  NOR2X0_RVT U2364 ( .A1(n2109), .A2(n2108), .Y(m2stg_frac1_array_in[49]) );
  AO22X1_RVT U2365 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[48]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[47]), .Y(n2111) );
  AO22X1_RVT U2366 ( .A1(mul_frac_in1[51]), .A2(m2stg_frac1_sng_norm), .A3(
        mul_frac_in1[50]), .A4(m2stg_frac1_sng_dnrm), .Y(n2110) );
  NOR2X0_RVT U2367 ( .A1(n2111), .A2(n2110), .Y(m2stg_frac1_array_in[48]) );
  AO22X1_RVT U2368 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[47]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[46]), .Y(n2113) );
  AO22X1_RVT U2369 ( .A1(mul_frac_in1[50]), .A2(m2stg_frac1_sng_norm), .A3(
        m2stg_frac1_sng_dnrm), .A4(mul_frac_in1[49]), .Y(n2112) );
  NOR2X0_RVT U2370 ( .A1(n2113), .A2(n2112), .Y(m2stg_frac1_array_in[47]) );
  AO22X1_RVT U2371 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[46]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[45]), .Y(n2115) );
  AO22X1_RVT U2372 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[48]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[49]), .Y(n2114) );
  NOR2X0_RVT U2373 ( .A1(n2115), .A2(n2114), .Y(m2stg_frac1_array_in[46]) );
  AO22X1_RVT U2374 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[45]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[44]), .Y(n2117) );
  AO22X1_RVT U2375 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[47]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[48]), .Y(n2116) );
  NOR2X0_RVT U2376 ( .A1(n2117), .A2(n2116), .Y(m2stg_frac1_array_in[45]) );
  AO22X1_RVT U2377 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[44]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[43]), .Y(n2119) );
  AO22X1_RVT U2378 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[46]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[47]), .Y(n2118) );
  NOR2X0_RVT U2379 ( .A1(n2119), .A2(n2118), .Y(m2stg_frac1_array_in[44]) );
  AO22X1_RVT U2380 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[43]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[42]), .Y(n2121) );
  AO22X1_RVT U2381 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[45]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[46]), .Y(n2120) );
  NOR2X0_RVT U2382 ( .A1(n2121), .A2(n2120), .Y(m2stg_frac1_array_in[43]) );
  AO22X1_RVT U2383 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[42]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[41]), .Y(n2123) );
  AO22X1_RVT U2384 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[44]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[45]), .Y(n2122) );
  NOR2X0_RVT U2385 ( .A1(n2123), .A2(n2122), .Y(m2stg_frac1_array_in[42]) );
  AO22X1_RVT U2386 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[41]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[40]), .Y(n2125) );
  AO22X1_RVT U2387 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[43]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[44]), .Y(n2124) );
  NOR2X0_RVT U2388 ( .A1(n2125), .A2(n2124), .Y(m2stg_frac1_array_in[41]) );
  AO22X1_RVT U2389 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[40]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[39]), .Y(n2127) );
  AO22X1_RVT U2390 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[42]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[43]), .Y(n2126) );
  NOR2X0_RVT U2391 ( .A1(n2127), .A2(n2126), .Y(m2stg_frac1_array_in[40]) );
  AO22X1_RVT U2392 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[39]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[38]), .Y(n2129) );
  AO22X1_RVT U2393 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[41]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[42]), .Y(n2128) );
  NOR2X0_RVT U2394 ( .A1(n2129), .A2(n2128), .Y(m2stg_frac1_array_in[39]) );
  AO22X1_RVT U2395 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[38]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[37]), .Y(n2131) );
  AO22X1_RVT U2396 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[40]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[41]), .Y(n2130) );
  NOR2X0_RVT U2397 ( .A1(n2131), .A2(n2130), .Y(m2stg_frac1_array_in[38]) );
  AO22X1_RVT U2398 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[37]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[36]), .Y(n2133) );
  AO22X1_RVT U2399 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[39]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[40]), .Y(n2132) );
  NOR2X0_RVT U2400 ( .A1(n2133), .A2(n2132), .Y(m2stg_frac1_array_in[37]) );
  AO22X1_RVT U2401 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[36]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[35]), .Y(n2135) );
  AO22X1_RVT U2402 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[38]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[39]), .Y(n2134) );
  NOR2X0_RVT U2403 ( .A1(n2135), .A2(n2134), .Y(m2stg_frac1_array_in[36]) );
  AO22X1_RVT U2404 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[35]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[34]), .Y(n2137) );
  AO22X1_RVT U2405 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[37]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[38]), .Y(n2136) );
  NOR2X0_RVT U2406 ( .A1(n2137), .A2(n2136), .Y(m2stg_frac1_array_in[35]) );
  AO22X1_RVT U2407 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[34]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[33]), .Y(n2139) );
  AO22X1_RVT U2408 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[36]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[37]), .Y(n2138) );
  NOR2X0_RVT U2409 ( .A1(n2139), .A2(n2138), .Y(m2stg_frac1_array_in[34]) );
  AO22X1_RVT U2410 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[33]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[32]), .Y(n2141) );
  AO22X1_RVT U2411 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[35]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[36]), .Y(n2140) );
  NOR2X0_RVT U2412 ( .A1(n2141), .A2(n2140), .Y(m2stg_frac1_array_in[33]) );
  AO22X1_RVT U2413 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[32]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[31]), .Y(n2143) );
  AO22X1_RVT U2414 ( .A1(m2stg_frac1_sng_dnrm), .A2(mul_frac_in1[34]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[35]), .Y(n2142) );
  NOR2X0_RVT U2415 ( .A1(n2143), .A2(n2142), .Y(m2stg_frac1_array_in[32]) );
  AO22X1_RVT U2416 ( .A1(m2stg_frac1_dbl_dnrm), .A2(mul_frac_in1[30]), .A3(
        m2stg_frac1_sng_dnrm), .A4(mul_frac_in1[33]), .Y(n2145) );
  AO22X1_RVT U2417 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[31]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[34]), .Y(n2144) );
  NOR2X0_RVT U2418 ( .A1(n2145), .A2(n2144), .Y(m2stg_frac1_array_in[31]) );
  AO22X1_RVT U2419 ( .A1(m2stg_frac1_dbl_dnrm), .A2(mul_frac_in1[29]), .A3(
        m2stg_frac1_sng_dnrm), .A4(mul_frac_in1[32]), .Y(n2147) );
  AO22X1_RVT U2420 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[30]), .A3(
        m2stg_frac1_sng_norm), .A4(mul_frac_in1[33]), .Y(n2146) );
  NOR2X0_RVT U2421 ( .A1(n2147), .A2(n2146), .Y(m2stg_frac1_array_in[30]) );
  AOI222X1_RVT U2422 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[29]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[28]), .A5(m2stg_frac1_sng_norm), .A6(mul_frac_in1[32]), .Y(m2stg_frac1_array_in[29]) );
  AOI22X1_RVT U2423 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[28]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[27]), .Y(
        m2stg_frac1_array_in[28]) );
  AOI22X1_RVT U2424 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[27]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[26]), .Y(
        m2stg_frac1_array_in[27]) );
  AOI22X1_RVT U2425 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[26]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[25]), .Y(
        m2stg_frac1_array_in[26]) );
  AOI22X1_RVT U2426 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[25]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[24]), .Y(
        m2stg_frac1_array_in[25]) );
  AOI22X1_RVT U2427 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[24]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[23]), .Y(
        m2stg_frac1_array_in[24]) );
  AOI22X1_RVT U2428 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[23]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[22]), .Y(
        m2stg_frac1_array_in[23]) );
  AOI22X1_RVT U2429 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[22]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[21]), .Y(
        m2stg_frac1_array_in[22]) );
  AOI22X1_RVT U2430 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[21]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[20]), .Y(
        m2stg_frac1_array_in[21]) );
  AOI22X1_RVT U2431 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[20]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[19]), .Y(
        m2stg_frac1_array_in[20]) );
  AOI22X1_RVT U2432 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[19]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[18]), .Y(
        m2stg_frac1_array_in[19]) );
  AOI22X1_RVT U2433 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[18]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[17]), .Y(
        m2stg_frac1_array_in[18]) );
  AOI22X1_RVT U2434 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[17]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[16]), .Y(
        m2stg_frac1_array_in[17]) );
  AOI22X1_RVT U2435 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[16]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[15]), .Y(
        m2stg_frac1_array_in[16]) );
  AOI22X1_RVT U2436 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[15]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[14]), .Y(
        m2stg_frac1_array_in[15]) );
  AOI22X1_RVT U2437 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[14]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[13]), .Y(
        m2stg_frac1_array_in[14]) );
  AOI22X1_RVT U2438 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[13]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[12]), .Y(
        m2stg_frac1_array_in[13]) );
  AOI22X1_RVT U2439 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[12]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[11]), .Y(
        m2stg_frac1_array_in[12]) );
  AOI22X1_RVT U2440 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[11]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[10]), .Y(
        m2stg_frac1_array_in[11]) );
  AOI22X1_RVT U2441 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[10]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[9]), .Y(
        m2stg_frac1_array_in[10]) );
  AOI22X1_RVT U2442 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[9]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[8]), .Y(
        m2stg_frac1_array_in[9]) );
  AOI22X1_RVT U2443 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[8]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[7]), .Y(
        m2stg_frac1_array_in[8]) );
  AOI22X1_RVT U2444 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[7]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[6]), .Y(
        m2stg_frac1_array_in[7]) );
  AOI22X1_RVT U2445 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[6]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[5]), .Y(
        m2stg_frac1_array_in[6]) );
  AOI22X1_RVT U2446 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[5]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[4]), .Y(
        m2stg_frac1_array_in[5]) );
  AOI22X1_RVT U2447 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[4]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[3]), .Y(
        m2stg_frac1_array_in[4]) );
  AOI22X1_RVT U2448 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[3]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[2]), .Y(
        m2stg_frac1_array_in[3]) );
  AOI22X1_RVT U2449 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[2]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[1]), .Y(
        m2stg_frac1_array_in[2]) );
  AOI22X1_RVT U2450 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[1]), .A3(
        m2stg_frac1_dbl_dnrm), .A4(mul_frac_in1[0]), .Y(
        m2stg_frac1_array_in[1]) );
  NAND2X0_RVT U2451 ( .A1(m2stg_frac1_dbl_norm), .A2(mul_frac_in1[0]), .Y(
        m2stg_frac1_array_in[0]) );
endmodule


module mul_bodec_0 ( x, b, b0, b1, b2, b3, b4, b5, b6, b7 );
  input [15:0] b;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  input x;
  wire   b_12, b_10, b_8, b_6, b_4, b_2, b_0, \b[1] , \b[3] , \b[5] , \b[7] ,
         \b[9] , \b[11] , \b[13] , \b[15] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15;
  assign b_12 = b[12];
  assign b_10 = b[10];
  assign b_8 = b[8];
  assign b_6 = b[6];
  assign b_4 = b[4];
  assign b_2 = b[2];
  assign b_0 = b[0];
  assign b0[2] = \b[1] ;
  assign \b[1]  = b[1];
  assign b1[2] = \b[3] ;
  assign \b[3]  = b[3];
  assign b2[2] = \b[5] ;
  assign \b[5]  = b[5];
  assign b3[2] = \b[7] ;
  assign \b[7]  = b[7];
  assign b4[2] = \b[9] ;
  assign \b[9]  = b[9];
  assign b5[2] = \b[11] ;
  assign \b[11]  = b[11];
  assign b6[2] = \b[13] ;
  assign \b[13]  = b[13];
  assign b7[2] = \b[15] ;
  assign \b[15]  = b[15];

  INVX0_RVT U1 ( .A(\b[15] ), .Y(n15) );
  INVX1_RVT U2 ( .A(\b[1] ), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(b_0), .A2(n2), .Y(b0[0]) );
  OR2X1_RVT U4 ( .A1(\b[1] ), .A2(b_0), .Y(b0[1]) );
  INVX1_RVT U5 ( .A(\b[3] ), .Y(n4) );
  INVX1_RVT U6 ( .A(b_2), .Y(n1) );
  OA222X1_RVT U7 ( .A1(\b[1] ), .A2(\b[3] ), .A3(n2), .A4(b_2), .A5(n4), .A6(
        n1), .Y(b1[0]) );
  INVX1_RVT U8 ( .A(\b[5] ), .Y(n6) );
  INVX1_RVT U9 ( .A(b_4), .Y(n3) );
  OA222X1_RVT U10 ( .A1(\b[3] ), .A2(\b[5] ), .A3(n4), .A4(b_4), .A5(n6), .A6(
        n3), .Y(b2[0]) );
  INVX1_RVT U11 ( .A(\b[7] ), .Y(n8) );
  INVX1_RVT U12 ( .A(b_6), .Y(n5) );
  OA222X1_RVT U13 ( .A1(\b[5] ), .A2(\b[7] ), .A3(n6), .A4(b_6), .A5(n8), .A6(
        n5), .Y(b3[0]) );
  INVX1_RVT U14 ( .A(\b[9] ), .Y(n10) );
  INVX1_RVT U15 ( .A(b_8), .Y(n7) );
  OA222X1_RVT U16 ( .A1(\b[7] ), .A2(\b[9] ), .A3(n8), .A4(b_8), .A5(n10), 
        .A6(n7), .Y(b4[0]) );
  INVX1_RVT U17 ( .A(\b[11] ), .Y(n12) );
  INVX1_RVT U18 ( .A(b_10), .Y(n9) );
  OA222X1_RVT U19 ( .A1(\b[9] ), .A2(\b[11] ), .A3(n10), .A4(b_10), .A5(n12), 
        .A6(n9), .Y(b5[0]) );
  INVX1_RVT U20 ( .A(\b[13] ), .Y(n14) );
  INVX1_RVT U21 ( .A(b_12), .Y(n11) );
  OA222X1_RVT U22 ( .A1(\b[11] ), .A2(\b[13] ), .A3(n12), .A4(b_12), .A5(n14), 
        .A6(n11), .Y(b6[0]) );
  INVX1_RVT U23 ( .A(b[14]), .Y(n13) );
  OA222X1_RVT U24 ( .A1(\b[13] ), .A2(\b[15] ), .A3(n14), .A4(b[14]), .A5(n15), 
        .A6(n13), .Y(b7[0]) );
  AO222X1_RVT U25 ( .A1(\b[1] ), .A2(n4), .A3(n2), .A4(b_2), .A5(\b[3] ), .A6(
        n1), .Y(b1[1]) );
  AO222X1_RVT U26 ( .A1(\b[3] ), .A2(n6), .A3(n4), .A4(b_4), .A5(\b[5] ), .A6(
        n3), .Y(b2[1]) );
  AO222X1_RVT U27 ( .A1(\b[5] ), .A2(n8), .A3(n6), .A4(b_6), .A5(\b[7] ), .A6(
        n5), .Y(b3[1]) );
  AO222X1_RVT U28 ( .A1(\b[7] ), .A2(n10), .A3(n8), .A4(b_8), .A5(\b[9] ), 
        .A6(n7), .Y(b4[1]) );
  AO222X1_RVT U29 ( .A1(\b[9] ), .A2(n12), .A3(n10), .A4(b_10), .A5(\b[11] ), 
        .A6(n9), .Y(b5[1]) );
  AO222X1_RVT U30 ( .A1(\b[11] ), .A2(n14), .A3(n12), .A4(b_12), .A5(\b[13] ), 
        .A6(n11), .Y(b6[1]) );
  AO222X1_RVT U31 ( .A1(\b[13] ), .A2(n15), .A3(n14), .A4(b[14]), .A5(\b[15] ), 
        .A6(n13), .Y(b7[1]) );
endmodule


module dp_mux2es_SIZE3_0 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module clken_buf_1 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module clken_buf_2 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module dp_mux2es_SIZE3_1 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AND2X1_RVT U2 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
  AND2X1_RVT U3 ( .A1(in0[1]), .A2(n1), .Y(dout[1]) );
  AND2X1_RVT U4 ( .A1(in0[0]), .A2(n1), .Y(dout[0]) );
endmodule


module dp_mux2es_SIZE3_2 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AND2X1_RVT U2 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
  AND2X1_RVT U3 ( .A1(in0[1]), .A2(n1), .Y(dout[1]) );
  AND2X1_RVT U4 ( .A1(in0[0]), .A2(n1), .Y(dout[0]) );
endmodule


module dp_mux2es_SIZE3_3 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AND2X1_RVT U2 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
  AND2X1_RVT U3 ( .A1(in0[1]), .A2(n1), .Y(dout[1]) );
  AND2X1_RVT U4 ( .A1(in0[0]), .A2(n1), .Y(dout[0]) );
endmodule


module dp_mux2es_SIZE3_4 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AND2X1_RVT U2 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
  AND2X1_RVT U3 ( .A1(in0[1]), .A2(n1), .Y(dout[1]) );
  AND2X1_RVT U4 ( .A1(in0[0]), .A2(n1), .Y(dout[0]) );
endmodule


module dp_mux2es_SIZE3_5 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AND2X1_RVT U2 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
  AND2X1_RVT U3 ( .A1(in0[1]), .A2(n1), .Y(dout[1]) );
  AND2X1_RVT U4 ( .A1(in0[0]), .A2(n1), .Y(dout[0]) );
endmodule


module dp_mux2es_SIZE3_6 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AND2X1_RVT U4 ( .A1(in0[2]), .A2(n1), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_7 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_8 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_9 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_10 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_11 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_12 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_13 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_14 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module dp_mux2es_SIZE3_15 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   n1;

  INVX0_RVT U1 ( .A(sel), .Y(n1) );
  AO22X1_RVT U2 ( .A1(sel), .A2(in1[0]), .A3(n1), .A4(in0[0]), .Y(dout[0]) );
  AO22X1_RVT U3 ( .A1(sel), .A2(in1[1]), .A3(n1), .A4(in0[1]), .Y(dout[1]) );
  AO22X1_RVT U4 ( .A1(sel), .A2(in1[2]), .A3(n1), .A4(in0[2]), .Y(dout[2]) );
endmodule


module mul_bodec_1 ( x, b, b0, b1, b2, b3, b4, b5, b6, b7 );
  input [15:0] b;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  input x;
  wire   b_4, b_2, b_0, \b[1] , \b[3] , n1, n2, n3, n4, n5;
  assign b_4 = b[4];
  assign b_2 = b[2];
  assign b_0 = b[0];
  assign b0[2] = \b[1] ;
  assign \b[1]  = b[1];
  assign b1[2] = \b[3] ;
  assign \b[3]  = b[3];

  INVX0_RVT U1 ( .A(x), .Y(n3) );
  INVX0_RVT U2 ( .A(\b[3] ), .Y(n1) );
  AND2X1_RVT U3 ( .A1(\b[3] ), .A2(b_4), .Y(b2[0]) );
  OR2X1_RVT U4 ( .A1(\b[3] ), .A2(b_4), .Y(b2[1]) );
  INVX1_RVT U5 ( .A(b_0), .Y(n4) );
  INVX1_RVT U6 ( .A(\b[1] ), .Y(n5) );
  OA222X1_RVT U7 ( .A1(b_0), .A2(\b[1] ), .A3(n4), .A4(x), .A5(n5), .A6(n3), 
        .Y(b0[0]) );
  INVX1_RVT U8 ( .A(b_2), .Y(n2) );
  OA222X1_RVT U9 ( .A1(\b[1] ), .A2(\b[3] ), .A3(n5), .A4(b_2), .A5(n1), .A6(
        n2), .Y(b1[0]) );
  AO222X1_RVT U10 ( .A1(\b[1] ), .A2(n2), .A3(n5), .A4(\b[3] ), .A5(b_2), .A6(
        n1), .Y(b1[1]) );
  AO222X1_RVT U11 ( .A1(b_0), .A2(n5), .A3(n4), .A4(x), .A5(\b[1] ), .A6(n3), 
        .Y(b0[1]) );
endmodule


module mul_bodec_2 ( x, b, b0, b1, b2, b3, b4, b5, b6, b7 );
  input [15:0] b;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  input x;
  wire   b_12, b_10, b_8, b_6, b_4, b_2, b_0, \b[1] , \b[3] , \b[5] , \b[7] ,
         \b[9] , \b[11] , \b[13] , \b[15] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17;
  assign b_12 = b[12];
  assign b_10 = b[10];
  assign b_8 = b[8];
  assign b_6 = b[6];
  assign b_4 = b[4];
  assign b_2 = b[2];
  assign b_0 = b[0];
  assign b0[2] = \b[1] ;
  assign \b[1]  = b[1];
  assign b1[2] = \b[3] ;
  assign \b[3]  = b[3];
  assign b2[2] = \b[5] ;
  assign \b[5]  = b[5];
  assign b3[2] = \b[7] ;
  assign \b[7]  = b[7];
  assign b4[2] = \b[9] ;
  assign \b[9]  = b[9];
  assign b5[2] = \b[11] ;
  assign \b[11]  = b[11];
  assign b6[2] = \b[13] ;
  assign \b[13]  = b[13];
  assign b7[2] = \b[15] ;
  assign \b[15]  = b[15];

  INVX0_RVT U1 ( .A(\b[15] ), .Y(n14) );
  INVX1_RVT U2 ( .A(b_0), .Y(n16) );
  INVX1_RVT U3 ( .A(\b[1] ), .Y(n17) );
  INVX1_RVT U4 ( .A(x), .Y(n15) );
  OA222X1_RVT U5 ( .A1(b_0), .A2(\b[1] ), .A3(n16), .A4(x), .A5(n17), .A6(n15), 
        .Y(b0[0]) );
  INVX1_RVT U6 ( .A(\b[3] ), .Y(n3) );
  INVX1_RVT U7 ( .A(b_2), .Y(n1) );
  OA222X1_RVT U8 ( .A1(\b[1] ), .A2(\b[3] ), .A3(n17), .A4(b_2), .A5(n3), .A6(
        n1), .Y(b1[0]) );
  INVX1_RVT U9 ( .A(\b[5] ), .Y(n5) );
  INVX1_RVT U10 ( .A(b_4), .Y(n2) );
  OA222X1_RVT U11 ( .A1(\b[3] ), .A2(\b[5] ), .A3(n3), .A4(b_4), .A5(n5), .A6(
        n2), .Y(b2[0]) );
  INVX1_RVT U12 ( .A(\b[7] ), .Y(n7) );
  INVX1_RVT U13 ( .A(b_6), .Y(n4) );
  OA222X1_RVT U14 ( .A1(\b[5] ), .A2(\b[7] ), .A3(n5), .A4(b_6), .A5(n7), .A6(
        n4), .Y(b3[0]) );
  INVX1_RVT U15 ( .A(\b[9] ), .Y(n9) );
  INVX1_RVT U16 ( .A(b_8), .Y(n6) );
  OA222X1_RVT U17 ( .A1(\b[7] ), .A2(\b[9] ), .A3(n7), .A4(b_8), .A5(n9), .A6(
        n6), .Y(b4[0]) );
  INVX1_RVT U18 ( .A(\b[11] ), .Y(n11) );
  INVX1_RVT U19 ( .A(b_10), .Y(n8) );
  OA222X1_RVT U20 ( .A1(\b[9] ), .A2(\b[11] ), .A3(n9), .A4(b_10), .A5(n11), 
        .A6(n8), .Y(b5[0]) );
  INVX1_RVT U21 ( .A(\b[13] ), .Y(n13) );
  INVX1_RVT U22 ( .A(b_12), .Y(n10) );
  OA222X1_RVT U23 ( .A1(\b[11] ), .A2(\b[13] ), .A3(n11), .A4(b_12), .A5(n13), 
        .A6(n10), .Y(b6[0]) );
  INVX1_RVT U24 ( .A(b[14]), .Y(n12) );
  OA222X1_RVT U25 ( .A1(\b[13] ), .A2(\b[15] ), .A3(n13), .A4(b[14]), .A5(n14), 
        .A6(n12), .Y(b7[0]) );
  AO222X1_RVT U26 ( .A1(\b[1] ), .A2(n3), .A3(n17), .A4(b_2), .A5(\b[3] ), 
        .A6(n1), .Y(b1[1]) );
  AO222X1_RVT U27 ( .A1(\b[3] ), .A2(n5), .A3(n3), .A4(b_4), .A5(\b[5] ), .A6(
        n2), .Y(b2[1]) );
  AO222X1_RVT U28 ( .A1(\b[5] ), .A2(n7), .A3(n5), .A4(b_6), .A5(\b[7] ), .A6(
        n4), .Y(b3[1]) );
  AO222X1_RVT U29 ( .A1(\b[7] ), .A2(n9), .A3(n7), .A4(b_8), .A5(\b[9] ), .A6(
        n6), .Y(b4[1]) );
  AO222X1_RVT U30 ( .A1(\b[9] ), .A2(n11), .A3(n9), .A4(b_10), .A5(\b[11] ), 
        .A6(n8), .Y(b5[1]) );
  AO222X1_RVT U31 ( .A1(\b[11] ), .A2(n13), .A3(n11), .A4(b_12), .A5(\b[13] ), 
        .A6(n10), .Y(b6[1]) );
  AO222X1_RVT U32 ( .A1(\b[13] ), .A2(n14), .A3(n13), .A4(b[14]), .A5(\b[15] ), 
        .A6(n12), .Y(b7[1]) );
  AO222X1_RVT U33 ( .A1(b_0), .A2(n17), .A3(n16), .A4(x), .A5(\b[1] ), .A6(n15), .Y(b0[1]) );
endmodule


module mul_bodec_3 ( x, b, b0, b1, b2, b3, b4, b5, b6, b7 );
  input [15:0] b;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  input x;
  wire   b_12, b_10, b_8, b_6, b_4, b_2, b_0, \b[1] , \b[3] , \b[5] , \b[7] ,
         \b[9] , \b[11] , \b[13] , \b[15] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17;
  assign b_12 = b[12];
  assign b_10 = b[10];
  assign b_8 = b[8];
  assign b_6 = b[6];
  assign b_4 = b[4];
  assign b_2 = b[2];
  assign b_0 = b[0];
  assign b0[2] = \b[1] ;
  assign \b[1]  = b[1];
  assign b1[2] = \b[3] ;
  assign \b[3]  = b[3];
  assign b2[2] = \b[5] ;
  assign \b[5]  = b[5];
  assign b3[2] = \b[7] ;
  assign \b[7]  = b[7];
  assign b4[2] = \b[9] ;
  assign \b[9]  = b[9];
  assign b5[2] = \b[11] ;
  assign \b[11]  = b[11];
  assign b6[2] = \b[13] ;
  assign \b[13]  = b[13];
  assign b7[2] = \b[15] ;
  assign \b[15]  = b[15];

  INVX0_RVT U1 ( .A(x), .Y(n15) );
  INVX0_RVT U2 ( .A(b_0), .Y(n16) );
  INVX0_RVT U3 ( .A(\b[15] ), .Y(n14) );
  INVX1_RVT U4 ( .A(\b[1] ), .Y(n17) );
  OA222X1_RVT U5 ( .A1(b_0), .A2(\b[1] ), .A3(n16), .A4(x), .A5(n17), .A6(n15), 
        .Y(b0[0]) );
  INVX1_RVT U6 ( .A(\b[3] ), .Y(n3) );
  INVX1_RVT U7 ( .A(b_2), .Y(n1) );
  OA222X1_RVT U8 ( .A1(\b[1] ), .A2(\b[3] ), .A3(n17), .A4(b_2), .A5(n3), .A6(
        n1), .Y(b1[0]) );
  INVX1_RVT U9 ( .A(\b[5] ), .Y(n5) );
  INVX1_RVT U10 ( .A(b_4), .Y(n2) );
  OA222X1_RVT U11 ( .A1(\b[3] ), .A2(\b[5] ), .A3(n3), .A4(b_4), .A5(n5), .A6(
        n2), .Y(b2[0]) );
  INVX1_RVT U12 ( .A(\b[7] ), .Y(n7) );
  INVX1_RVT U13 ( .A(b_6), .Y(n4) );
  OA222X1_RVT U14 ( .A1(\b[5] ), .A2(\b[7] ), .A3(n5), .A4(b_6), .A5(n7), .A6(
        n4), .Y(b3[0]) );
  INVX1_RVT U15 ( .A(\b[9] ), .Y(n9) );
  INVX1_RVT U16 ( .A(b_8), .Y(n6) );
  OA222X1_RVT U17 ( .A1(\b[7] ), .A2(\b[9] ), .A3(n7), .A4(b_8), .A5(n9), .A6(
        n6), .Y(b4[0]) );
  INVX1_RVT U18 ( .A(\b[11] ), .Y(n11) );
  INVX1_RVT U19 ( .A(b_10), .Y(n8) );
  OA222X1_RVT U20 ( .A1(\b[9] ), .A2(\b[11] ), .A3(n9), .A4(b_10), .A5(n11), 
        .A6(n8), .Y(b5[0]) );
  INVX1_RVT U21 ( .A(\b[13] ), .Y(n13) );
  INVX1_RVT U22 ( .A(b_12), .Y(n10) );
  OA222X1_RVT U23 ( .A1(\b[11] ), .A2(\b[13] ), .A3(n11), .A4(b_12), .A5(n13), 
        .A6(n10), .Y(b6[0]) );
  INVX1_RVT U24 ( .A(b[14]), .Y(n12) );
  OA222X1_RVT U25 ( .A1(\b[13] ), .A2(\b[15] ), .A3(n13), .A4(b[14]), .A5(n14), 
        .A6(n12), .Y(b7[0]) );
  AO222X1_RVT U26 ( .A1(\b[1] ), .A2(n3), .A3(n17), .A4(b_2), .A5(\b[3] ), 
        .A6(n1), .Y(b1[1]) );
  AO222X1_RVT U27 ( .A1(\b[3] ), .A2(n5), .A3(n3), .A4(b_4), .A5(\b[5] ), .A6(
        n2), .Y(b2[1]) );
  AO222X1_RVT U28 ( .A1(\b[5] ), .A2(n7), .A3(n5), .A4(b_6), .A5(\b[7] ), .A6(
        n4), .Y(b3[1]) );
  AO222X1_RVT U29 ( .A1(\b[7] ), .A2(n9), .A3(n7), .A4(b_8), .A5(\b[9] ), .A6(
        n6), .Y(b4[1]) );
  AO222X1_RVT U30 ( .A1(\b[9] ), .A2(n11), .A3(n9), .A4(b_10), .A5(\b[11] ), 
        .A6(n8), .Y(b5[1]) );
  AO222X1_RVT U31 ( .A1(\b[11] ), .A2(n13), .A3(n11), .A4(b_12), .A5(\b[13] ), 
        .A6(n10), .Y(b6[1]) );
  AO222X1_RVT U32 ( .A1(\b[13] ), .A2(n14), .A3(n13), .A4(b[14]), .A5(\b[15] ), 
        .A6(n12), .Y(b7[1]) );
  AO222X1_RVT U33 ( .A1(b_0), .A2(n17), .A3(n16), .A4(x), .A5(\b[1] ), .A6(n15), .Y(b0[1]) );
endmodule


module dff_SIZE1_2 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE32_1 ( din, clk, q, se, si, so );
  input [31:0] din;
  output [31:0] q;
  input [31:0] si;
  output [31:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, n1;
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
endmodule


module dff_SIZE3_16 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_15 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_14 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_13 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_12 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_11 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_10 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_9 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_8 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_7 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_6 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_5 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_4 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_3 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_2 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE3_1 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module mul_booth ( head, b_in, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, 
        b11, b12, b13, b14, b15, b16, clk, se, si, so, mul_step, tm_l );
  input [63:0] b_in;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  output [2:0] b8;
  output [2:0] b9;
  output [2:0] b10;
  output [2:0] b11;
  output [2:0] b12;
  output [2:0] b13;
  output [2:0] b14;
  output [2:0] b15;
  input head, clk, se, si, mul_step, tm_l;
  output b16, so;
  wire   clk_enb0, clk_enb1, n3, n1, n2, net210894, net210895, net210896,
         net210897, net210898, net210899, net210900, net210901, net210902,
         net210903, net210904, net210905, net210906, net210907, net210908,
         net210909, net210910, net210911, net210912, net210913, net210914,
         net210915, net210916, net210917, net210918, net210919, net210920,
         net210921, net210922, net210923, net210924, net210925, net210926,
         net210927, net210928, net210929, net210930, net210931;
  wire   [2:0] b0_in0;
  wire   [2:0] b1_in0;
  wire   [2:0] b2_in0;
  wire   [2:0] b3_in0;
  wire   [2:0] b4_in0;
  wire   [2:0] b5_in0;
  wire   [2:0] b6_in0;
  wire   [2:0] b7_in0;
  wire   [2:0] b8_in0;
  wire   [2:0] b9_in0;
  wire   [2:0] b10_in0;
  wire   [2:0] b11_in0;
  wire   [2:0] b12_in0;
  wire   [2:0] b13_in0;
  wire   [2:0] b14_in0;
  wire   [2:0] b15_in0;
  wire   [63:31] b;
  wire   [2:0] b0_in1;
  wire   [2:0] b1_in1;
  wire   [2:0] b2_in1;
  wire   [2:0] b3_in1;
  wire   [2:0] b4_in1;
  wire   [2:0] b5_in1;
  wire   [2:0] b6_in1;
  wire   [2:0] b7_in1;
  wire   [2:0] b8_in1;
  wire   [2:0] b9_in1;
  wire   [2:0] b10_in1;
  wire   [2:0] b0_outmx;
  wire   [2:0] b1_outmx;
  wire   [2:0] b2_outmx;
  wire   [2:0] b3_outmx;
  wire   [2:0] b4_outmx;
  wire   [2:0] b5_outmx;
  wire   [2:0] b6_outmx;
  wire   [2:0] b7_outmx;
  wire   [2:0] b8_outmx;
  wire   [2:0] b9_outmx;
  wire   [2:0] b10_outmx;
  wire   [2:0] b11_outmx;
  wire   [2:0] b12_outmx;
  wire   [2:0] b13_outmx;
  wire   [2:0] b14_outmx;
  wire   [2:0] b15_outmx;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  mul_bodec_0 encode0_a ( .x(1'b0), .b(b_in[15:0]), .b0(b0_in0), .b1(b1_in0), 
        .b2(b2_in0), .b3(b3_in0), .b4(b4_in0), .b5(b5_in0), .b6(b6_in0), .b7(
        b7_in0) );
  mul_bodec_3 encode0_b ( .x(b_in[15]), .b(b_in[31:16]), .b0(b8_in0), .b1(
        b9_in0), .b2(b10_in0), .b3(b11_in0), .b4(b12_in0), .b5(b13_in0), .b6(
        b14_in0), .b7(b15_in0) );
  clken_buf_2 ckbuf_0 ( .clk(clk_enb0), .rclk(clk), .enb_l(n2), .tmb_l(tm_l)
         );
  clken_buf_1 ckbuf_1 ( .clk(clk_enb1), .rclk(clk), .enb_l(n3), .tmb_l(tm_l)
         );
  dff_SIZE1_2 hld_dff0 ( .din(b_in[31]), .clk(clk_enb1), .q(b[31]), .se(se), 
        .si(1'b0) );
  dff_SIZE32_1 hld_dff ( .din({net210921, net210922, net210923, net210924, 
        net210925, net210926, net210927, net210928, net210929, net210930, 
        net210931, b_in[52:32]}), .clk(clk_enb1), .q({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, b[52:32]}), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  mul_bodec_2 encode1_a ( .x(b[31]), .b(b[47:32]), .b0(b0_in1), .b1(b1_in1), 
        .b2(b2_in1), .b3(b3_in1), .b4(b4_in1), .b5(b5_in1), .b6(b6_in1), .b7(
        b7_in1) );
  mul_bodec_1 encode1_b ( .x(b[47]), .b({net210910, net210911, net210912, 
        net210913, net210914, net210915, net210916, net210917, net210918, 
        net210919, net210920, b[52:48]}), .b0(b8_in1), .b1(b9_in1), .b2({
        SYNOPSYS_UNCONNECTED__11, b10_in1[1:0]}) );
  dp_mux2es_SIZE3_0 out_mux0 ( .dout(b0_outmx), .in0(b0_in0), .in1(b0_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_15 out_mux1 ( .dout(b1_outmx), .in0(b1_in0), .in1(b1_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_14 out_mux2 ( .dout(b2_outmx), .in0(b2_in0), .in1(b2_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_13 out_mux3 ( .dout(b3_outmx), .in0(b3_in0), .in1(b3_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_12 out_mux4 ( .dout(b4_outmx), .in0(b4_in0), .in1(b4_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_11 out_mux5 ( .dout(b5_outmx), .in0(b5_in0), .in1(b5_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_10 out_mux6 ( .dout(b6_outmx), .in0(b6_in0), .in1(b6_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_9 out_mux7 ( .dout(b7_outmx), .in0(b7_in0), .in1(b7_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_8 out_mux8 ( .dout(b8_outmx), .in0(b8_in0), .in1(b8_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_7 out_mux9 ( .dout(b9_outmx), .in0(b9_in0), .in1(b9_in1), 
        .sel(n1) );
  dp_mux2es_SIZE3_6 out_mux10 ( .dout(b10_outmx), .in0(b10_in0), .in1({
        net210909, b10_in1[1:0]}), .sel(n1) );
  dp_mux2es_SIZE3_5 out_mux11 ( .dout(b11_outmx), .in0(b11_in0), .in1({
        net210906, net210907, net210908}), .sel(n1) );
  dp_mux2es_SIZE3_4 out_mux12 ( .dout(b12_outmx), .in0(b12_in0), .in1({
        net210903, net210904, net210905}), .sel(n1) );
  dp_mux2es_SIZE3_3 out_mux13 ( .dout(b13_outmx), .in0(b13_in0), .in1({
        net210900, net210901, net210902}), .sel(n1) );
  dp_mux2es_SIZE3_2 out_mux14 ( .dout(b14_outmx), .in0(b14_in0), .in1({
        net210897, net210898, net210899}), .sel(n1) );
  dp_mux2es_SIZE3_1 out_mux15 ( .dout(b15_outmx), .in0(b15_in0), .in1({
        net210894, net210895, net210896}), .sel(n1) );
  dff_SIZE3_16 out_dff0 ( .din(b0_outmx), .clk(clk_enb0), .q(b0), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_15 out_dff1 ( .din(b1_outmx), .clk(clk_enb0), .q(b1), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_14 out_dff2 ( .din(b2_outmx), .clk(clk_enb0), .q(b2), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_13 out_dff3 ( .din(b3_outmx), .clk(clk_enb0), .q(b3), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_12 out_dff4 ( .din(b4_outmx), .clk(clk_enb0), .q(b4), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_11 out_dff5 ( .din(b5_outmx), .clk(clk_enb0), .q(b5), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_10 out_dff6 ( .din(b6_outmx), .clk(clk_enb0), .q(b6), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_9 out_dff7 ( .din(b7_outmx), .clk(clk_enb0), .q(b7), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_8 out_dff8 ( .din(b8_outmx), .clk(clk_enb0), .q(b8), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_7 out_dff9 ( .din(b9_outmx), .clk(clk_enb0), .q(b9), .se(se), .si(
        {1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_6 out_dff10 ( .din(b10_outmx), .clk(clk_enb0), .q(b10), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_5 out_dff11 ( .din(b11_outmx), .clk(clk_enb0), .q(b11), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_4 out_dff12 ( .din(b12_outmx), .clk(clk_enb0), .q(b12), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_3 out_dff13 ( .din(b13_outmx), .clk(clk_enb0), .q(b13), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_2 out_dff14 ( .din(b14_outmx), .clk(clk_enb0), .q(b14), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE3_1 out_dff15 ( .din(b15_outmx), .clk(clk_enb0), .q(b15), .se(se), 
        .si({1'b0, 1'b0, 1'b0}) );
  INVX0_RVT U2 ( .A(mul_step), .Y(n2) );
  INVX1_RVT U3 ( .A(head), .Y(n1) );
  NAND2X0_RVT U5 ( .A1(head), .A2(mul_step), .Y(n3) );
endmodule


module mul_negen_0 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa42_0 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa32_0 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ha_0 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ppgensign_0 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1148 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1149 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_393 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_394 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_395 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   a;
  assign cout = a;

  INVX1_RVT U1 ( .A(a), .Y(sum) );
endmodule


module mul_csa32_396 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   a;
  assign sum = a;

endmodule


module mul_ppgensign_16 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_0 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net42, net47, p1_l_65, net38, net0118, p1_l_64, net43, net48,
         net210534, net210535, net210536, net210537;
  assign sum[5] = 1'b0;

  mul_ppgensign_0 p0_64_ ( .p_l(net42), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_16 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ppgen_1149 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_1148 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_csa32_396 sc1_67_ ( .sum(sum[3]), .a(net0118), .b(1'b0), .c(net210537)
         );
  mul_csa32_395 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(1'b1), 
        .c(net210536) );
  mul_csa32_394 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net210535) );
  mul_csa32_393 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net210534) );
endmodule


module mul_ppgen_1144 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1145 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_392 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_0 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210533;

  mul_csa32_392 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210533) );
  mul_ppgen_1145 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1144 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_961 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_962 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_963 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_964 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_965 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_966 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_11 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_11 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_12 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_331 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_332 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_0 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_12 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_11 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_332 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_331 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_11 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_966 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_965 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_964 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(
        p0_l_1) );
  mul_ppgen_963 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(
        p0_l_0) );
  mul_ppgen_962 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_961 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_967 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_968 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_333 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_301 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210199;

  mul_csa32_333 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210199) );
  mul_ppgen_968 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_967 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_970 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_971 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_334 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_302 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210198;

  mul_csa32_334 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210198) );
  mul_ppgen_971 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_970 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_973 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_974 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_335 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_303 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210197;

  mul_csa32_335 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210197) );
  mul_ppgen_974 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_973 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_976 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_977 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_336 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_304 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210196;

  mul_csa32_336 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210196) );
  mul_ppgen_977 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_976 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_979 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_980 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_337 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_305 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210195;

  mul_csa32_337 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210195) );
  mul_ppgen_980 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_979 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_982 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_983 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_338 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_306 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210194;

  mul_csa32_338 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210194) );
  mul_ppgen_983 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_982 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_985 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_986 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_339 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_307 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210193;

  mul_csa32_339 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210193) );
  mul_ppgen_986 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_985 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_988 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_989 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_340 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_308 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210192;

  mul_csa32_340 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210192) );
  mul_ppgen_989 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_988 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_991 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_992 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_341 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_309 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210191;

  mul_csa32_341 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210191) );
  mul_ppgen_992 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_991 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_994 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_995 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_342 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_310 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210190;

  mul_csa32_342 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210190) );
  mul_ppgen_995 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_994 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_997 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_998 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_343 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_311 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210189;

  mul_csa32_343 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210189) );
  mul_ppgen_998 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_997 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1000 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1001 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_344 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_312 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210188;

  mul_csa32_344 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210188) );
  mul_ppgen_1001 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1000 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1003 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1004 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_345 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_313 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210187;

  mul_csa32_345 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210187) );
  mul_ppgen_1004 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1003 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1006 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1007 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_346 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_314 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210186;

  mul_csa32_346 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210186) );
  mul_ppgen_1007 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1006 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1009 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1010 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_347 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_315 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210185;

  mul_csa32_347 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210185) );
  mul_ppgen_1010 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1009 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1012 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1013 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_348 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_316 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210184;

  mul_csa32_348 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210184) );
  mul_ppgen_1013 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1012 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1015 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1016 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_349 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_317 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210183;

  mul_csa32_349 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210183) );
  mul_ppgen_1016 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1015 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1018 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1019 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_350 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_318 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210182;

  mul_csa32_350 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210182) );
  mul_ppgen_1019 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1018 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1021 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1022 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_351 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_319 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210181;

  mul_csa32_351 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210181) );
  mul_ppgen_1022 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1021 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1024 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1025 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_352 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_320 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210180;

  mul_csa32_352 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210180) );
  mul_ppgen_1025 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1024 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1027 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1028 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_353 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_321 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210179;

  mul_csa32_353 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210179) );
  mul_ppgen_1028 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1027 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1030 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1031 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_354 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_322 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210178;

  mul_csa32_354 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210178) );
  mul_ppgen_1031 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1030 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1033 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1034 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_355 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_323 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210177;

  mul_csa32_355 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210177) );
  mul_ppgen_1034 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1033 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1036 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1037 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_356 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_324 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210176;

  mul_csa32_356 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210176) );
  mul_ppgen_1037 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1036 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1039 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1040 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_357 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_325 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210175;

  mul_csa32_357 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210175) );
  mul_ppgen_1040 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1039 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1042 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1043 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_358 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_326 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210174;

  mul_csa32_358 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210174) );
  mul_ppgen_1043 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1042 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1045 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1046 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_359 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_327 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210173;

  mul_csa32_359 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210173) );
  mul_ppgen_1046 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1045 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1048 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1049 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_360 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_328 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210172;

  mul_csa32_360 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210172) );
  mul_ppgen_1049 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1048 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1051 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1052 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_361 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_329 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210171;

  mul_csa32_361 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210171) );
  mul_ppgen_1052 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1051 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1054 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1055 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_362 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_330 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210170;

  mul_csa32_362 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210170) );
  mul_ppgen_1055 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1054 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1057 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1058 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_363 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_331 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210169;

  mul_csa32_363 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210169) );
  mul_ppgen_1058 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1057 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1060 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1061 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_364 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_332 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210168;

  mul_csa32_364 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210168) );
  mul_ppgen_1061 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1060 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1063 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1064 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_365 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_333 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210167;

  mul_csa32_365 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210167) );
  mul_ppgen_1064 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1063 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1066 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1067 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_366 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_334 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210166;

  mul_csa32_366 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210166) );
  mul_ppgen_1067 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1066 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1069 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1070 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_367 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_335 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210165;

  mul_csa32_367 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210165) );
  mul_ppgen_1070 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1069 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1072 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1073 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_368 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_336 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210164;

  mul_csa32_368 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210164) );
  mul_ppgen_1073 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1072 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1075 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1076 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_369 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_337 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210163;

  mul_csa32_369 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210163) );
  mul_ppgen_1076 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1075 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1078 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1079 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_370 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_338 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210162;

  mul_csa32_370 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210162) );
  mul_ppgen_1079 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1078 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1081 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1082 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_371 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_339 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210161;

  mul_csa32_371 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210161) );
  mul_ppgen_1082 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1081 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1084 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1085 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_372 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_340 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210160;

  mul_csa32_372 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210160) );
  mul_ppgen_1085 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1084 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1087 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1088 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_373 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_341 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210159;

  mul_csa32_373 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210159) );
  mul_ppgen_1088 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1087 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1090 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1091 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_374 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_342 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210158;

  mul_csa32_374 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210158) );
  mul_ppgen_1091 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1090 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1093 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1094 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_375 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_343 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210157;

  mul_csa32_375 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210157) );
  mul_ppgen_1094 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1093 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1096 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1097 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_376 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_344 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210156;

  mul_csa32_376 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210156) );
  mul_ppgen_1097 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1096 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1099 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1100 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_377 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_345 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210155;

  mul_csa32_377 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210155) );
  mul_ppgen_1100 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1099 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1102 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1103 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_378 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_346 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210154;

  mul_csa32_378 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210154) );
  mul_ppgen_1103 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1102 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1105 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1106 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_379 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_347 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210153;

  mul_csa32_379 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210153) );
  mul_ppgen_1106 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1105 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1108 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1109 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_380 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_348 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210152;

  mul_csa32_380 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210152) );
  mul_ppgen_1109 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1108 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1111 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1112 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_381 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_349 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210151;

  mul_csa32_381 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210151) );
  mul_ppgen_1112 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1111 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1114 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1115 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_382 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_350 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210150;

  mul_csa32_382 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210150) );
  mul_ppgen_1115 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1114 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1117 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1118 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_383 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_351 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210149;

  mul_csa32_383 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210149) );
  mul_ppgen_1118 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1117 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1120 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1121 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_384 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_352 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210148;

  mul_csa32_384 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210148) );
  mul_ppgen_1121 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1120 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1123 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1124 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_385 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_353 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210147;

  mul_csa32_385 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210147) );
  mul_ppgen_1124 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1123 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1126 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1127 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_386 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_354 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210146;

  mul_csa32_386 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210146) );
  mul_ppgen_1127 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1126 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1129 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1130 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_387 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_355 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210145;

  mul_csa32_387 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210145) );
  mul_ppgen_1130 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1129 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1132 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1133 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_388 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_356 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210144;

  mul_csa32_388 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210144) );
  mul_ppgen_1133 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1132 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1135 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1136 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_389 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_357 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210143;

  mul_csa32_389 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210143) );
  mul_ppgen_1136 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1135 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1138 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1139 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_390 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_358 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210142;

  mul_csa32_390 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210142) );
  mul_ppgen_1139 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1138 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_1141 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_1142 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_391 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_359 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210141;

  mul_csa32_391 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210141) );
  mul_ppgen_1142 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_1141 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_0 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210540, net210541, net210542, net210543, net210544, net210545,
         net210546, net210547, net210548, net210549, net210550, net210551,
         net210552, net210553, net210554, net210555, net210556, net210557,
         net210558, net210559, net210560, net210561, net210562, net210563,
         net210564, net210565, net210566, net210567, net210568, net210569,
         net210570, net210571, net210572, net210573, net210574, net210575,
         net210576, net210577, net210578, net210579, net210580, net210581,
         net210582, net210583, net210584, net210585, net210586, net210587,
         net210588, net210589, net210590, net210591, net210592, net210593,
         net210594, net210595, net210596, net210597, net210598, net210599,
         net210600, net210601, net210602, net210603, net210604, net210605,
         net210606, net210607, net210608, net210609, net210610, net210611,
         net210612, net210613, net210614, net210615, net210616, net210617,
         net210618, net210619, net210620, net210621, net210622, net210623,
         net210624, net210625, net210626, net210627, net210628, net210629,
         net210630, net210631, net210632, net210633, net210634, net210635,
         net210636, net210637, net210638, net210639, net210640, net210641,
         net210642, net210643, net210644, net210645, net210646, net210647,
         net210648, net210649, net210650, net210651, net210652, net210653,
         net210654, net210655, net210656, net210657, net210658, net210659,
         net210660, net210661, net210662, net210663, net210664, net210665,
         net210666, net210667, net210668, net210669, net210670, net210671,
         net210672, net210673, net210674, net210675, net210676, net210677,
         net210678, net210679, net210680, net210681, net210682, net210683,
         net210684, net210685, net210686, net210687, net210688, net210689,
         net210690, net210691, net210692, net210693, net210694, net210695,
         net210696, net210697, net210698, net210699, net210700, net210701,
         net210702, net210703, net210704, net210705, net210706, net210707,
         net210708, net210709, net210710, net210711, net210712, net210713,
         net210714, net210715, net210716, net210717, net210718, net210719,
         net210720, net210721, net210722, net210723, net210724, net210725,
         net210726, net210727, net210728, net210729, net210730, net210731,
         net210732, net210733, net210734, net210735, net210736, net210737,
         net210738, net210739, net210740, net210741, net210742, net210743,
         net210744, net210745, net210746, net210747, net210748, net210749,
         net210750, net210751, net210752, net210753, net210754, net210755,
         net210756, net210757, net210758, net210759, net210760, net210761,
         net210762, net210763, net210764, net210765, net210766, net210767,
         net210768, net210769, net210770, net210771, net210772, net210773,
         net210774, net210775, net210776, net210777, net210778, net210779,
         net210780, net210781, net210782, net210783, net210784;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  mul_ppgen3sign_0 I2 ( .cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, cout[66:64]}), .sum({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, sum[67:64]}), .am1(a[63]), .am2(a[62]), .am3(
        a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2({net210779, net210780, 
        net210781}), .bot(net210782), .head(net210783), .p0m1_l(p0_l[63]), 
        .p1m1_l(p1_l[63]), .p2m1_l(net210784) );
  mul_ppgen3_0 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), .b0(b0), .b1(b1), 
        .b2({net210775, net210776, net210777}), .p0m1_l(p0_l[62]), .p1m1_l(
        p1_l[62]), .p2m1_l(net210778) );
  mul_ppgen3_359 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), .b0(b0), .b1(b1), 
        .b2({net210771, net210772, net210773}), .p0m1_l(p0_l[61]), .p1m1_l(
        p1_l[61]), .p2m1_l(net210774) );
  mul_ppgen3_358 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), .b0(b0), .b1(b1), 
        .b2({net210767, net210768, net210769}), .p0m1_l(p0_l[60]), .p1m1_l(
        p1_l[60]), .p2m1_l(net210770) );
  mul_ppgen3_357 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), .b0(b0), .b1(b1), 
        .b2({net210763, net210764, net210765}), .p0m1_l(p0_l[59]), .p1m1_l(
        p1_l[59]), .p2m1_l(net210766) );
  mul_ppgen3_356 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), .b0(b0), .b1(b1), 
        .b2({net210759, net210760, net210761}), .p0m1_l(p0_l[58]), .p1m1_l(
        p1_l[58]), .p2m1_l(net210762) );
  mul_ppgen3_355 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), .b0(b0), .b1(b1), 
        .b2({net210755, net210756, net210757}), .p0m1_l(p0_l[57]), .p1m1_l(
        p1_l[57]), .p2m1_l(net210758) );
  mul_ppgen3_354 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), .b0(b0), .b1(b1), 
        .b2({net210751, net210752, net210753}), .p0m1_l(p0_l[56]), .p1m1_l(
        p1_l[56]), .p2m1_l(net210754) );
  mul_ppgen3_353 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), .b0(b0), .b1(b1), 
        .b2({net210747, net210748, net210749}), .p0m1_l(p0_l[55]), .p1m1_l(
        p1_l[55]), .p2m1_l(net210750) );
  mul_ppgen3_352 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), .b0(b0), .b1(b1), 
        .b2({net210743, net210744, net210745}), .p0m1_l(p0_l[54]), .p1m1_l(
        p1_l[54]), .p2m1_l(net210746) );
  mul_ppgen3_351 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), .b0(b0), .b1(b1), 
        .b2({net210739, net210740, net210741}), .p0m1_l(p0_l[53]), .p1m1_l(
        p1_l[53]), .p2m1_l(net210742) );
  mul_ppgen3_350 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), .b0(b0), .b1(b1), 
        .b2({net210735, net210736, net210737}), .p0m1_l(p0_l[52]), .p1m1_l(
        p1_l[52]), .p2m1_l(net210738) );
  mul_ppgen3_349 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), .b0(b0), .b1(b1), 
        .b2({net210731, net210732, net210733}), .p0m1_l(p0_l[51]), .p1m1_l(
        p1_l[51]), .p2m1_l(net210734) );
  mul_ppgen3_348 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), .b0(b0), .b1(b1), 
        .b2({net210727, net210728, net210729}), .p0m1_l(p0_l[50]), .p1m1_l(
        p1_l[50]), .p2m1_l(net210730) );
  mul_ppgen3_347 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), .b0(b0), .b1(b1), 
        .b2({net210723, net210724, net210725}), .p0m1_l(p0_l[49]), .p1m1_l(
        p1_l[49]), .p2m1_l(net210726) );
  mul_ppgen3_346 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), .b0(b0), .b1(b1), 
        .b2({net210719, net210720, net210721}), .p0m1_l(p0_l[48]), .p1m1_l(
        p1_l[48]), .p2m1_l(net210722) );
  mul_ppgen3_345 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), .b0(b0), .b1(b1), 
        .b2({net210715, net210716, net210717}), .p0m1_l(p0_l[47]), .p1m1_l(
        p1_l[47]), .p2m1_l(net210718) );
  mul_ppgen3_344 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), .b0(b0), .b1(b1), 
        .b2({net210711, net210712, net210713}), .p0m1_l(p0_l[46]), .p1m1_l(
        p1_l[46]), .p2m1_l(net210714) );
  mul_ppgen3_343 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), .b0(b0), .b1(b1), 
        .b2({net210707, net210708, net210709}), .p0m1_l(p0_l[45]), .p1m1_l(
        p1_l[45]), .p2m1_l(net210710) );
  mul_ppgen3_342 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), .b0(b0), .b1(b1), 
        .b2({net210703, net210704, net210705}), .p0m1_l(p0_l[44]), .p1m1_l(
        p1_l[44]), .p2m1_l(net210706) );
  mul_ppgen3_341 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), .b0(b0), .b1(b1), 
        .b2({net210699, net210700, net210701}), .p0m1_l(p0_l[43]), .p1m1_l(
        p1_l[43]), .p2m1_l(net210702) );
  mul_ppgen3_340 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), .b0(b0), .b1(b1), 
        .b2({net210695, net210696, net210697}), .p0m1_l(p0_l[42]), .p1m1_l(
        p1_l[42]), .p2m1_l(net210698) );
  mul_ppgen3_339 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), .b0(b0), .b1(b1), 
        .b2({net210691, net210692, net210693}), .p0m1_l(p0_l[41]), .p1m1_l(
        p1_l[41]), .p2m1_l(net210694) );
  mul_ppgen3_338 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), .b0(b0), .b1(b1), 
        .b2({net210687, net210688, net210689}), .p0m1_l(p0_l[40]), .p1m1_l(
        p1_l[40]), .p2m1_l(net210690) );
  mul_ppgen3_337 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), .b0(b0), .b1(b1), 
        .b2({net210683, net210684, net210685}), .p0m1_l(p0_l[39]), .p1m1_l(
        p1_l[39]), .p2m1_l(net210686) );
  mul_ppgen3_336 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), .b0(b0), .b1(b1), 
        .b2({net210679, net210680, net210681}), .p0m1_l(p0_l[38]), .p1m1_l(
        p1_l[38]), .p2m1_l(net210682) );
  mul_ppgen3_335 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), .b0(b0), .b1(b1), 
        .b2({net210675, net210676, net210677}), .p0m1_l(p0_l[37]), .p1m1_l(
        p1_l[37]), .p2m1_l(net210678) );
  mul_ppgen3_334 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), .b0(b0), .b1(b1), 
        .b2({net210671, net210672, net210673}), .p0m1_l(p0_l[36]), .p1m1_l(
        p1_l[36]), .p2m1_l(net210674) );
  mul_ppgen3_333 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), .b0(b0), .b1(b1), 
        .b2({net210667, net210668, net210669}), .p0m1_l(p0_l[35]), .p1m1_l(
        p1_l[35]), .p2m1_l(net210670) );
  mul_ppgen3_332 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), .b0(b0), .b1(b1), 
        .b2({net210663, net210664, net210665}), .p0m1_l(p0_l[34]), .p1m1_l(
        p1_l[34]), .p2m1_l(net210666) );
  mul_ppgen3_331 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), .b0(b0), .b1(b1), 
        .b2({net210659, net210660, net210661}), .p0m1_l(p0_l[33]), .p1m1_l(
        p1_l[33]), .p2m1_l(net210662) );
  mul_ppgen3_330 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), .b0(b0), .b1(b1), 
        .b2({net210655, net210656, net210657}), .p0m1_l(p0_l[32]), .p1m1_l(
        p1_l[32]), .p2m1_l(net210658) );
  mul_ppgen3_329 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), .b0(b0), .b1(b1), 
        .b2({net210651, net210652, net210653}), .p0m1_l(p0_l[31]), .p1m1_l(
        p1_l[31]), .p2m1_l(net210654) );
  mul_ppgen3_328 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), .b0(b0), .b1(b1), 
        .b2({net210647, net210648, net210649}), .p0m1_l(p0_l[30]), .p1m1_l(
        p1_l[30]), .p2m1_l(net210650) );
  mul_ppgen3_327 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), .b0(b0), .b1(b1), 
        .b2({net210643, net210644, net210645}), .p0m1_l(p0_l[29]), .p1m1_l(
        p1_l[29]), .p2m1_l(net210646) );
  mul_ppgen3_326 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), .b0(b0), .b1(b1), 
        .b2({net210639, net210640, net210641}), .p0m1_l(p0_l[28]), .p1m1_l(
        p1_l[28]), .p2m1_l(net210642) );
  mul_ppgen3_325 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), .b0(b0), .b1(b1), 
        .b2({net210635, net210636, net210637}), .p0m1_l(p0_l[27]), .p1m1_l(
        p1_l[27]), .p2m1_l(net210638) );
  mul_ppgen3_324 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), .b0(b0), .b1(b1), 
        .b2({net210631, net210632, net210633}), .p0m1_l(p0_l[26]), .p1m1_l(
        p1_l[26]), .p2m1_l(net210634) );
  mul_ppgen3_323 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), .b0(b0), .b1(b1), 
        .b2({net210627, net210628, net210629}), .p0m1_l(p0_l[25]), .p1m1_l(
        p1_l[25]), .p2m1_l(net210630) );
  mul_ppgen3_322 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), .b0(b0), .b1(b1), 
        .b2({net210623, net210624, net210625}), .p0m1_l(p0_l[24]), .p1m1_l(
        p1_l[24]), .p2m1_l(net210626) );
  mul_ppgen3_321 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), .b0(b0), .b1(b1), 
        .b2({net210619, net210620, net210621}), .p0m1_l(p0_l[23]), .p1m1_l(
        p1_l[23]), .p2m1_l(net210622) );
  mul_ppgen3_320 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), .b0(b0), .b1(b1), 
        .b2({net210615, net210616, net210617}), .p0m1_l(p0_l[22]), .p1m1_l(
        p1_l[22]), .p2m1_l(net210618) );
  mul_ppgen3_319 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), .b0(b0), .b1(b1), 
        .b2({net210611, net210612, net210613}), .p0m1_l(p0_l[21]), .p1m1_l(
        p1_l[21]), .p2m1_l(net210614) );
  mul_ppgen3_318 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), .b0(b0), .b1(b1), 
        .b2({net210607, net210608, net210609}), .p0m1_l(p0_l[20]), .p1m1_l(
        p1_l[20]), .p2m1_l(net210610) );
  mul_ppgen3_317 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), .b0(b0), .b1(b1), 
        .b2({net210603, net210604, net210605}), .p0m1_l(p0_l[19]), .p1m1_l(
        p1_l[19]), .p2m1_l(net210606) );
  mul_ppgen3_316 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), .b0(b0), .b1(b1), 
        .b2({net210599, net210600, net210601}), .p0m1_l(p0_l[18]), .p1m1_l(
        p1_l[18]), .p2m1_l(net210602) );
  mul_ppgen3_315 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), .b0(b0), .b1(b1), 
        .b2({net210595, net210596, net210597}), .p0m1_l(p0_l[17]), .p1m1_l(
        p1_l[17]), .p2m1_l(net210598) );
  mul_ppgen3_314 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), .b0(b0), .b1(b1), 
        .b2({net210591, net210592, net210593}), .p0m1_l(p0_l[16]), .p1m1_l(
        p1_l[16]), .p2m1_l(net210594) );
  mul_ppgen3_313 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), .b0(b0), .b1(b1), 
        .b2({net210587, net210588, net210589}), .p0m1_l(p0_l[15]), .p1m1_l(
        p1_l[15]), .p2m1_l(net210590) );
  mul_ppgen3_312 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), .b0(b0), .b1(b1), 
        .b2({net210583, net210584, net210585}), .p0m1_l(p0_l[14]), .p1m1_l(
        p1_l[14]), .p2m1_l(net210586) );
  mul_ppgen3_311 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), .b0(b0), .b1(b1), 
        .b2({net210579, net210580, net210581}), .p0m1_l(p0_l[13]), .p1m1_l(
        p1_l[13]), .p2m1_l(net210582) );
  mul_ppgen3_310 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), .b0(b0), .b1(b1), 
        .b2({net210575, net210576, net210577}), .p0m1_l(p0_l[12]), .p1m1_l(
        p1_l[12]), .p2m1_l(net210578) );
  mul_ppgen3_309 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), .b0(b0), .b1(b1), 
        .b2({net210571, net210572, net210573}), .p0m1_l(p0_l[11]), .p1m1_l(
        p1_l[11]), .p2m1_l(net210574) );
  mul_ppgen3_308 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), .b0(b0), .b1(b1), 
        .b2({net210567, net210568, net210569}), .p0m1_l(p0_l[10]), .p1m1_l(
        p1_l[10]), .p2m1_l(net210570) );
  mul_ppgen3_307 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), .b0(b0), .b1(b1), 
        .b2({net210563, net210564, net210565}), .p0m1_l(p0_l[9]), .p1m1_l(
        p1_l[9]), .p2m1_l(net210566) );
  mul_ppgen3_306 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), .sum(
        sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), .b1(b1), .b2({
        net210559, net210560, net210561}), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), 
        .p2m1_l(net210562) );
  mul_ppgen3_305 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), .sum(
        sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), .b1(b1), .b2({
        net210555, net210556, net210557}), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), 
        .p2m1_l(net210558) );
  mul_ppgen3_304 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), .sum(
        sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), .b1(b1), .b2({
        net210551, net210552, net210553}), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), 
        .p2m1_l(net210554) );
  mul_ppgen3_303 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), .sum(
        sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), .b1(b1), .b2({
        net210547, net210548, net210549}), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), 
        .p2m1_l(net210550) );
  mul_ppgen3_302 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), .sum(
        sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), .b1(b1), .b2({
        net210543, net210544, net210545}), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), 
        .p2m1_l(net210546) );
  mul_ppgen3_301 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), .sum(
        sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), .b1(b1), .b2({
        net210540, net210541, net210542}), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), 
        .p2m1_l(1'b1) );
  mul_ppgen3lsb4_0 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ppgen_763 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_764 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_765 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_766 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_767 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_768 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_8 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_csa32_261 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_262 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_263 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_264 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgensign_10 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_11 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_12 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_4 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net088, net0117, net42, net47, p2_l_67, net073, p1_l_65, net38,
         net0118, p2_l_66, net078, p2_l_65, net8, p2_l_64, net15, p1_l_64,
         net43, net48, net35, n1;

  mul_ppgensign_12 p0_64_ ( .p_l(net088), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_11 p2_68_ ( .p_l(sum[5]), .z(net073), .b(b2), .pm1_l(p2_l_67)
         );
  mul_ppgensign_10 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ha_8 sc1_68_ ( .cout(cout[4]), .sum(sum[4]), .a(1'b1), .b(net073) );
  mul_ppgen_768 p2_67_ ( .p_l(p2_l_67), .z(net078), .a(am1), .b(b2), .pm1_l(
        p2_l_66) );
  mul_ppgen_767 p2_66_ ( .p_l(p2_l_66), .z(net8), .a(am2), .b(b2), .pm1_l(
        p2_l_65) );
  mul_ppgen_766 p2_65_ ( .p_l(p2_l_65), .z(net15), .a(am3), .b(b2), .pm1_l(
        p2_l_64) );
  mul_ppgen_765 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_764 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_ppgen_763 p2_64_ ( .p_l(p2_l_64), .z(net35), .a(am4), .b(b2), .pm1_l(
        p2m1_l) );
  mul_csa32_264 sc1_67_ ( .sum(sum[3]), .cout(cout[3]), .a(net0118), .b(
        net0117), .c(net078) );
  mul_csa32_263 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(n1), .c(
        net8) );
  mul_csa32_262 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net15) );
  mul_csa32_261 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net35) );
  NAND2X0_RVT U2 ( .A1(net088), .A2(head), .Y(n1) );
  INVX1_RVT U3 ( .A(n1), .Y(net0117) );
  OA21X1_RVT U5 ( .A1(net088), .A2(head), .A3(n1), .Y(net42) );
endmodule


module mul_ppgen_577 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_578 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_579 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_580 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_581 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_582 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_7 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_7 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_8 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_199 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_200 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_4 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_8 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_7 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_200 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_199 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_7 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_582 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_581 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_580 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(
        p0_l_1) );
  mul_ppgen_579 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(
        p0_l_0) );
  mul_ppgen_578 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_577 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_583 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_584 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_585 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_csa32_201 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_181 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043, net210201;

  mul_csa32_201 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_585 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(net210201) );
  mul_ppgen_584 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_583 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_586 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_587 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_588 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_202 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_182 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_202 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_588 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_587 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_586 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_589 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_590 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_591 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_203 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_183 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_203 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_591 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_590 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_589 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_592 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_593 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_594 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_204 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_184 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_204 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_594 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_593 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_592 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_595 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_596 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_597 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_205 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_185 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_205 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_597 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_596 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_595 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_598 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_599 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_600 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_206 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_186 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_206 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_600 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_599 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_598 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_601 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_602 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_603 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_207 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_187 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_207 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_603 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_602 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_601 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_604 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_605 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_606 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_208 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_188 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_208 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_606 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_605 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_604 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_607 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_608 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_609 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_209 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_189 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_209 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_609 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_608 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_607 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_610 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_611 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_612 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_210 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_190 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_210 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_612 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_611 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_610 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_613 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_614 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_615 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_211 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_191 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_211 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_615 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_614 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_613 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_616 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_617 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_618 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_212 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_192 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_212 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_618 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_617 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_616 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_619 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_620 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_621 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_213 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_193 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_213 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_621 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_620 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_619 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_622 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_623 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_624 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_214 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_194 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_214 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_624 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_623 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_622 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_625 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_626 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_627 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_215 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_195 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_215 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_627 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_626 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_625 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_628 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_629 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_630 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_216 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_196 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_216 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_630 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_629 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_628 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_631 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_632 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_633 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_217 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_197 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_217 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_633 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_632 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_631 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_634 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_635 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_636 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_218 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_198 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_218 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_636 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_635 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_634 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_637 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_638 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_639 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_219 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_199 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_219 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_639 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_638 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_637 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_640 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_641 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_642 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_220 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_200 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_220 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_642 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_641 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_640 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_643 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_644 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_645 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_221 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_201 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_221 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_645 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_644 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_643 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_646 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_647 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_648 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_222 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_202 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_222 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_648 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_647 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_646 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_649 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_650 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_651 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_223 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_203 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_223 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_651 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_650 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_649 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_652 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_653 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_654 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_224 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_204 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_224 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_654 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_653 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_652 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_655 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_656 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_657 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_225 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_205 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_225 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_657 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_656 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_655 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_658 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_659 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_660 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_226 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_206 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_226 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_660 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_659 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_658 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_661 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_662 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_663 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_227 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_207 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_227 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_663 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_662 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_661 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_664 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_665 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_666 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_228 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_208 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_228 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_666 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_665 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_664 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_667 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_668 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_669 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_229 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_209 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_229 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_669 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_668 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_667 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_670 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_671 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_672 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_230 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_210 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_230 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_672 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_671 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_670 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_673 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_674 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_675 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_231 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_211 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_231 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_675 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_674 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_673 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_676 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_677 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_678 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_232 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_212 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_232 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_678 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_677 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_676 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_679 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_680 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_681 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_233 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_213 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_233 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_681 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_680 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_679 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_682 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_683 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_684 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_234 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_214 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_234 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_684 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_683 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_682 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_685 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_686 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_687 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_235 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_215 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_235 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_687 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_686 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_685 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_688 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_689 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_690 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_236 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_216 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_236 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_690 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_689 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_688 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_691 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_692 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_693 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_237 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_217 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_237 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_693 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_692 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_691 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_694 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_695 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_696 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_238 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_218 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_238 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_696 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_695 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_694 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_697 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_698 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_699 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_239 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_219 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_239 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_699 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_698 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_697 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_700 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_701 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_702 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_240 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_220 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_240 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_702 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_701 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_700 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_703 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_704 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_705 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_241 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_221 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_241 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_705 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_704 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_703 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_706 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_707 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_708 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_242 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_222 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_242 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_708 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_707 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_706 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_709 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_710 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_711 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_243 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_223 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_243 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_711 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_710 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_709 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_712 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_713 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_714 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_244 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_224 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_244 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_714 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_713 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_712 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_715 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_716 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_717 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_245 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_225 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_245 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_717 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_716 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_715 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_718 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_719 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_720 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_246 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_226 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_246 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_720 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_719 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_718 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_721 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_722 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_723 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_247 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_227 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_247 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_723 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_722 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_721 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_724 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_725 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_726 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_248 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_228 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_248 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_726 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_725 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_724 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_727 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_728 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_729 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_249 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_229 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_249 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_729 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_728 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_727 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_730 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_731 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_732 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_250 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_230 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_250 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_732 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_731 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_730 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_733 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_734 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_735 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_251 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_231 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_251 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_735 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_734 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_733 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_736 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_737 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_738 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_252 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_232 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_252 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_738 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_737 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_736 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_739 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_740 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_741 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_253 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_233 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_253 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_741 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_740 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_739 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_742 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_743 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_744 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_254 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_234 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_254 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_744 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_743 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_742 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_745 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_746 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_747 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_255 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_235 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_255 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_747 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_746 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_745 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_748 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_749 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_750 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_256 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_236 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_256 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_750 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_749 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_748 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_751 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_752 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_753 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_257 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_237 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_257 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_753 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_752 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_751 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_754 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_755 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_756 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_258 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_238 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_258 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_756 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_755 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_754 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_757 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_758 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_759 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_259 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_239 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_259 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_759 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_758 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_757 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_760 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_761 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_762 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_260 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_240 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_260 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_762 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_761 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_760 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_4 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210279;
  wire   [63:4] p2_l;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;

  mul_ppgen3sign_4 I2 ( .cout(cout[68:64]), .sum(sum[69:64]), .am1(a[63]), 
        .am2(a[62]), .am3(a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2(b2), 
        .bot(net210279), .head(head), .p0m1_l(p0_l[63]), .p1m1_l(p1_l[63]), 
        .p2m1_l(p2_l[63]) );
  mul_ppgen3_240 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .p2_l(p2_l[63]), .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[62]), .p1m1_l(p1_l[62]), 
        .p2m1_l(p2_l[62]) );
  mul_ppgen3_239 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .p2_l(p2_l[62]), .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[61]), .p1m1_l(p1_l[61]), 
        .p2m1_l(p2_l[61]) );
  mul_ppgen3_238 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .p2_l(p2_l[61]), .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[60]), .p1m1_l(p1_l[60]), 
        .p2m1_l(p2_l[60]) );
  mul_ppgen3_237 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .p2_l(p2_l[60]), .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[59]), .p1m1_l(p1_l[59]), 
        .p2m1_l(p2_l[59]) );
  mul_ppgen3_236 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .p2_l(p2_l[59]), .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[58]), .p1m1_l(p1_l[58]), 
        .p2m1_l(p2_l[58]) );
  mul_ppgen3_235 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .p2_l(p2_l[58]), .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[57]), .p1m1_l(p1_l[57]), 
        .p2m1_l(p2_l[57]) );
  mul_ppgen3_234 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .p2_l(p2_l[57]), .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[56]), .p1m1_l(p1_l[56]), 
        .p2m1_l(p2_l[56]) );
  mul_ppgen3_233 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .p2_l(p2_l[56]), .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[55]), .p1m1_l(p1_l[55]), 
        .p2m1_l(p2_l[55]) );
  mul_ppgen3_232 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .p2_l(p2_l[55]), .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[54]), .p1m1_l(p1_l[54]), 
        .p2m1_l(p2_l[54]) );
  mul_ppgen3_231 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .p2_l(p2_l[54]), .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[53]), .p1m1_l(p1_l[53]), 
        .p2m1_l(p2_l[53]) );
  mul_ppgen3_230 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .p2_l(p2_l[53]), .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[52]), .p1m1_l(p1_l[52]), 
        .p2m1_l(p2_l[52]) );
  mul_ppgen3_229 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .p2_l(p2_l[52]), .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[51]), .p1m1_l(p1_l[51]), 
        .p2m1_l(p2_l[51]) );
  mul_ppgen3_228 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .p2_l(p2_l[51]), .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[50]), .p1m1_l(p1_l[50]), 
        .p2m1_l(p2_l[50]) );
  mul_ppgen3_227 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .p2_l(p2_l[50]), .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[49]), .p1m1_l(p1_l[49]), 
        .p2m1_l(p2_l[49]) );
  mul_ppgen3_226 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .p2_l(p2_l[49]), .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[48]), .p1m1_l(p1_l[48]), 
        .p2m1_l(p2_l[48]) );
  mul_ppgen3_225 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .p2_l(p2_l[48]), .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[47]), .p1m1_l(p1_l[47]), 
        .p2m1_l(p2_l[47]) );
  mul_ppgen3_224 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .p2_l(p2_l[47]), .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[46]), .p1m1_l(p1_l[46]), 
        .p2m1_l(p2_l[46]) );
  mul_ppgen3_223 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .p2_l(p2_l[46]), .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[45]), .p1m1_l(p1_l[45]), 
        .p2m1_l(p2_l[45]) );
  mul_ppgen3_222 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .p2_l(p2_l[45]), .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[44]), .p1m1_l(p1_l[44]), 
        .p2m1_l(p2_l[44]) );
  mul_ppgen3_221 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .p2_l(p2_l[44]), .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[43]), .p1m1_l(p1_l[43]), 
        .p2m1_l(p2_l[43]) );
  mul_ppgen3_220 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .p2_l(p2_l[43]), .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[42]), .p1m1_l(p1_l[42]), 
        .p2m1_l(p2_l[42]) );
  mul_ppgen3_219 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .p2_l(p2_l[42]), .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[41]), .p1m1_l(p1_l[41]), 
        .p2m1_l(p2_l[41]) );
  mul_ppgen3_218 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .p2_l(p2_l[41]), .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[40]), .p1m1_l(p1_l[40]), 
        .p2m1_l(p2_l[40]) );
  mul_ppgen3_217 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .p2_l(p2_l[40]), .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[39]), .p1m1_l(p1_l[39]), 
        .p2m1_l(p2_l[39]) );
  mul_ppgen3_216 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .p2_l(p2_l[39]), .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[38]), .p1m1_l(p1_l[38]), 
        .p2m1_l(p2_l[38]) );
  mul_ppgen3_215 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .p2_l(p2_l[38]), .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[37]), .p1m1_l(p1_l[37]), 
        .p2m1_l(p2_l[37]) );
  mul_ppgen3_214 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .p2_l(p2_l[37]), .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[36]), .p1m1_l(p1_l[36]), 
        .p2m1_l(p2_l[36]) );
  mul_ppgen3_213 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .p2_l(p2_l[36]), .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[35]), .p1m1_l(p1_l[35]), 
        .p2m1_l(p2_l[35]) );
  mul_ppgen3_212 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .p2_l(p2_l[35]), .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[34]), .p1m1_l(p1_l[34]), 
        .p2m1_l(p2_l[34]) );
  mul_ppgen3_211 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .p2_l(p2_l[34]), .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[33]), .p1m1_l(p1_l[33]), 
        .p2m1_l(p2_l[33]) );
  mul_ppgen3_210 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .p2_l(p2_l[33]), .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[32]), .p1m1_l(p1_l[32]), 
        .p2m1_l(p2_l[32]) );
  mul_ppgen3_209 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .p2_l(p2_l[32]), .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[31]), .p1m1_l(p1_l[31]), 
        .p2m1_l(p2_l[31]) );
  mul_ppgen3_208 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .p2_l(p2_l[31]), .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[30]), .p1m1_l(p1_l[30]), 
        .p2m1_l(p2_l[30]) );
  mul_ppgen3_207 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .p2_l(p2_l[30]), .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[29]), .p1m1_l(p1_l[29]), 
        .p2m1_l(p2_l[29]) );
  mul_ppgen3_206 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .p2_l(p2_l[29]), .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[28]), .p1m1_l(p1_l[28]), 
        .p2m1_l(p2_l[28]) );
  mul_ppgen3_205 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .p2_l(p2_l[28]), .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[27]), .p1m1_l(p1_l[27]), 
        .p2m1_l(p2_l[27]) );
  mul_ppgen3_204 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .p2_l(p2_l[27]), .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[26]), .p1m1_l(p1_l[26]), 
        .p2m1_l(p2_l[26]) );
  mul_ppgen3_203 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .p2_l(p2_l[26]), .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[25]), .p1m1_l(p1_l[25]), 
        .p2m1_l(p2_l[25]) );
  mul_ppgen3_202 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .p2_l(p2_l[25]), .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[24]), .p1m1_l(p1_l[24]), 
        .p2m1_l(p2_l[24]) );
  mul_ppgen3_201 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .p2_l(p2_l[24]), .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[23]), .p1m1_l(p1_l[23]), 
        .p2m1_l(p2_l[23]) );
  mul_ppgen3_200 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .p2_l(p2_l[23]), .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[22]), .p1m1_l(p1_l[22]), 
        .p2m1_l(p2_l[22]) );
  mul_ppgen3_199 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .p2_l(p2_l[22]), .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[21]), .p1m1_l(p1_l[21]), 
        .p2m1_l(p2_l[21]) );
  mul_ppgen3_198 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .p2_l(p2_l[21]), .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[20]), .p1m1_l(p1_l[20]), 
        .p2m1_l(p2_l[20]) );
  mul_ppgen3_197 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .p2_l(p2_l[20]), .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[19]), .p1m1_l(p1_l[19]), 
        .p2m1_l(p2_l[19]) );
  mul_ppgen3_196 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .p2_l(p2_l[19]), .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[18]), .p1m1_l(p1_l[18]), 
        .p2m1_l(p2_l[18]) );
  mul_ppgen3_195 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .p2_l(p2_l[18]), .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[17]), .p1m1_l(p1_l[17]), 
        .p2m1_l(p2_l[17]) );
  mul_ppgen3_194 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .p2_l(p2_l[17]), .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[16]), .p1m1_l(p1_l[16]), 
        .p2m1_l(p2_l[16]) );
  mul_ppgen3_193 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .p2_l(p2_l[16]), .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[15]), .p1m1_l(p1_l[15]), 
        .p2m1_l(p2_l[15]) );
  mul_ppgen3_192 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .p2_l(p2_l[15]), .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[14]), .p1m1_l(p1_l[14]), 
        .p2m1_l(p2_l[14]) );
  mul_ppgen3_191 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .p2_l(p2_l[14]), .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[13]), .p1m1_l(p1_l[13]), 
        .p2m1_l(p2_l[13]) );
  mul_ppgen3_190 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .p2_l(p2_l[13]), .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[12]), .p1m1_l(p1_l[12]), 
        .p2m1_l(p2_l[12]) );
  mul_ppgen3_189 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .p2_l(p2_l[12]), .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[11]), .p1m1_l(p1_l[11]), 
        .p2m1_l(p2_l[11]) );
  mul_ppgen3_188 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .p2_l(p2_l[11]), .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[10]), .p1m1_l(p1_l[10]), 
        .p2m1_l(p2_l[10]) );
  mul_ppgen3_187 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .p2_l(p2_l[10]), .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[9]), .p1m1_l(p1_l[9]), 
        .p2m1_l(p2_l[9]) );
  mul_ppgen3_186 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), 
        .p2_l(p2_l[9]), .sum(sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), .p2m1_l(p2_l[8]) );
  mul_ppgen3_185 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), 
        .p2_l(p2_l[8]), .sum(sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), .p2m1_l(p2_l[7]) );
  mul_ppgen3_184 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), 
        .p2_l(p2_l[7]), .sum(sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), .p2m1_l(p2_l[6]) );
  mul_ppgen3_183 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), 
        .p2_l(p2_l[6]), .sum(sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), .p2m1_l(p2_l[5]) );
  mul_ppgen3_182 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), 
        .p2_l(p2_l[5]), .sum(sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), .p2m1_l(p2_l[4]) );
  mul_ppgen3_181 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), 
        .p2_l(p2_l[4]), .sum(sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), .p2m1_l(1'b1) );
  mul_ppgen3lsb4_4 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ppgen_955 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_956 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_957 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_958 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_959 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_960 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_10 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_csa32_327 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_328 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_329 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  OR2X1_RVT U1 ( .A1(a), .A2(c), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(a), .A2(c), .Y(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(cout), .Y(sum) );
endmodule


module mul_csa32_330 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ppgensign_13 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_14 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_15 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_5 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net42, net47, p2_l_67, net073, p1_l_65, net38, net0118, p2_l_66,
         net078, p2_l_65, net8, p2_l_64, net15, p1_l_64, net43, net48, net35;

  mul_ppgensign_15 p0_64_ ( .p_l(net42), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_14 p2_68_ ( .p_l(sum[5]), .z(net073), .b(b2), .pm1_l(p2_l_67)
         );
  mul_ppgensign_13 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ha_10 sc1_68_ ( .cout(cout[4]), .sum(sum[4]), .a(1'b1), .b(net073) );
  mul_ppgen_960 p2_67_ ( .p_l(p2_l_67), .z(net078), .a(am1), .b(b2), .pm1_l(
        p2_l_66) );
  mul_ppgen_959 p2_66_ ( .p_l(p2_l_66), .z(net8), .a(am2), .b(b2), .pm1_l(
        p2_l_65) );
  mul_ppgen_958 p2_65_ ( .p_l(p2_l_65), .z(net15), .a(am3), .b(b2), .pm1_l(
        p2_l_64) );
  mul_ppgen_957 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_956 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_ppgen_955 p2_64_ ( .p_l(p2_l_64), .z(net35), .a(am4), .b(b2), .pm1_l(
        p2m1_l) );
  mul_csa32_330 sc1_67_ ( .sum(sum[3]), .cout(cout[3]), .a(net0118), .b(1'b0), 
        .c(net078) );
  mul_csa32_329 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(1'b1), 
        .c(net8) );
  mul_csa32_328 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net15) );
  mul_csa32_327 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net35) );
endmodule


module mul_ppgen_769 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_770 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_771 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_772 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_773 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_774 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_9 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_9 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_10 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_265 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_266 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_5 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_10 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_9 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_266 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_265 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_9 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_774 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_773 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_772 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(
        p0_l_1) );
  mul_ppgen_771 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(
        p0_l_0) );
  mul_ppgen_770 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_769 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_775 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_776 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_777 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_csa32_267 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_241 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043, net210200;

  mul_csa32_267 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_777 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(net210200) );
  mul_ppgen_776 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_775 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_778 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_779 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_780 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_268 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_242 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_268 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_780 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_779 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_778 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_781 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_782 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_783 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_269 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_243 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_269 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_783 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_782 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_781 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_784 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_785 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_786 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_270 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_244 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_270 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_786 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_785 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_784 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_787 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_788 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_789 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_271 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_245 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_271 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_789 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_788 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_787 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_790 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_791 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_792 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_272 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_246 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_272 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_792 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_791 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_790 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_793 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_794 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_795 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_273 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_247 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_273 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_795 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_794 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_793 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_796 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_797 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_798 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_274 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_248 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_274 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_798 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_797 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_796 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_799 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_800 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_801 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_275 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_249 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_275 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_801 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_800 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_799 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_802 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_803 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_804 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_276 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_250 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_276 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_804 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_803 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_802 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_805 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_806 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_807 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_277 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_251 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_277 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_807 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_806 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_805 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_808 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_809 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_810 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_278 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_252 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_278 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_810 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_809 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_808 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_811 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_812 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_813 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_279 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_253 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_279 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_813 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_812 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_811 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_814 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_815 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_816 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_280 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_254 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_280 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_816 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_815 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_814 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_817 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_818 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_819 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_281 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_255 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_281 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_819 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_818 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_817 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_820 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_821 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_822 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_282 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_256 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_282 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_822 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_821 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_820 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_823 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_824 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_825 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_283 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_257 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_283 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_825 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_824 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_823 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_826 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_827 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_828 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_284 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_258 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_284 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_828 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_827 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_826 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_829 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_830 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_831 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_285 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_259 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_285 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_831 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_830 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_829 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_832 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_833 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_834 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_286 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_260 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_286 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_834 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_833 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_832 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_835 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_836 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_837 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_287 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_261 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_287 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_837 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_836 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_835 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_838 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_839 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_840 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_288 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_262 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_288 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_840 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_839 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_838 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_841 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_842 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_843 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_289 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_263 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_289 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_843 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_842 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_841 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_844 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_845 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_846 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_290 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_264 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_290 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_846 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_845 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_844 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_847 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_848 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_849 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_291 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_265 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_291 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_849 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_848 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_847 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_850 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_851 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_852 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_292 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_266 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_292 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_852 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_851 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_850 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_853 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_854 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_855 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_293 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_267 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_293 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_855 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_854 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_853 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_856 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_857 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_858 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_294 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_268 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_294 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_858 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_857 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_856 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_859 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_860 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_861 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_295 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_269 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_295 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_861 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_860 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_859 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_862 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_863 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_864 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_296 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_270 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_296 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_864 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_863 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_862 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_865 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_866 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_867 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_297 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_271 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_297 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_867 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_866 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_865 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_868 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_869 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_870 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_298 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_272 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_298 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_870 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_869 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_868 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_871 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_872 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_873 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_299 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_273 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_299 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_873 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_872 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_871 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_874 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_875 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_876 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_300 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_274 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_300 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_876 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_875 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_874 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_877 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_878 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_879 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_301 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_275 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_301 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_879 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_878 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_877 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_880 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_881 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_882 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_302 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_276 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_302 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_882 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_881 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_880 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_883 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_884 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_885 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_303 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_277 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_303 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_885 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_884 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_883 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_886 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_887 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_888 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_304 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_278 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_304 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_888 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_887 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_886 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_889 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_890 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_891 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_305 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_279 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_305 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_891 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_890 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_889 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_892 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_893 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_894 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_306 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_280 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_306 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_894 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_893 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_892 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_895 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_896 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_897 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_307 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_281 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_307 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_897 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_896 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_895 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_898 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_899 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_900 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_308 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_282 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_308 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_900 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_899 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_898 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_901 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_902 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_903 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_309 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_283 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_309 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_903 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_902 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_901 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_904 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_905 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_906 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_310 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_284 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_310 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_906 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_905 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_904 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_907 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_908 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_909 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_311 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_285 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_311 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_909 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_908 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_907 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_910 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_911 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_912 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_312 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_286 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_312 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_912 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_911 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_910 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_913 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_914 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_915 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_313 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_287 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_313 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_915 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_914 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_913 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_916 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_917 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_918 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_314 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_288 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_314 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_918 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_917 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_916 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_919 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_920 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_921 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_315 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_289 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_315 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_921 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_920 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_919 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_922 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_923 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_924 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_316 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_290 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_316 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_924 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_923 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_922 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_925 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_926 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_927 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_317 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_291 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_317 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_927 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_926 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_925 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_928 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_929 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_930 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_318 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_292 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_318 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_930 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_929 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_928 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_931 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_932 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_933 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_319 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_293 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_319 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_933 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_932 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_931 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_934 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_935 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_936 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_320 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_294 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_320 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_936 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_935 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_934 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_937 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_938 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_939 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_321 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_295 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_321 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_939 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_938 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_937 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_940 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_941 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_942 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_322 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_296 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_322 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_942 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_941 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_940 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_943 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_944 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_945 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_323 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_297 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_323 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_945 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_944 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_943 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_946 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_947 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_948 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_324 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_298 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_324 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_948 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_947 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_946 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_949 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_950 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_951 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_325 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_299 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_325 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_951 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_950 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_949 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_952 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_953 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_954 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_326 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_300 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_326 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_954 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_953 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_952 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_5 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210277, net210278;
  wire   [63:4] p2_l;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;

  mul_ppgen3sign_5 I2 ( .cout(cout[68:64]), .sum(sum[69:64]), .am1(a[63]), 
        .am2(a[62]), .am3(a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2(b2), 
        .bot(net210277), .head(net210278), .p0m1_l(p0_l[63]), .p1m1_l(p1_l[63]), .p2m1_l(p2_l[63]) );
  mul_ppgen3_300 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .p2_l(p2_l[63]), .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[62]), .p1m1_l(p1_l[62]), 
        .p2m1_l(p2_l[62]) );
  mul_ppgen3_299 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .p2_l(p2_l[62]), .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[61]), .p1m1_l(p1_l[61]), 
        .p2m1_l(p2_l[61]) );
  mul_ppgen3_298 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .p2_l(p2_l[61]), .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[60]), .p1m1_l(p1_l[60]), 
        .p2m1_l(p2_l[60]) );
  mul_ppgen3_297 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .p2_l(p2_l[60]), .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[59]), .p1m1_l(p1_l[59]), 
        .p2m1_l(p2_l[59]) );
  mul_ppgen3_296 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .p2_l(p2_l[59]), .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[58]), .p1m1_l(p1_l[58]), 
        .p2m1_l(p2_l[58]) );
  mul_ppgen3_295 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .p2_l(p2_l[58]), .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[57]), .p1m1_l(p1_l[57]), 
        .p2m1_l(p2_l[57]) );
  mul_ppgen3_294 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .p2_l(p2_l[57]), .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[56]), .p1m1_l(p1_l[56]), 
        .p2m1_l(p2_l[56]) );
  mul_ppgen3_293 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .p2_l(p2_l[56]), .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[55]), .p1m1_l(p1_l[55]), 
        .p2m1_l(p2_l[55]) );
  mul_ppgen3_292 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .p2_l(p2_l[55]), .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[54]), .p1m1_l(p1_l[54]), 
        .p2m1_l(p2_l[54]) );
  mul_ppgen3_291 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .p2_l(p2_l[54]), .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[53]), .p1m1_l(p1_l[53]), 
        .p2m1_l(p2_l[53]) );
  mul_ppgen3_290 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .p2_l(p2_l[53]), .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[52]), .p1m1_l(p1_l[52]), 
        .p2m1_l(p2_l[52]) );
  mul_ppgen3_289 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .p2_l(p2_l[52]), .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[51]), .p1m1_l(p1_l[51]), 
        .p2m1_l(p2_l[51]) );
  mul_ppgen3_288 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .p2_l(p2_l[51]), .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[50]), .p1m1_l(p1_l[50]), 
        .p2m1_l(p2_l[50]) );
  mul_ppgen3_287 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .p2_l(p2_l[50]), .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[49]), .p1m1_l(p1_l[49]), 
        .p2m1_l(p2_l[49]) );
  mul_ppgen3_286 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .p2_l(p2_l[49]), .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[48]), .p1m1_l(p1_l[48]), 
        .p2m1_l(p2_l[48]) );
  mul_ppgen3_285 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .p2_l(p2_l[48]), .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[47]), .p1m1_l(p1_l[47]), 
        .p2m1_l(p2_l[47]) );
  mul_ppgen3_284 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .p2_l(p2_l[47]), .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[46]), .p1m1_l(p1_l[46]), 
        .p2m1_l(p2_l[46]) );
  mul_ppgen3_283 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .p2_l(p2_l[46]), .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[45]), .p1m1_l(p1_l[45]), 
        .p2m1_l(p2_l[45]) );
  mul_ppgen3_282 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .p2_l(p2_l[45]), .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[44]), .p1m1_l(p1_l[44]), 
        .p2m1_l(p2_l[44]) );
  mul_ppgen3_281 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .p2_l(p2_l[44]), .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[43]), .p1m1_l(p1_l[43]), 
        .p2m1_l(p2_l[43]) );
  mul_ppgen3_280 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .p2_l(p2_l[43]), .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[42]), .p1m1_l(p1_l[42]), 
        .p2m1_l(p2_l[42]) );
  mul_ppgen3_279 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .p2_l(p2_l[42]), .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[41]), .p1m1_l(p1_l[41]), 
        .p2m1_l(p2_l[41]) );
  mul_ppgen3_278 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .p2_l(p2_l[41]), .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[40]), .p1m1_l(p1_l[40]), 
        .p2m1_l(p2_l[40]) );
  mul_ppgen3_277 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .p2_l(p2_l[40]), .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[39]), .p1m1_l(p1_l[39]), 
        .p2m1_l(p2_l[39]) );
  mul_ppgen3_276 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .p2_l(p2_l[39]), .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[38]), .p1m1_l(p1_l[38]), 
        .p2m1_l(p2_l[38]) );
  mul_ppgen3_275 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .p2_l(p2_l[38]), .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[37]), .p1m1_l(p1_l[37]), 
        .p2m1_l(p2_l[37]) );
  mul_ppgen3_274 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .p2_l(p2_l[37]), .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[36]), .p1m1_l(p1_l[36]), 
        .p2m1_l(p2_l[36]) );
  mul_ppgen3_273 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .p2_l(p2_l[36]), .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[35]), .p1m1_l(p1_l[35]), 
        .p2m1_l(p2_l[35]) );
  mul_ppgen3_272 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .p2_l(p2_l[35]), .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[34]), .p1m1_l(p1_l[34]), 
        .p2m1_l(p2_l[34]) );
  mul_ppgen3_271 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .p2_l(p2_l[34]), .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[33]), .p1m1_l(p1_l[33]), 
        .p2m1_l(p2_l[33]) );
  mul_ppgen3_270 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .p2_l(p2_l[33]), .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[32]), .p1m1_l(p1_l[32]), 
        .p2m1_l(p2_l[32]) );
  mul_ppgen3_269 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .p2_l(p2_l[32]), .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[31]), .p1m1_l(p1_l[31]), 
        .p2m1_l(p2_l[31]) );
  mul_ppgen3_268 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .p2_l(p2_l[31]), .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[30]), .p1m1_l(p1_l[30]), 
        .p2m1_l(p2_l[30]) );
  mul_ppgen3_267 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .p2_l(p2_l[30]), .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[29]), .p1m1_l(p1_l[29]), 
        .p2m1_l(p2_l[29]) );
  mul_ppgen3_266 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .p2_l(p2_l[29]), .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[28]), .p1m1_l(p1_l[28]), 
        .p2m1_l(p2_l[28]) );
  mul_ppgen3_265 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .p2_l(p2_l[28]), .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[27]), .p1m1_l(p1_l[27]), 
        .p2m1_l(p2_l[27]) );
  mul_ppgen3_264 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .p2_l(p2_l[27]), .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[26]), .p1m1_l(p1_l[26]), 
        .p2m1_l(p2_l[26]) );
  mul_ppgen3_263 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .p2_l(p2_l[26]), .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[25]), .p1m1_l(p1_l[25]), 
        .p2m1_l(p2_l[25]) );
  mul_ppgen3_262 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .p2_l(p2_l[25]), .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[24]), .p1m1_l(p1_l[24]), 
        .p2m1_l(p2_l[24]) );
  mul_ppgen3_261 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .p2_l(p2_l[24]), .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[23]), .p1m1_l(p1_l[23]), 
        .p2m1_l(p2_l[23]) );
  mul_ppgen3_260 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .p2_l(p2_l[23]), .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[22]), .p1m1_l(p1_l[22]), 
        .p2m1_l(p2_l[22]) );
  mul_ppgen3_259 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .p2_l(p2_l[22]), .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[21]), .p1m1_l(p1_l[21]), 
        .p2m1_l(p2_l[21]) );
  mul_ppgen3_258 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .p2_l(p2_l[21]), .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[20]), .p1m1_l(p1_l[20]), 
        .p2m1_l(p2_l[20]) );
  mul_ppgen3_257 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .p2_l(p2_l[20]), .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[19]), .p1m1_l(p1_l[19]), 
        .p2m1_l(p2_l[19]) );
  mul_ppgen3_256 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .p2_l(p2_l[19]), .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[18]), .p1m1_l(p1_l[18]), 
        .p2m1_l(p2_l[18]) );
  mul_ppgen3_255 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .p2_l(p2_l[18]), .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[17]), .p1m1_l(p1_l[17]), 
        .p2m1_l(p2_l[17]) );
  mul_ppgen3_254 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .p2_l(p2_l[17]), .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[16]), .p1m1_l(p1_l[16]), 
        .p2m1_l(p2_l[16]) );
  mul_ppgen3_253 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .p2_l(p2_l[16]), .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[15]), .p1m1_l(p1_l[15]), 
        .p2m1_l(p2_l[15]) );
  mul_ppgen3_252 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .p2_l(p2_l[15]), .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[14]), .p1m1_l(p1_l[14]), 
        .p2m1_l(p2_l[14]) );
  mul_ppgen3_251 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .p2_l(p2_l[14]), .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[13]), .p1m1_l(p1_l[13]), 
        .p2m1_l(p2_l[13]) );
  mul_ppgen3_250 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .p2_l(p2_l[13]), .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[12]), .p1m1_l(p1_l[12]), 
        .p2m1_l(p2_l[12]) );
  mul_ppgen3_249 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .p2_l(p2_l[12]), .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[11]), .p1m1_l(p1_l[11]), 
        .p2m1_l(p2_l[11]) );
  mul_ppgen3_248 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .p2_l(p2_l[11]), .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[10]), .p1m1_l(p1_l[10]), 
        .p2m1_l(p2_l[10]) );
  mul_ppgen3_247 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .p2_l(p2_l[10]), .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[9]), .p1m1_l(p1_l[9]), 
        .p2m1_l(p2_l[9]) );
  mul_ppgen3_246 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), 
        .p2_l(p2_l[9]), .sum(sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), .p2m1_l(p2_l[8]) );
  mul_ppgen3_245 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), 
        .p2_l(p2_l[8]), .sum(sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), .p2m1_l(p2_l[7]) );
  mul_ppgen3_244 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), 
        .p2_l(p2_l[7]), .sum(sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), .p2m1_l(p2_l[6]) );
  mul_ppgen3_243 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), 
        .p2_l(p2_l[6]), .sum(sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), .p2m1_l(p2_l[5]) );
  mul_ppgen3_242 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), 
        .p2_l(p2_l[5]), .sum(sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), .p2m1_l(p2_l[4]) );
  mul_ppgen3_241 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), 
        .p2_l(p2_l[4]), .sum(sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), .p2m1_l(1'b1) );
  mul_ppgen3lsb4_5 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ha_62 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_63 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_64 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_65 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_66 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_ha_67 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_68 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_71 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_72 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_73 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_74 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_15 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_795 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_796 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_797 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_798 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_799 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_800 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_801 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_802 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_803 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_804 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_805 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_806 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_807 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_808 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_809 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_810 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_811 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_812 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_813 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_814 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_815 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_816 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_817 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_818 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_819 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_820 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_821 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_822 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_823 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_824 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_825 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_826 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_827 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_828 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_829 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_830 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_831 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_832 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_833 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_834 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_835 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_836 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_837 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_838 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_839 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_840 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_841 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_842 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_843 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_844 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_845 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_846 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_847 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_848 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_849 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_850 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_851 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_852 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_853 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_854 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_855 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_856 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_857 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_858 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_859 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_860 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_861 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_862 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_863 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_864 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_865 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_866 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_867 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  OR2X1_RVT U1 ( .A1(b), .A2(a), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(cout), .Y(sum) );
endmodule


module mul_csa32_868 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_869 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_870 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_871 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_872 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_873 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_874 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_875 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_876 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_877 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_878 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_879 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_880 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_881 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_882 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_883 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_884 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_885 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_886 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_887 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_888 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_889 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_890 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_891 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_892 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_893 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_894 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_895 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_896 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_897 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_898 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_899 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_900 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_901 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_902 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_903 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_904 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_905 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_906 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_907 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_908 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_909 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_910 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_911 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_912 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_913 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_914 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_915 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_916 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_917 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_918 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_919 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_920 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_921 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_922 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_923 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_924 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_925 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_926 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_927 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa42_116 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(n1), .Y(carry) );
  NAND2X0_RVT U2 ( .A1(n2), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(n2), .A2(b), .A3(n1), .Y(sum) );
  FADDX1_RVT U4 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n2) );
endmodule


module mul_csa42_117 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_118 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_119 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_120 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_121 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_122 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_123 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_124 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_125 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_126 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_127 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_128 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_129 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_130 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_131 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_132 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_133 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_134 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_135 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_136 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_137 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_138 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_139 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_140 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_141 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_142 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_143 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_144 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_145 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_146 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_147 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_148 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_149 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_150 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_151 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_152 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_153 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_154 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_155 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_156 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_157 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_158 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_159 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_160 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_161 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_162 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_163 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_164 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_165 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_166 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_167 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_168 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_169 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_170 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_171 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_172 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_173 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_174 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_175 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_176 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;


  FADDX1_RVT U1 ( .A(c), .B(b), .CI(cin), .CO(carry), .S(sum) );
endmodule


module mul_csa42_177 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_178 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_179 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_180 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_array1_0 ( cout, sum, a, b0, b1, b2, b3, b4, b5, b6, b7, b8, bot, 
        head );
  output [81:4] cout;
  output [81:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input [2:0] b3;
  input [2:0] b4;
  input [2:0] b5;
  input [2:0] b6;
  input [2:0] b7;
  input [2:0] b8;
  input bot, head;
  wire   net210890, net210891, net210892, net210893;
  wire   [1:0] b5n;
  wire   [1:0] b2n;
  wire   [76:10] s_2;
  wire   [75:11] co;
  wire   [70:2] c_1;
  wire   [76:10] c_2;
  wire   [69:0] s1;
  wire   [70:4] s_1;
  wire   [68:1] c1;
  wire   [68:1] c2;
  wire   [69:0] s2;
  wire   [68:1] c0;
  wire   [69:2] s0;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  mul_negen_0 p1n ( .n0(b5n[0]), .n1(b5n[1]), .b(b5) );
  mul_negen_15 p0n ( .n0(b2n[0]), .n1(b2n[1]), .b(b2) );
  mul_csa42_0 sc3_71_ ( .sum(sum[71]), .carry(cout[71]), .cout(co[71]), .a(
        c_1[70]), .b(c_2[70]), .c(s_2[71]), .d(s1[65]), .cin(co[70]) );
  mul_csa42_180 sc3_75_ ( .sum(sum[75]), .carry(cout[75]), .cout(co[75]), .a(
        1'b0), .b(c_2[74]), .c(s_2[75]), .d(s1[69]), .cin(co[74]) );
  mul_csa42_179 sc3_74_ ( .sum(sum[74]), .carry(cout[74]), .cout(co[74]), .a(
        1'b0), .b(c_2[73]), .c(s_2[74]), .d(s1[68]), .cin(co[73]) );
  mul_csa42_178 sc3_73_ ( .sum(sum[73]), .carry(cout[73]), .cout(co[73]), .a(
        1'b0), .b(c_2[72]), .c(s_2[73]), .d(s1[67]), .cin(co[72]) );
  mul_csa42_177 sc3_72_ ( .sum(sum[72]), .carry(cout[72]), .cout(co[72]), .a(
        1'b0), .b(c_2[71]), .c(s_2[72]), .d(s1[66]), .cin(co[71]) );
  mul_csa42_176 sc3_76_ ( .sum(sum[76]), .carry(cout[76]), .a(1'b0), .b(
        c_2[75]), .c(s_2[76]), .d(1'b0), .cin(co[75]) );
  mul_csa42_175 sc3_70_ ( .sum(sum[70]), .carry(cout[70]), .cout(co[70]), .a(
        c_1[69]), .b(c_2[69]), .c(s_2[70]), .d(s_1[70]), .cin(co[69]) );
  mul_csa42_174 sc3_69_ ( .sum(sum[69]), .carry(cout[69]), .cout(co[69]), .a(
        c_1[68]), .b(c_2[68]), .c(s_2[69]), .d(s_1[69]), .cin(co[68]) );
  mul_csa42_173 sc3_68_ ( .sum(sum[68]), .carry(cout[68]), .cout(co[68]), .a(
        c_1[67]), .b(c_2[67]), .c(s_2[68]), .d(s_1[68]), .cin(co[67]) );
  mul_csa42_172 sc3_67_ ( .sum(sum[67]), .carry(cout[67]), .cout(co[67]), .a(
        c_1[66]), .b(c_2[66]), .c(s_2[67]), .d(s_1[67]), .cin(co[66]) );
  mul_csa42_171 sc3_66_ ( .sum(sum[66]), .carry(cout[66]), .cout(co[66]), .a(
        c_1[65]), .b(c_2[65]), .c(s_2[66]), .d(s_1[66]), .cin(co[65]) );
  mul_csa42_170 sc3_65_ ( .sum(sum[65]), .carry(cout[65]), .cout(co[65]), .a(
        c_1[64]), .b(c_2[64]), .c(s_2[65]), .d(s_1[65]), .cin(co[64]) );
  mul_csa42_169 sc3_64_ ( .sum(sum[64]), .carry(cout[64]), .cout(co[64]), .a(
        c_1[63]), .b(c_2[63]), .c(s_2[64]), .d(s_1[64]), .cin(co[63]) );
  mul_csa42_168 sc3_63_ ( .sum(sum[63]), .carry(cout[63]), .cout(co[63]), .a(
        c_1[62]), .b(c_2[62]), .c(s_2[63]), .d(s_1[63]), .cin(co[62]) );
  mul_csa42_167 sc3_62_ ( .sum(sum[62]), .carry(cout[62]), .cout(co[62]), .a(
        c_1[61]), .b(c_2[61]), .c(s_2[62]), .d(s_1[62]), .cin(co[61]) );
  mul_csa42_166 sc3_61_ ( .sum(sum[61]), .carry(cout[61]), .cout(co[61]), .a(
        c_1[60]), .b(c_2[60]), .c(s_2[61]), .d(s_1[61]), .cin(co[60]) );
  mul_csa42_165 sc3_60_ ( .sum(sum[60]), .carry(cout[60]), .cout(co[60]), .a(
        c_1[59]), .b(c_2[59]), .c(s_2[60]), .d(s_1[60]), .cin(co[59]) );
  mul_csa42_164 sc3_59_ ( .sum(sum[59]), .carry(cout[59]), .cout(co[59]), .a(
        c_1[58]), .b(c_2[58]), .c(s_2[59]), .d(s_1[59]), .cin(co[58]) );
  mul_csa42_163 sc3_58_ ( .sum(sum[58]), .carry(cout[58]), .cout(co[58]), .a(
        c_1[57]), .b(c_2[57]), .c(s_2[58]), .d(s_1[58]), .cin(co[57]) );
  mul_csa42_162 sc3_57_ ( .sum(sum[57]), .carry(cout[57]), .cout(co[57]), .a(
        c_1[56]), .b(c_2[56]), .c(s_2[57]), .d(s_1[57]), .cin(co[56]) );
  mul_csa42_161 sc3_56_ ( .sum(sum[56]), .carry(cout[56]), .cout(co[56]), .a(
        c_1[55]), .b(c_2[55]), .c(s_2[56]), .d(s_1[56]), .cin(co[55]) );
  mul_csa42_160 sc3_55_ ( .sum(sum[55]), .carry(cout[55]), .cout(co[55]), .a(
        c_1[54]), .b(c_2[54]), .c(s_2[55]), .d(s_1[55]), .cin(co[54]) );
  mul_csa42_159 sc3_54_ ( .sum(sum[54]), .carry(cout[54]), .cout(co[54]), .a(
        c_1[53]), .b(c_2[53]), .c(s_2[54]), .d(s_1[54]), .cin(co[53]) );
  mul_csa42_158 sc3_53_ ( .sum(sum[53]), .carry(cout[53]), .cout(co[53]), .a(
        c_1[52]), .b(c_2[52]), .c(s_2[53]), .d(s_1[53]), .cin(co[52]) );
  mul_csa42_157 sc3_52_ ( .sum(sum[52]), .carry(cout[52]), .cout(co[52]), .a(
        c_1[51]), .b(c_2[51]), .c(s_2[52]), .d(s_1[52]), .cin(co[51]) );
  mul_csa42_156 sc3_51_ ( .sum(sum[51]), .carry(cout[51]), .cout(co[51]), .a(
        c_1[50]), .b(c_2[50]), .c(s_2[51]), .d(s_1[51]), .cin(co[50]) );
  mul_csa42_155 sc3_50_ ( .sum(sum[50]), .carry(cout[50]), .cout(co[50]), .a(
        c_1[49]), .b(c_2[49]), .c(s_2[50]), .d(s_1[50]), .cin(co[49]) );
  mul_csa42_154 sc3_49_ ( .sum(sum[49]), .carry(cout[49]), .cout(co[49]), .a(
        c_1[48]), .b(c_2[48]), .c(s_2[49]), .d(s_1[49]), .cin(co[48]) );
  mul_csa42_153 sc3_48_ ( .sum(sum[48]), .carry(cout[48]), .cout(co[48]), .a(
        c_1[47]), .b(c_2[47]), .c(s_2[48]), .d(s_1[48]), .cin(co[47]) );
  mul_csa42_152 sc3_47_ ( .sum(sum[47]), .carry(cout[47]), .cout(co[47]), .a(
        c_1[46]), .b(c_2[46]), .c(s_2[47]), .d(s_1[47]), .cin(co[46]) );
  mul_csa42_151 sc3_46_ ( .sum(sum[46]), .carry(cout[46]), .cout(co[46]), .a(
        c_1[45]), .b(c_2[45]), .c(s_2[46]), .d(s_1[46]), .cin(co[45]) );
  mul_csa42_150 sc3_45_ ( .sum(sum[45]), .carry(cout[45]), .cout(co[45]), .a(
        c_1[44]), .b(c_2[44]), .c(s_2[45]), .d(s_1[45]), .cin(co[44]) );
  mul_csa42_149 sc3_44_ ( .sum(sum[44]), .carry(cout[44]), .cout(co[44]), .a(
        c_1[43]), .b(c_2[43]), .c(s_2[44]), .d(s_1[44]), .cin(co[43]) );
  mul_csa42_148 sc3_43_ ( .sum(sum[43]), .carry(cout[43]), .cout(co[43]), .a(
        c_1[42]), .b(c_2[42]), .c(s_2[43]), .d(s_1[43]), .cin(co[42]) );
  mul_csa42_147 sc3_42_ ( .sum(sum[42]), .carry(cout[42]), .cout(co[42]), .a(
        c_1[41]), .b(c_2[41]), .c(s_2[42]), .d(s_1[42]), .cin(co[41]) );
  mul_csa42_146 sc3_41_ ( .sum(sum[41]), .carry(cout[41]), .cout(co[41]), .a(
        c_1[40]), .b(c_2[40]), .c(s_2[41]), .d(s_1[41]), .cin(co[40]) );
  mul_csa42_145 sc3_40_ ( .sum(sum[40]), .carry(cout[40]), .cout(co[40]), .a(
        c_1[39]), .b(c_2[39]), .c(s_2[40]), .d(s_1[40]), .cin(co[39]) );
  mul_csa42_144 sc3_39_ ( .sum(sum[39]), .carry(cout[39]), .cout(co[39]), .a(
        c_1[38]), .b(c_2[38]), .c(s_2[39]), .d(s_1[39]), .cin(co[38]) );
  mul_csa42_143 sc3_38_ ( .sum(sum[38]), .carry(cout[38]), .cout(co[38]), .a(
        c_1[37]), .b(c_2[37]), .c(s_2[38]), .d(s_1[38]), .cin(co[37]) );
  mul_csa42_142 sc3_37_ ( .sum(sum[37]), .carry(cout[37]), .cout(co[37]), .a(
        c_1[36]), .b(c_2[36]), .c(s_2[37]), .d(s_1[37]), .cin(co[36]) );
  mul_csa42_141 sc3_36_ ( .sum(sum[36]), .carry(cout[36]), .cout(co[36]), .a(
        c_1[35]), .b(c_2[35]), .c(s_2[36]), .d(s_1[36]), .cin(co[35]) );
  mul_csa42_140 sc3_35_ ( .sum(sum[35]), .carry(cout[35]), .cout(co[35]), .a(
        c_1[34]), .b(c_2[34]), .c(s_2[35]), .d(s_1[35]), .cin(co[34]) );
  mul_csa42_139 sc3_34_ ( .sum(sum[34]), .carry(cout[34]), .cout(co[34]), .a(
        c_1[33]), .b(c_2[33]), .c(s_2[34]), .d(s_1[34]), .cin(co[33]) );
  mul_csa42_138 sc3_33_ ( .sum(sum[33]), .carry(cout[33]), .cout(co[33]), .a(
        c_1[32]), .b(c_2[32]), .c(s_2[33]), .d(s_1[33]), .cin(co[32]) );
  mul_csa42_137 sc3_32_ ( .sum(sum[32]), .carry(cout[32]), .cout(co[32]), .a(
        c_1[31]), .b(c_2[31]), .c(s_2[32]), .d(s_1[32]), .cin(co[31]) );
  mul_csa42_136 sc3_31_ ( .sum(sum[31]), .carry(cout[31]), .cout(co[31]), .a(
        c_1[30]), .b(c_2[30]), .c(s_2[31]), .d(s_1[31]), .cin(co[30]) );
  mul_csa42_135 sc3_30_ ( .sum(sum[30]), .carry(cout[30]), .cout(co[30]), .a(
        c_1[29]), .b(c_2[29]), .c(s_2[30]), .d(s_1[30]), .cin(co[29]) );
  mul_csa42_134 sc3_29_ ( .sum(sum[29]), .carry(cout[29]), .cout(co[29]), .a(
        c_1[28]), .b(c_2[28]), .c(s_2[29]), .d(s_1[29]), .cin(co[28]) );
  mul_csa42_133 sc3_28_ ( .sum(sum[28]), .carry(cout[28]), .cout(co[28]), .a(
        c_1[27]), .b(c_2[27]), .c(s_2[28]), .d(s_1[28]), .cin(co[27]) );
  mul_csa42_132 sc3_27_ ( .sum(sum[27]), .carry(cout[27]), .cout(co[27]), .a(
        c_1[26]), .b(c_2[26]), .c(s_2[27]), .d(s_1[27]), .cin(co[26]) );
  mul_csa42_131 sc3_26_ ( .sum(sum[26]), .carry(cout[26]), .cout(co[26]), .a(
        c_1[25]), .b(c_2[25]), .c(s_2[26]), .d(s_1[26]), .cin(co[25]) );
  mul_csa42_130 sc3_25_ ( .sum(sum[25]), .carry(cout[25]), .cout(co[25]), .a(
        c_1[24]), .b(c_2[24]), .c(s_2[25]), .d(s_1[25]), .cin(co[24]) );
  mul_csa42_129 sc3_24_ ( .sum(sum[24]), .carry(cout[24]), .cout(co[24]), .a(
        c_1[23]), .b(c_2[23]), .c(s_2[24]), .d(s_1[24]), .cin(co[23]) );
  mul_csa42_128 sc3_23_ ( .sum(sum[23]), .carry(cout[23]), .cout(co[23]), .a(
        c_1[22]), .b(c_2[22]), .c(s_2[23]), .d(s_1[23]), .cin(co[22]) );
  mul_csa42_127 sc3_22_ ( .sum(sum[22]), .carry(cout[22]), .cout(co[22]), .a(
        c_1[21]), .b(c_2[21]), .c(s_2[22]), .d(s_1[22]), .cin(co[21]) );
  mul_csa42_126 sc3_21_ ( .sum(sum[21]), .carry(cout[21]), .cout(co[21]), .a(
        c_1[20]), .b(c_2[20]), .c(s_2[21]), .d(s_1[21]), .cin(co[20]) );
  mul_csa42_125 sc3_20_ ( .sum(sum[20]), .carry(cout[20]), .cout(co[20]), .a(
        c_1[19]), .b(c_2[19]), .c(s_2[20]), .d(s_1[20]), .cin(co[19]) );
  mul_csa42_124 sc3_19_ ( .sum(sum[19]), .carry(cout[19]), .cout(co[19]), .a(
        c_1[18]), .b(c_2[18]), .c(s_2[19]), .d(s_1[19]), .cin(co[18]) );
  mul_csa42_123 sc3_18_ ( .sum(sum[18]), .carry(cout[18]), .cout(co[18]), .a(
        c_1[17]), .b(c_2[17]), .c(s_2[18]), .d(s_1[18]), .cin(co[17]) );
  mul_csa42_122 sc3_17_ ( .sum(sum[17]), .carry(cout[17]), .cout(co[17]), .a(
        c_1[16]), .b(c_2[16]), .c(s_2[17]), .d(s_1[17]), .cin(co[16]) );
  mul_csa42_121 sc3_16_ ( .sum(sum[16]), .carry(cout[16]), .cout(co[16]), .a(
        c_1[15]), .b(c_2[15]), .c(s_2[16]), .d(s_1[16]), .cin(co[15]) );
  mul_csa42_120 sc3_15_ ( .sum(sum[15]), .carry(cout[15]), .cout(co[15]), .a(
        c_1[14]), .b(c_2[14]), .c(s_2[15]), .d(s_1[15]), .cin(co[14]) );
  mul_csa42_119 sc3_14_ ( .sum(sum[14]), .carry(cout[14]), .cout(co[14]), .a(
        c_1[13]), .b(c_2[13]), .c(s_2[14]), .d(s_1[14]), .cin(co[13]) );
  mul_csa42_118 sc3_13_ ( .sum(sum[13]), .carry(cout[13]), .cout(co[13]), .a(
        c_1[12]), .b(c_2[12]), .c(s_2[13]), .d(s_1[13]), .cin(co[12]) );
  mul_csa42_117 sc3_12_ ( .sum(sum[12]), .carry(cout[12]), .cout(co[12]), .a(
        c_1[11]), .b(c_2[11]), .c(s_2[12]), .d(s_1[12]), .cin(co[11]) );
  mul_csa42_116 sc3_11_ ( .sum(sum[11]), .carry(cout[11]), .cout(co[11]), .a(
        c_1[10]), .b(c_2[10]), .c(s_2[11]), .d(s_1[11]), .cin(1'b0) );
  mul_csa32_0 sc2_2_70_ ( .sum(s_2[70]), .cout(c_2[70]), .a(s2[58]), .b(c2[57]), .c(c1[63]) );
  mul_csa32_927 sc2_2_69_ ( .sum(s_2[69]), .cout(c_2[69]), .a(s2[57]), .b(
        c2[56]), .c(c1[62]) );
  mul_csa32_926 sc2_2_68_ ( .sum(s_2[68]), .cout(c_2[68]), .a(s2[56]), .b(
        c2[55]), .c(c1[61]) );
  mul_csa32_925 sc2_2_67_ ( .sum(s_2[67]), .cout(c_2[67]), .a(s2[55]), .b(
        c2[54]), .c(c1[60]) );
  mul_csa32_924 sc2_2_66_ ( .sum(s_2[66]), .cout(c_2[66]), .a(s2[54]), .b(
        c2[53]), .c(c1[59]) );
  mul_csa32_923 sc2_2_65_ ( .sum(s_2[65]), .cout(c_2[65]), .a(s2[53]), .b(
        c2[52]), .c(c1[58]) );
  mul_csa32_922 sc2_2_64_ ( .sum(s_2[64]), .cout(c_2[64]), .a(s2[52]), .b(
        c2[51]), .c(c1[57]) );
  mul_csa32_921 sc2_2_63_ ( .sum(s_2[63]), .cout(c_2[63]), .a(s2[51]), .b(
        c2[50]), .c(c1[56]) );
  mul_csa32_920 sc2_2_62_ ( .sum(s_2[62]), .cout(c_2[62]), .a(s2[50]), .b(
        c2[49]), .c(c1[55]) );
  mul_csa32_919 sc2_2_61_ ( .sum(s_2[61]), .cout(c_2[61]), .a(s2[49]), .b(
        c2[48]), .c(c1[54]) );
  mul_csa32_918 sc2_2_60_ ( .sum(s_2[60]), .cout(c_2[60]), .a(s2[48]), .b(
        c2[47]), .c(c1[53]) );
  mul_csa32_917 sc2_2_59_ ( .sum(s_2[59]), .cout(c_2[59]), .a(s2[47]), .b(
        c2[46]), .c(c1[52]) );
  mul_csa32_916 sc2_2_58_ ( .sum(s_2[58]), .cout(c_2[58]), .a(s2[46]), .b(
        c2[45]), .c(c1[51]) );
  mul_csa32_915 sc2_2_57_ ( .sum(s_2[57]), .cout(c_2[57]), .a(s2[45]), .b(
        c2[44]), .c(c1[50]) );
  mul_csa32_914 sc2_2_56_ ( .sum(s_2[56]), .cout(c_2[56]), .a(s2[44]), .b(
        c2[43]), .c(c1[49]) );
  mul_csa32_913 sc2_2_55_ ( .sum(s_2[55]), .cout(c_2[55]), .a(s2[43]), .b(
        c2[42]), .c(c1[48]) );
  mul_csa32_912 sc2_2_54_ ( .sum(s_2[54]), .cout(c_2[54]), .a(s2[42]), .b(
        c2[41]), .c(c1[47]) );
  mul_csa32_911 sc2_2_53_ ( .sum(s_2[53]), .cout(c_2[53]), .a(s2[41]), .b(
        c2[40]), .c(c1[46]) );
  mul_csa32_910 sc2_2_52_ ( .sum(s_2[52]), .cout(c_2[52]), .a(s2[40]), .b(
        c2[39]), .c(c1[45]) );
  mul_csa32_909 sc2_2_51_ ( .sum(s_2[51]), .cout(c_2[51]), .a(s2[39]), .b(
        c2[38]), .c(c1[44]) );
  mul_csa32_908 sc2_2_50_ ( .sum(s_2[50]), .cout(c_2[50]), .a(s2[38]), .b(
        c2[37]), .c(c1[43]) );
  mul_csa32_907 sc2_2_49_ ( .sum(s_2[49]), .cout(c_2[49]), .a(s2[37]), .b(
        c2[36]), .c(c1[42]) );
  mul_csa32_906 sc2_2_48_ ( .sum(s_2[48]), .cout(c_2[48]), .a(s2[36]), .b(
        c2[35]), .c(c1[41]) );
  mul_csa32_905 sc2_2_47_ ( .sum(s_2[47]), .cout(c_2[47]), .a(s2[35]), .b(
        c2[34]), .c(c1[40]) );
  mul_csa32_904 sc2_2_46_ ( .sum(s_2[46]), .cout(c_2[46]), .a(s2[34]), .b(
        c2[33]), .c(c1[39]) );
  mul_csa32_903 sc2_2_45_ ( .sum(s_2[45]), .cout(c_2[45]), .a(s2[33]), .b(
        c2[32]), .c(c1[38]) );
  mul_csa32_902 sc2_2_44_ ( .sum(s_2[44]), .cout(c_2[44]), .a(s2[32]), .b(
        c2[31]), .c(c1[37]) );
  mul_csa32_901 sc2_2_43_ ( .sum(s_2[43]), .cout(c_2[43]), .a(s2[31]), .b(
        c2[30]), .c(c1[36]) );
  mul_csa32_900 sc2_2_42_ ( .sum(s_2[42]), .cout(c_2[42]), .a(s2[30]), .b(
        c2[29]), .c(c1[35]) );
  mul_csa32_899 sc2_2_41_ ( .sum(s_2[41]), .cout(c_2[41]), .a(s2[29]), .b(
        c2[28]), .c(c1[34]) );
  mul_csa32_898 sc2_2_40_ ( .sum(s_2[40]), .cout(c_2[40]), .a(s2[28]), .b(
        c2[27]), .c(c1[33]) );
  mul_csa32_897 sc2_2_39_ ( .sum(s_2[39]), .cout(c_2[39]), .a(s2[27]), .b(
        c2[26]), .c(c1[32]) );
  mul_csa32_896 sc2_2_38_ ( .sum(s_2[38]), .cout(c_2[38]), .a(s2[26]), .b(
        c2[25]), .c(c1[31]) );
  mul_csa32_895 sc2_2_37_ ( .sum(s_2[37]), .cout(c_2[37]), .a(s2[25]), .b(
        c2[24]), .c(c1[30]) );
  mul_csa32_894 sc2_2_36_ ( .sum(s_2[36]), .cout(c_2[36]), .a(s2[24]), .b(
        c2[23]), .c(c1[29]) );
  mul_csa32_893 sc2_2_35_ ( .sum(s_2[35]), .cout(c_2[35]), .a(s2[23]), .b(
        c2[22]), .c(c1[28]) );
  mul_csa32_892 sc2_2_34_ ( .sum(s_2[34]), .cout(c_2[34]), .a(s2[22]), .b(
        c2[21]), .c(c1[27]) );
  mul_csa32_891 sc2_2_33_ ( .sum(s_2[33]), .cout(c_2[33]), .a(s2[21]), .b(
        c2[20]), .c(c1[26]) );
  mul_csa32_890 sc2_2_32_ ( .sum(s_2[32]), .cout(c_2[32]), .a(s2[20]), .b(
        c2[19]), .c(c1[25]) );
  mul_csa32_889 sc2_2_31_ ( .sum(s_2[31]), .cout(c_2[31]), .a(s2[19]), .b(
        c2[18]), .c(c1[24]) );
  mul_csa32_888 sc2_2_30_ ( .sum(s_2[30]), .cout(c_2[30]), .a(s2[18]), .b(
        c2[17]), .c(c1[23]) );
  mul_csa32_887 sc2_2_29_ ( .sum(s_2[29]), .cout(c_2[29]), .a(s2[17]), .b(
        c2[16]), .c(c1[22]) );
  mul_csa32_886 sc2_2_28_ ( .sum(s_2[28]), .cout(c_2[28]), .a(s2[16]), .b(
        c2[15]), .c(c1[21]) );
  mul_csa32_885 sc2_2_27_ ( .sum(s_2[27]), .cout(c_2[27]), .a(s2[15]), .b(
        c2[14]), .c(c1[20]) );
  mul_csa32_884 sc2_2_26_ ( .sum(s_2[26]), .cout(c_2[26]), .a(s2[14]), .b(
        c2[13]), .c(c1[19]) );
  mul_csa32_883 sc2_2_25_ ( .sum(s_2[25]), .cout(c_2[25]), .a(s2[13]), .b(
        c2[12]), .c(c1[18]) );
  mul_csa32_882 sc2_2_24_ ( .sum(s_2[24]), .cout(c_2[24]), .a(s2[12]), .b(
        c2[11]), .c(c1[17]) );
  mul_csa32_881 sc2_2_23_ ( .sum(s_2[23]), .cout(c_2[23]), .a(s2[11]), .b(
        c2[10]), .c(c1[16]) );
  mul_csa32_880 sc2_2_22_ ( .sum(s_2[22]), .cout(c_2[22]), .a(s2[10]), .b(
        c2[9]), .c(c1[15]) );
  mul_csa32_879 sc2_2_21_ ( .sum(s_2[21]), .cout(c_2[21]), .a(s2[9]), .b(c2[8]), .c(c1[14]) );
  mul_csa32_878 sc2_2_20_ ( .sum(s_2[20]), .cout(c_2[20]), .a(s2[8]), .b(c2[7]), .c(c1[13]) );
  mul_csa32_877 sc2_2_19_ ( .sum(s_2[19]), .cout(c_2[19]), .a(s2[7]), .b(c2[6]), .c(c1[12]) );
  mul_csa32_876 sc2_2_18_ ( .sum(s_2[18]), .cout(c_2[18]), .a(s2[6]), .b(c2[5]), .c(c1[11]) );
  mul_csa32_875 sc2_2_17_ ( .sum(s_2[17]), .cout(c_2[17]), .a(s2[5]), .b(c2[4]), .c(c1[10]) );
  mul_csa32_874 sc2_2_16_ ( .sum(s_2[16]), .cout(c_2[16]), .a(s2[4]), .b(c2[3]), .c(c1[9]) );
  mul_csa32_873 sc2_2_15_ ( .sum(s_2[15]), .cout(c_2[15]), .a(s2[3]), .b(c2[2]), .c(c1[8]) );
  mul_csa32_872 sc2_2_14_ ( .sum(s_2[14]), .cout(c_2[14]), .a(s2[2]), .b(c2[1]), .c(c1[7]) );
  mul_csa32_871 sc2_2_13_ ( .sum(s_2[13]), .cout(c_2[13]), .a(s2[1]), .b(s1[7]), .c(c1[6]) );
  mul_csa32_870 sc2_2_12_ ( .sum(s_2[12]), .cout(c_2[12]), .a(s2[0]), .b(s1[6]), .c(c1[5]) );
  mul_csa32_869 sc2_2_11_ ( .sum(s_2[11]), .cout(c_2[11]), .a(b5n[1]), .b(
        s1[5]), .c(c1[4]) );
  mul_csa32_868 sc2_2_10_ ( .sum(s_2[10]), .cout(c_2[10]), .a(b5n[0]), .b(
        s1[4]), .c(c1[3]) );
  mul_csa32_867 sc2_2_76_ ( .sum(s_2[76]), .cout(c_2[76]), .a(s2[64]), .b(
        c2[63]), .c(1'b1) );
  mul_csa32_866 sc2_2_77_ ( .sum(sum[77]), .cout(cout[77]), .a(s2[65]), .b(
        c2[64]), .c(c_2[76]) );
  mul_csa32_865 sc2_1_9_ ( .sum(s_1[9]), .cout(c_1[9]), .a(s0[9]), .b(c0[8]), 
        .c(s1[3]) );
  mul_csa32_864 sc2_1_8_ ( .sum(s_1[8]), .cout(c_1[8]), .a(s0[8]), .b(c0[7]), 
        .c(s1[2]) );
  mul_csa32_863 sc2_1_3_ ( .sum(sum[3]), .cout(c_1[3]), .a(s0[3]), .b(c0[2]), 
        .c(c_1[2]) );
  mul_csa32_862 sc3_10_ ( .sum(sum[10]), .cout(cout[10]), .a(c_1[9]), .b(
        s_1[10]), .c(s_2[10]) );
  mul_csa32_861 sc3_9_ ( .sum(sum[9]), .cout(cout[9]), .a(c_1[8]), .b(s_1[9]), 
        .c(c1[2]) );
  mul_csa32_860 sc3_8_ ( .sum(sum[8]), .cout(cout[8]), .a(c_1[7]), .b(s_1[8]), 
        .c(c1[1]) );
  mul_csa32_859 sc2_2_71_ ( .sum(s_2[71]), .cout(c_2[71]), .a(s2[59]), .b(
        c2[58]), .c(c1[64]) );
  mul_csa32_858 sc2_2_75_ ( .sum(s_2[75]), .cout(c_2[75]), .a(s2[63]), .b(
        c2[62]), .c(c1[68]) );
  mul_csa32_857 sc2_2_74_ ( .sum(s_2[74]), .cout(c_2[74]), .a(s2[62]), .b(
        c2[61]), .c(c1[67]) );
  mul_csa32_856 sc2_2_73_ ( .sum(s_2[73]), .cout(c_2[73]), .a(s2[61]), .b(
        c2[60]), .c(c1[66]) );
  mul_csa32_855 sc2_2_72_ ( .sum(s_2[72]), .cout(c_2[72]), .a(s2[60]), .b(
        c2[59]), .c(c1[65]) );
  mul_csa32_854 sc2_1_69_ ( .sum(s_1[69]), .cout(c_1[69]), .a(s0[69]), .b(
        c0[68]), .c(s1[63]) );
  mul_csa32_853 sc2_1_68_ ( .sum(s_1[68]), .cout(c_1[68]), .a(s0[68]), .b(
        c0[67]), .c(s1[62]) );
  mul_csa32_852 sc2_1_67_ ( .sum(s_1[67]), .cout(c_1[67]), .a(s0[67]), .b(
        c0[66]), .c(s1[61]) );
  mul_csa32_851 sc2_1_66_ ( .sum(s_1[66]), .cout(c_1[66]), .a(s0[66]), .b(
        c0[65]), .c(s1[60]) );
  mul_csa32_850 sc2_1_65_ ( .sum(s_1[65]), .cout(c_1[65]), .a(s0[65]), .b(
        c0[64]), .c(s1[59]) );
  mul_csa32_849 sc2_1_64_ ( .sum(s_1[64]), .cout(c_1[64]), .a(s0[64]), .b(
        c0[63]), .c(s1[58]) );
  mul_csa32_848 sc2_1_63_ ( .sum(s_1[63]), .cout(c_1[63]), .a(s0[63]), .b(
        c0[62]), .c(s1[57]) );
  mul_csa32_847 sc2_1_62_ ( .sum(s_1[62]), .cout(c_1[62]), .a(s0[62]), .b(
        c0[61]), .c(s1[56]) );
  mul_csa32_846 sc2_1_61_ ( .sum(s_1[61]), .cout(c_1[61]), .a(s0[61]), .b(
        c0[60]), .c(s1[55]) );
  mul_csa32_845 sc2_1_60_ ( .sum(s_1[60]), .cout(c_1[60]), .a(s0[60]), .b(
        c0[59]), .c(s1[54]) );
  mul_csa32_844 sc2_1_59_ ( .sum(s_1[59]), .cout(c_1[59]), .a(s0[59]), .b(
        c0[58]), .c(s1[53]) );
  mul_csa32_843 sc2_1_58_ ( .sum(s_1[58]), .cout(c_1[58]), .a(s0[58]), .b(
        c0[57]), .c(s1[52]) );
  mul_csa32_842 sc2_1_57_ ( .sum(s_1[57]), .cout(c_1[57]), .a(s0[57]), .b(
        c0[56]), .c(s1[51]) );
  mul_csa32_841 sc2_1_56_ ( .sum(s_1[56]), .cout(c_1[56]), .a(s0[56]), .b(
        c0[55]), .c(s1[50]) );
  mul_csa32_840 sc2_1_55_ ( .sum(s_1[55]), .cout(c_1[55]), .a(s0[55]), .b(
        c0[54]), .c(s1[49]) );
  mul_csa32_839 sc2_1_54_ ( .sum(s_1[54]), .cout(c_1[54]), .a(s0[54]), .b(
        c0[53]), .c(s1[48]) );
  mul_csa32_838 sc2_1_53_ ( .sum(s_1[53]), .cout(c_1[53]), .a(s0[53]), .b(
        c0[52]), .c(s1[47]) );
  mul_csa32_837 sc2_1_52_ ( .sum(s_1[52]), .cout(c_1[52]), .a(s0[52]), .b(
        c0[51]), .c(s1[46]) );
  mul_csa32_836 sc2_1_51_ ( .sum(s_1[51]), .cout(c_1[51]), .a(s0[51]), .b(
        c0[50]), .c(s1[45]) );
  mul_csa32_835 sc2_1_50_ ( .sum(s_1[50]), .cout(c_1[50]), .a(s0[50]), .b(
        c0[49]), .c(s1[44]) );
  mul_csa32_834 sc2_1_49_ ( .sum(s_1[49]), .cout(c_1[49]), .a(s0[49]), .b(
        c0[48]), .c(s1[43]) );
  mul_csa32_833 sc2_1_48_ ( .sum(s_1[48]), .cout(c_1[48]), .a(s0[48]), .b(
        c0[47]), .c(s1[42]) );
  mul_csa32_832 sc2_1_47_ ( .sum(s_1[47]), .cout(c_1[47]), .a(s0[47]), .b(
        c0[46]), .c(s1[41]) );
  mul_csa32_831 sc2_1_46_ ( .sum(s_1[46]), .cout(c_1[46]), .a(s0[46]), .b(
        c0[45]), .c(s1[40]) );
  mul_csa32_830 sc2_1_45_ ( .sum(s_1[45]), .cout(c_1[45]), .a(s0[45]), .b(
        c0[44]), .c(s1[39]) );
  mul_csa32_829 sc2_1_44_ ( .sum(s_1[44]), .cout(c_1[44]), .a(s0[44]), .b(
        c0[43]), .c(s1[38]) );
  mul_csa32_828 sc2_1_43_ ( .sum(s_1[43]), .cout(c_1[43]), .a(s0[43]), .b(
        c0[42]), .c(s1[37]) );
  mul_csa32_827 sc2_1_42_ ( .sum(s_1[42]), .cout(c_1[42]), .a(s0[42]), .b(
        c0[41]), .c(s1[36]) );
  mul_csa32_826 sc2_1_41_ ( .sum(s_1[41]), .cout(c_1[41]), .a(s0[41]), .b(
        c0[40]), .c(s1[35]) );
  mul_csa32_825 sc2_1_40_ ( .sum(s_1[40]), .cout(c_1[40]), .a(s0[40]), .b(
        c0[39]), .c(s1[34]) );
  mul_csa32_824 sc2_1_39_ ( .sum(s_1[39]), .cout(c_1[39]), .a(s0[39]), .b(
        c0[38]), .c(s1[33]) );
  mul_csa32_823 sc2_1_38_ ( .sum(s_1[38]), .cout(c_1[38]), .a(s0[38]), .b(
        c0[37]), .c(s1[32]) );
  mul_csa32_822 sc2_1_37_ ( .sum(s_1[37]), .cout(c_1[37]), .a(s0[37]), .b(
        c0[36]), .c(s1[31]) );
  mul_csa32_821 sc2_1_36_ ( .sum(s_1[36]), .cout(c_1[36]), .a(s0[36]), .b(
        c0[35]), .c(s1[30]) );
  mul_csa32_820 sc2_1_35_ ( .sum(s_1[35]), .cout(c_1[35]), .a(s0[35]), .b(
        c0[34]), .c(s1[29]) );
  mul_csa32_819 sc2_1_34_ ( .sum(s_1[34]), .cout(c_1[34]), .a(s0[34]), .b(
        c0[33]), .c(s1[28]) );
  mul_csa32_818 sc2_1_33_ ( .sum(s_1[33]), .cout(c_1[33]), .a(s0[33]), .b(
        c0[32]), .c(s1[27]) );
  mul_csa32_817 sc2_1_32_ ( .sum(s_1[32]), .cout(c_1[32]), .a(s0[32]), .b(
        c0[31]), .c(s1[26]) );
  mul_csa32_816 sc2_1_31_ ( .sum(s_1[31]), .cout(c_1[31]), .a(s0[31]), .b(
        c0[30]), .c(s1[25]) );
  mul_csa32_815 sc2_1_30_ ( .sum(s_1[30]), .cout(c_1[30]), .a(s0[30]), .b(
        c0[29]), .c(s1[24]) );
  mul_csa32_814 sc2_1_29_ ( .sum(s_1[29]), .cout(c_1[29]), .a(s0[29]), .b(
        c0[28]), .c(s1[23]) );
  mul_csa32_813 sc2_1_28_ ( .sum(s_1[28]), .cout(c_1[28]), .a(s0[28]), .b(
        c0[27]), .c(s1[22]) );
  mul_csa32_812 sc2_1_27_ ( .sum(s_1[27]), .cout(c_1[27]), .a(s0[27]), .b(
        c0[26]), .c(s1[21]) );
  mul_csa32_811 sc2_1_26_ ( .sum(s_1[26]), .cout(c_1[26]), .a(s0[26]), .b(
        c0[25]), .c(s1[20]) );
  mul_csa32_810 sc2_1_25_ ( .sum(s_1[25]), .cout(c_1[25]), .a(s0[25]), .b(
        c0[24]), .c(s1[19]) );
  mul_csa32_809 sc2_1_24_ ( .sum(s_1[24]), .cout(c_1[24]), .a(s0[24]), .b(
        c0[23]), .c(s1[18]) );
  mul_csa32_808 sc2_1_23_ ( .sum(s_1[23]), .cout(c_1[23]), .a(s0[23]), .b(
        c0[22]), .c(s1[17]) );
  mul_csa32_807 sc2_1_22_ ( .sum(s_1[22]), .cout(c_1[22]), .a(s0[22]), .b(
        c0[21]), .c(s1[16]) );
  mul_csa32_806 sc2_1_21_ ( .sum(s_1[21]), .cout(c_1[21]), .a(s0[21]), .b(
        c0[20]), .c(s1[15]) );
  mul_csa32_805 sc2_1_20_ ( .sum(s_1[20]), .cout(c_1[20]), .a(s0[20]), .b(
        c0[19]), .c(s1[14]) );
  mul_csa32_804 sc2_1_19_ ( .sum(s_1[19]), .cout(c_1[19]), .a(s0[19]), .b(
        c0[18]), .c(s1[13]) );
  mul_csa32_803 sc2_1_18_ ( .sum(s_1[18]), .cout(c_1[18]), .a(s0[18]), .b(
        c0[17]), .c(s1[12]) );
  mul_csa32_802 sc2_1_17_ ( .sum(s_1[17]), .cout(c_1[17]), .a(s0[17]), .b(
        c0[16]), .c(s1[11]) );
  mul_csa32_801 sc2_1_16_ ( .sum(s_1[16]), .cout(c_1[16]), .a(s0[16]), .b(
        c0[15]), .c(s1[10]) );
  mul_csa32_800 sc2_1_15_ ( .sum(s_1[15]), .cout(c_1[15]), .a(s0[15]), .b(
        c0[14]), .c(s1[9]) );
  mul_csa32_799 sc2_1_14_ ( .sum(s_1[14]), .cout(c_1[14]), .a(s0[14]), .b(
        c0[13]), .c(s1[8]) );
  mul_csa32_798 sc2_1_7_ ( .sum(s_1[7]), .cout(c_1[7]), .a(s0[7]), .b(c0[6]), 
        .c(s1[1]) );
  mul_csa32_797 sc2_1_6_ ( .sum(s_1[6]), .cout(c_1[6]), .a(s0[6]), .b(c0[5]), 
        .c(s1[0]) );
  mul_csa32_796 sc2_1_5_ ( .sum(s_1[5]), .cout(c_1[5]), .a(s0[5]), .b(c0[4]), 
        .c(b2n[1]) );
  mul_csa32_795 sc2_1_4_ ( .sum(s_1[4]), .cout(c_1[4]), .a(s0[4]), .b(c0[3]), 
        .c(b2n[0]) );
  mul_ha_0 sc2_1_10_ ( .cout(c_1[10]), .sum(s_1[10]), .a(s0[10]), .b(c0[9]) );
  mul_ha_74 sc3_7_ ( .cout(cout[7]), .sum(sum[7]), .a(c_1[6]), .b(s_1[7]) );
  mul_ha_73 sc3_6_ ( .cout(cout[6]), .sum(sum[6]), .a(c_1[5]), .b(s_1[6]) );
  mul_ha_72 sc3_5_ ( .cout(cout[5]), .sum(sum[5]), .a(c_1[4]), .b(s_1[5]) );
  mul_ha_71 sc3_4_ ( .cout(cout[4]), .sum(sum[4]), .a(c_1[3]), .b(s_1[4]) );
  mul_ha_68 sc2_2_79_ ( .cout(cout[79]), .sum(sum[79]), .a(s2[67]), .b(c2[66])
         );
  mul_ha_67 sc2_2_78_ ( .cout(cout[78]), .sum(sum[78]), .a(s2[66]), .b(c2[65])
         );
  mul_ha_66 sc2_1_70_ ( .cout(c_1[70]), .sum(s_1[70]), .a(1'b1), .b(s1[64]) );
  mul_ha_65 sc2_1_2_ ( .cout(c_1[2]), .sum(sum[2]), .a(s0[2]), .b(c0[1]) );
  mul_ha_64 sc2_1_13_ ( .cout(c_1[13]), .sum(s_1[13]), .a(s0[13]), .b(c0[12])
         );
  mul_ha_63 sc2_1_12_ ( .cout(c_1[12]), .sum(s_1[12]), .a(s0[12]), .b(c0[11])
         );
  mul_ha_62 sc2_1_11_ ( .cout(c_1[11]), .sum(s_1[11]), .a(s0[11]), .b(c0[10])
         );
  mul_ppgenrow3_0 I2 ( .cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        c2[66:1]}), .sum({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        s2[67:0]}), .a(a), .b0(b6), .b1(b7), .b2({net210890, net210891, 
        net210892}), .bot(net210893), .head(1'b0) );
  mul_ppgenrow3_5 I1 ( .cout(c1), .sum(s1), .a(a), .b0(b3), .b1(b4), .b2(b5), 
        .bot(1'b1), .head(1'b0) );
  mul_ppgenrow3_4 I0 ( .cout(c0), .sum({s0, sum[1:0]}), .a(a), .b0(b0), .b1(b1), .b2(b2), .bot(1'b1), .head(head) );
endmodule


module mul_ha_14 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   a;
  assign sum = a;

endmodule


module mul_ha_15 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_16 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_17 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_18 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_20 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_21 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_22 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_23 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_24 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_25 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_26 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_27 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_28 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_29 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_30 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_31 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_32 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_33 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_34 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_35 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_36 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_37 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_38 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_39 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_40 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_41 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_42 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_43 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_44 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_45 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_47 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign sum = b;

endmodule


module mul_csa32_397 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_398 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_399 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   b;
  assign sum = b;

endmodule


module mul_csa32_400 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_401 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_402 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_403 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_404 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_405 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_406 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_407 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_408 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_409 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_410 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_411 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_412 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_413 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_414 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_415 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_416 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_417 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_418 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_419 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_420 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_421 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_422 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_423 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_424 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_425 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_426 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_427 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_428 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_429 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_430 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_431 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_432 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_433 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_434 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_435 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_436 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_437 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_438 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_439 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_440 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_441 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_442 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_443 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_444 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_445 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_446 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_447 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_448 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_449 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_450 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_451 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_452 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_453 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_454 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_455 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_456 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_457 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_458 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_459 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_460 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_461 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_462 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_463 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_464 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_465 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_466 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_467 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_468 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_469 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_470 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_471 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_472 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_473 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_474 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_475 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_476 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_477 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_478 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_479 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_480 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_481 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_482 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_483 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_484 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_485 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_486 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_487 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_488 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_489 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_490 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_491 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_492 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_493 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_494 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_495 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_496 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_497 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_498 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_499 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_500 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_501 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_502 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_503 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_504 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_505 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_506 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_507 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_508 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_509 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_510 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_511 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_512 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_513 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_514 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_515 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_516 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_517 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_518 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_519 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_520 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_521 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_522 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_523 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_524 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_525 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_526 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_527 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_528 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_529 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_530 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_531 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_532 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_533 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_534 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_535 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_536 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_537 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_538 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_539 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_540 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_541 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_542 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_543 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_544 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_545 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_546 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_547 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_548 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_549 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_550 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_551 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_552 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_553 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_554 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_555 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_556 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_557 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_558 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_559 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_560 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_561 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_562 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_563 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_564 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_565 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_566 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_567 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_568 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_569 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_570 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_571 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_572 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_573 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_574 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_575 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_576 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_577 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_578 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_579 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_580 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_581 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   b;
  assign sum = b;

endmodule


module mul_csa32_582 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_583 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_584 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_585 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_586 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_587 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_588 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_589 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_590 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_591 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_592 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_593 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_594 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_595 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_596 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_597 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_598 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_599 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_600 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_601 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_602 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_603 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_604 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_605 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_606 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_607 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_608 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_609 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_610 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_611 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_612 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_613 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_614 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_615 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_616 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_617 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_618 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_619 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_620 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_621 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_622 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_623 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_624 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_625 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_626 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_627 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_628 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_629 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_630 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_631 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_632 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_633 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_634 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_635 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_636 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_637 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_638 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_639 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_640 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_641 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_642 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_643 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_644 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_645 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_646 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_647 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_648 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_649 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_650 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_651 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_652 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_653 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_654 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_655 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_656 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_657 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_658 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_659 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_660 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(c), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(c), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa42_1 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(n2), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(carry) );
  OA21X1_RVT U3 ( .A1(n2), .A2(b), .A3(n1), .Y(sum) );
  FADDX1_RVT U4 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n2) );
endmodule


module mul_csa42_2 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_3 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_4 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_5 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_6 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_7 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_8 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_9 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_10 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_11 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_12 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_13 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_14 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_15 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_16 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_17 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_18 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_19 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_20 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_21 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_22 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_23 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_24 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_25 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_26 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_27 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_28 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_29 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_30 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_31 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_32 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_33 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_34 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_35 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_36 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_37 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_38 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_39 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_40 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_41 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_42 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_43 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_44 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_45 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_46 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_47 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_48 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_49 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;


  FADDX1_RVT U1 ( .A(c), .B(b), .CI(cin), .CO(carry), .S(sum) );
endmodule


module mul_array2 ( pcout, pcoutx2, psum, psumx2, a0c, a0s, a1c, a1s, areg, 
        bot, pc, ps, x2 );
  output [98:0] pcout;
  output [98:0] psum;
  input [81:4] a0c;
  input [81:0] a0s;
  input [81:4] a1c;
  input [81:0] a1s;
  input [96:0] areg;
  input [98:30] pc;
  input [98:31] ps;
  input bot, x2;
  output pcoutx2, psumx2;
  wire   net210786, net210787, net210788, net210789, net210790, net210791,
         net210792, net210793, net210794, net210795, net210796, net210797,
         net210798, net210799, net210800, net210801, net210802, net210803,
         net210804, net210805, net210806, net210807, net210808, net210809,
         net210810, net210811, net210812, net210813, net210814, net210815,
         net210816, net210817, net210818, net210819, net210820, net210821,
         net210822, net210823, net210824, net210825, net210826, net210827,
         net210828, net210829, net210830, net210831, net210832, net210833,
         net210834, net210835, net210836, net210837, net210838, net210839,
         net210840, net210841, net210842, net210843, net210844, net210845,
         net210846, net210847, net210848, net210849, net210850, net210851,
         net210852, net210853, net210854, net210855, net210856, net210857,
         net210858, net210859, net210860, net210861, net210862, net210863,
         net210864, net210865, net210866, net210867, net210868, net210869,
         net210870, net210871, net210872, net210873, net210874, net210875,
         net210876, net210877, net210878, net210879, net210880, net210881,
         net210882, net210883, net210884, net210885, net210886, net210887,
         net210888, net210889;
  wire   [67:20] co;
  wire   [81:15] c3;
  wire   [96:0] c2;
  wire   [96:0] s2;
  wire   [81:15] s3;
  wire   [82:0] s1;
  wire   [82:0] c1;

  mul_csa42_49 sc3_68_ ( .sum(s3[68]), .carry(c3[68]), .a(1'b0), .b(s2[68]), 
        .c(c2[67]), .d(1'b0), .cin(co[67]) );
  mul_csa42_48 sc3_67_ ( .sum(s3[67]), .carry(c3[67]), .cout(co[67]), .a(
        s1[67]), .b(s2[67]), .c(c2[66]), .d(1'b0), .cin(co[66]) );
  mul_csa42_47 sc3_66_ ( .sum(s3[66]), .carry(c3[66]), .cout(co[66]), .a(
        s1[66]), .b(s2[66]), .c(c2[65]), .d(c1[65]), .cin(co[65]) );
  mul_csa42_46 sc3_65_ ( .sum(s3[65]), .carry(c3[65]), .cout(co[65]), .a(
        s1[65]), .b(s2[65]), .c(c2[64]), .d(c1[64]), .cin(co[64]) );
  mul_csa42_45 sc3_64_ ( .sum(s3[64]), .carry(c3[64]), .cout(co[64]), .a(
        s1[64]), .b(s2[64]), .c(c2[63]), .d(c1[63]), .cin(co[63]) );
  mul_csa42_44 sc3_63_ ( .sum(s3[63]), .carry(c3[63]), .cout(co[63]), .a(
        s1[63]), .b(s2[63]), .c(c2[62]), .d(c1[62]), .cin(co[62]) );
  mul_csa42_43 sc3_62_ ( .sum(s3[62]), .carry(c3[62]), .cout(co[62]), .a(
        s1[62]), .b(s2[62]), .c(c2[61]), .d(c1[61]), .cin(co[61]) );
  mul_csa42_42 sc3_61_ ( .sum(s3[61]), .carry(c3[61]), .cout(co[61]), .a(
        s1[61]), .b(s2[61]), .c(c2[60]), .d(c1[60]), .cin(co[60]) );
  mul_csa42_41 sc3_60_ ( .sum(s3[60]), .carry(c3[60]), .cout(co[60]), .a(
        s1[60]), .b(s2[60]), .c(c2[59]), .d(c1[59]), .cin(co[59]) );
  mul_csa42_40 sc3_59_ ( .sum(s3[59]), .carry(c3[59]), .cout(co[59]), .a(
        s1[59]), .b(s2[59]), .c(c2[58]), .d(c1[58]), .cin(co[58]) );
  mul_csa42_39 sc3_58_ ( .sum(s3[58]), .carry(c3[58]), .cout(co[58]), .a(
        s1[58]), .b(s2[58]), .c(c2[57]), .d(c1[57]), .cin(co[57]) );
  mul_csa42_38 sc3_57_ ( .sum(s3[57]), .carry(c3[57]), .cout(co[57]), .a(
        s1[57]), .b(s2[57]), .c(c2[56]), .d(c1[56]), .cin(co[56]) );
  mul_csa42_37 sc3_56_ ( .sum(s3[56]), .carry(c3[56]), .cout(co[56]), .a(
        s1[56]), .b(s2[56]), .c(c2[55]), .d(c1[55]), .cin(co[55]) );
  mul_csa42_36 sc3_55_ ( .sum(s3[55]), .carry(c3[55]), .cout(co[55]), .a(
        s1[55]), .b(s2[55]), .c(c2[54]), .d(c1[54]), .cin(co[54]) );
  mul_csa42_35 sc3_54_ ( .sum(s3[54]), .carry(c3[54]), .cout(co[54]), .a(
        s1[54]), .b(s2[54]), .c(c2[53]), .d(c1[53]), .cin(co[53]) );
  mul_csa42_34 sc3_53_ ( .sum(s3[53]), .carry(c3[53]), .cout(co[53]), .a(
        s1[53]), .b(s2[53]), .c(c2[52]), .d(c1[52]), .cin(co[52]) );
  mul_csa42_33 sc3_52_ ( .sum(s3[52]), .carry(c3[52]), .cout(co[52]), .a(
        s1[52]), .b(s2[52]), .c(c2[51]), .d(c1[51]), .cin(co[51]) );
  mul_csa42_32 sc3_51_ ( .sum(s3[51]), .carry(c3[51]), .cout(co[51]), .a(
        s1[51]), .b(s2[51]), .c(c2[50]), .d(c1[50]), .cin(co[50]) );
  mul_csa42_31 sc3_50_ ( .sum(s3[50]), .carry(c3[50]), .cout(co[50]), .a(
        s1[50]), .b(s2[50]), .c(c2[49]), .d(c1[49]), .cin(co[49]) );
  mul_csa42_30 sc3_49_ ( .sum(s3[49]), .carry(c3[49]), .cout(co[49]), .a(
        s1[49]), .b(s2[49]), .c(c2[48]), .d(c1[48]), .cin(co[48]) );
  mul_csa42_29 sc3_48_ ( .sum(s3[48]), .carry(c3[48]), .cout(co[48]), .a(
        s1[48]), .b(s2[48]), .c(c2[47]), .d(c1[47]), .cin(co[47]) );
  mul_csa42_28 sc3_47_ ( .sum(s3[47]), .carry(c3[47]), .cout(co[47]), .a(
        s1[47]), .b(s2[47]), .c(c2[46]), .d(c1[46]), .cin(co[46]) );
  mul_csa42_27 sc3_46_ ( .sum(s3[46]), .carry(c3[46]), .cout(co[46]), .a(
        s1[46]), .b(s2[46]), .c(c2[45]), .d(c1[45]), .cin(co[45]) );
  mul_csa42_26 sc3_45_ ( .sum(s3[45]), .carry(c3[45]), .cout(co[45]), .a(
        s1[45]), .b(s2[45]), .c(c2[44]), .d(c1[44]), .cin(co[44]) );
  mul_csa42_25 sc3_44_ ( .sum(s3[44]), .carry(c3[44]), .cout(co[44]), .a(
        s1[44]), .b(s2[44]), .c(c2[43]), .d(c1[43]), .cin(co[43]) );
  mul_csa42_24 sc3_43_ ( .sum(s3[43]), .carry(c3[43]), .cout(co[43]), .a(
        s1[43]), .b(s2[43]), .c(c2[42]), .d(c1[42]), .cin(co[42]) );
  mul_csa42_23 sc3_42_ ( .sum(s3[42]), .carry(c3[42]), .cout(co[42]), .a(
        s1[42]), .b(s2[42]), .c(c2[41]), .d(c1[41]), .cin(co[41]) );
  mul_csa42_22 sc3_41_ ( .sum(s3[41]), .carry(c3[41]), .cout(co[41]), .a(
        s1[41]), .b(s2[41]), .c(c2[40]), .d(c1[40]), .cin(co[40]) );
  mul_csa42_21 sc3_40_ ( .sum(s3[40]), .carry(c3[40]), .cout(co[40]), .a(
        s1[40]), .b(s2[40]), .c(c2[39]), .d(c1[39]), .cin(co[39]) );
  mul_csa42_20 sc3_39_ ( .sum(s3[39]), .carry(c3[39]), .cout(co[39]), .a(
        s1[39]), .b(s2[39]), .c(c2[38]), .d(c1[38]), .cin(co[38]) );
  mul_csa42_19 sc3_38_ ( .sum(s3[38]), .carry(c3[38]), .cout(co[38]), .a(
        s1[38]), .b(s2[38]), .c(c2[37]), .d(c1[37]), .cin(co[37]) );
  mul_csa42_18 sc3_37_ ( .sum(s3[37]), .carry(c3[37]), .cout(co[37]), .a(
        s1[37]), .b(s2[37]), .c(c2[36]), .d(c1[36]), .cin(co[36]) );
  mul_csa42_17 sc3_36_ ( .sum(s3[36]), .carry(c3[36]), .cout(co[36]), .a(
        s1[36]), .b(s2[36]), .c(c2[35]), .d(c1[35]), .cin(co[35]) );
  mul_csa42_16 sc3_35_ ( .sum(s3[35]), .carry(c3[35]), .cout(co[35]), .a(
        s1[35]), .b(s2[35]), .c(c2[34]), .d(c1[34]), .cin(co[34]) );
  mul_csa42_15 sc3_34_ ( .sum(s3[34]), .carry(c3[34]), .cout(co[34]), .a(
        s1[34]), .b(s2[34]), .c(c2[33]), .d(c1[33]), .cin(co[33]) );
  mul_csa42_14 sc3_33_ ( .sum(s3[33]), .carry(c3[33]), .cout(co[33]), .a(
        s1[33]), .b(s2[33]), .c(c2[32]), .d(c1[32]), .cin(co[32]) );
  mul_csa42_13 sc3_32_ ( .sum(s3[32]), .carry(c3[32]), .cout(co[32]), .a(
        s1[32]), .b(s2[32]), .c(c2[31]), .d(c1[31]), .cin(co[31]) );
  mul_csa42_12 sc3_31_ ( .sum(s3[31]), .carry(c3[31]), .cout(co[31]), .a(
        s1[31]), .b(s2[31]), .c(c2[30]), .d(c1[30]), .cin(co[30]) );
  mul_csa42_11 sc3_30_ ( .sum(s3[30]), .carry(c3[30]), .cout(co[30]), .a(
        s1[30]), .b(s2[30]), .c(c2[29]), .d(c1[29]), .cin(co[29]) );
  mul_csa42_10 sc3_29_ ( .sum(s3[29]), .carry(c3[29]), .cout(co[29]), .a(
        s1[29]), .b(s2[29]), .c(c2[28]), .d(c1[28]), .cin(co[28]) );
  mul_csa42_9 sc3_28_ ( .sum(s3[28]), .carry(c3[28]), .cout(co[28]), .a(s1[28]), .b(s2[28]), .c(c2[27]), .d(c1[27]), .cin(co[27]) );
  mul_csa42_8 sc3_27_ ( .sum(s3[27]), .carry(c3[27]), .cout(co[27]), .a(s1[27]), .b(s2[27]), .c(c2[26]), .d(c1[26]), .cin(co[26]) );
  mul_csa42_7 sc3_26_ ( .sum(s3[26]), .carry(c3[26]), .cout(co[26]), .a(s1[26]), .b(s2[26]), .c(c2[25]), .d(c1[25]), .cin(co[25]) );
  mul_csa42_6 sc3_25_ ( .sum(s3[25]), .carry(c3[25]), .cout(co[25]), .a(s1[25]), .b(s2[25]), .c(c2[24]), .d(c1[24]), .cin(co[24]) );
  mul_csa42_5 sc3_24_ ( .sum(s3[24]), .carry(c3[24]), .cout(co[24]), .a(s1[24]), .b(s2[24]), .c(c2[23]), .d(c1[23]), .cin(co[23]) );
  mul_csa42_4 sc3_23_ ( .sum(s3[23]), .carry(c3[23]), .cout(co[23]), .a(s1[23]), .b(s2[23]), .c(c2[22]), .d(c1[22]), .cin(co[22]) );
  mul_csa42_3 sc3_22_ ( .sum(s3[22]), .carry(c3[22]), .cout(co[22]), .a(s1[22]), .b(s2[22]), .c(c2[21]), .d(c1[21]), .cin(co[21]) );
  mul_csa42_2 sc3_21_ ( .sum(s3[21]), .carry(c3[21]), .cout(co[21]), .a(s1[21]), .b(s2[21]), .c(c2[20]), .d(c1[20]), .cin(co[20]) );
  mul_csa42_1 sc3_20_ ( .sum(s3[20]), .carry(c3[20]), .cout(co[20]), .a(s1[20]), .b(s2[20]), .c(c2[19]), .d(c1[19]), .cin(1'b0) );
  mul_csa32_660 sc4_82_ ( .sum(psum[82]), .cout(pcout[82]), .a(net210889), .b(
        s2[82]), .c(c3[81]) );
  mul_csa32_659 sc4_68_ ( .sum(psum[68]), .cout(pcout[68]), .a(net210888), .b(
        s3[68]), .c(c3[67]) );
  mul_csa32_658 sc4_67_ ( .sum(psum[67]), .cout(pcout[67]), .a(net210887), .b(
        s3[67]), .c(c3[66]) );
  mul_csa32_657 sc4_66_ ( .sum(psum[66]), .cout(pcout[66]), .a(net210886), .b(
        s3[66]), .c(c3[65]) );
  mul_csa32_656 sc4_65_ ( .sum(psum[65]), .cout(pcout[65]), .a(net210885), .b(
        s3[65]), .c(c3[64]) );
  mul_csa32_655 sc4_64_ ( .sum(psum[64]), .cout(pcout[64]), .a(net210884), .b(
        s3[64]), .c(c3[63]) );
  mul_csa32_654 sc4_63_ ( .sum(psum[63]), .cout(pcout[63]), .a(net210883), .b(
        s3[63]), .c(c3[62]) );
  mul_csa32_653 sc4_62_ ( .sum(psum[62]), .cout(pcout[62]), .a(net210882), .b(
        s3[62]), .c(c3[61]) );
  mul_csa32_652 sc4_61_ ( .sum(psum[61]), .cout(pcout[61]), .a(net210881), .b(
        s3[61]), .c(c3[60]) );
  mul_csa32_651 sc4_60_ ( .sum(psum[60]), .cout(pcout[60]), .a(net210880), .b(
        s3[60]), .c(c3[59]) );
  mul_csa32_650 sc4_59_ ( .sum(psum[59]), .cout(pcout[59]), .a(net210879), .b(
        s3[59]), .c(c3[58]) );
  mul_csa32_649 sc4_58_ ( .sum(psum[58]), .cout(pcout[58]), .a(net210878), .b(
        s3[58]), .c(c3[57]) );
  mul_csa32_648 sc4_57_ ( .sum(psum[57]), .cout(pcout[57]), .a(net210877), .b(
        s3[57]), .c(c3[56]) );
  mul_csa32_647 sc4_56_ ( .sum(psum[56]), .cout(pcout[56]), .a(net210876), .b(
        s3[56]), .c(c3[55]) );
  mul_csa32_646 sc4_55_ ( .sum(psum[55]), .cout(pcout[55]), .a(net210875), .b(
        s3[55]), .c(c3[54]) );
  mul_csa32_645 sc4_54_ ( .sum(psum[54]), .cout(pcout[54]), .a(net210874), .b(
        s3[54]), .c(c3[53]) );
  mul_csa32_644 sc4_53_ ( .sum(psum[53]), .cout(pcout[53]), .a(net210873), .b(
        s3[53]), .c(c3[52]) );
  mul_csa32_643 sc4_52_ ( .sum(psum[52]), .cout(pcout[52]), .a(net210872), .b(
        s3[52]), .c(c3[51]) );
  mul_csa32_642 sc4_51_ ( .sum(psum[51]), .cout(pcout[51]), .a(net210871), .b(
        s3[51]), .c(c3[50]) );
  mul_csa32_641 sc4_50_ ( .sum(psum[50]), .cout(pcout[50]), .a(net210870), .b(
        s3[50]), .c(c3[49]) );
  mul_csa32_640 sc4_49_ ( .sum(psum[49]), .cout(pcout[49]), .a(net210869), .b(
        s3[49]), .c(c3[48]) );
  mul_csa32_639 sc4_48_ ( .sum(psum[48]), .cout(pcout[48]), .a(net210868), .b(
        s3[48]), .c(c3[47]) );
  mul_csa32_638 sc4_47_ ( .sum(psum[47]), .cout(pcout[47]), .a(net210867), .b(
        s3[47]), .c(c3[46]) );
  mul_csa32_637 sc4_46_ ( .sum(psum[46]), .cout(pcout[46]), .a(net210866), .b(
        s3[46]), .c(c3[45]) );
  mul_csa32_636 sc4_45_ ( .sum(psum[45]), .cout(pcout[45]), .a(net210865), .b(
        s3[45]), .c(c3[44]) );
  mul_csa32_635 sc4_44_ ( .sum(psum[44]), .cout(pcout[44]), .a(net210864), .b(
        s3[44]), .c(c3[43]) );
  mul_csa32_634 sc4_43_ ( .sum(psum[43]), .cout(pcout[43]), .a(net210863), .b(
        s3[43]), .c(c3[42]) );
  mul_csa32_633 sc4_42_ ( .sum(psum[42]), .cout(pcout[42]), .a(net210862), .b(
        s3[42]), .c(c3[41]) );
  mul_csa32_632 sc4_41_ ( .sum(psum[41]), .cout(pcout[41]), .a(net210861), .b(
        s3[41]), .c(c3[40]) );
  mul_csa32_631 sc4_40_ ( .sum(psum[40]), .cout(pcout[40]), .a(net210860), .b(
        s3[40]), .c(c3[39]) );
  mul_csa32_630 sc4_39_ ( .sum(psum[39]), .cout(pcout[39]), .a(net210859), .b(
        s3[39]), .c(c3[38]) );
  mul_csa32_629 sc4_38_ ( .sum(psum[38]), .cout(pcout[38]), .a(net210858), .b(
        s3[38]), .c(c3[37]) );
  mul_csa32_628 sc4_37_ ( .sum(psum[37]), .cout(pcout[37]), .a(net210857), .b(
        s3[37]), .c(c3[36]) );
  mul_csa32_627 sc4_36_ ( .sum(psum[36]), .cout(pcout[36]), .a(net210856), .b(
        s3[36]), .c(c3[35]) );
  mul_csa32_626 sc4_35_ ( .sum(psum[35]), .cout(pcout[35]), .a(net210855), .b(
        s3[35]), .c(c3[34]) );
  mul_csa32_625 sc4_34_ ( .sum(psum[34]), .cout(pcout[34]), .a(net210854), .b(
        s3[34]), .c(c3[33]) );
  mul_csa32_624 sc4_33_ ( .sum(psum[33]), .cout(pcout[33]), .a(net210853), .b(
        s3[33]), .c(c3[32]) );
  mul_csa32_623 sc4_32_ ( .sum(psum[32]), .cout(pcout[32]), .a(net210852), .b(
        s3[32]), .c(c3[31]) );
  mul_csa32_622 sc4_31_ ( .sum(psum[31]), .cout(pcout[31]), .a(net210851), .b(
        s3[31]), .c(c3[30]) );
  mul_csa32_621 sc4_30_ ( .sum(psum[30]), .cout(pcout[30]), .a(net210850), .b(
        s3[30]), .c(c3[29]) );
  mul_csa32_620 sc4_29_ ( .sum(psum[29]), .cout(pcout[29]), .a(net210849), .b(
        s3[29]), .c(c3[28]) );
  mul_csa32_619 sc4_28_ ( .sum(psum[28]), .cout(pcout[28]), .a(net210848), .b(
        s3[28]), .c(c3[27]) );
  mul_csa32_618 sc4_27_ ( .sum(psum[27]), .cout(pcout[27]), .a(net210847), .b(
        s3[27]), .c(c3[26]) );
  mul_csa32_617 sc4_26_ ( .sum(psum[26]), .cout(pcout[26]), .a(net210846), .b(
        s3[26]), .c(c3[25]) );
  mul_csa32_616 sc4_25_ ( .sum(psum[25]), .cout(pcout[25]), .a(net210845), .b(
        s3[25]), .c(c3[24]) );
  mul_csa32_615 sc4_24_ ( .sum(psum[24]), .cout(pcout[24]), .a(net210844), .b(
        s3[24]), .c(c3[23]) );
  mul_csa32_614 sc4_23_ ( .sum(psum[23]), .cout(pcout[23]), .a(net210843), .b(
        s3[23]), .c(c3[22]) );
  mul_csa32_613 sc4_22_ ( .sum(psum[22]), .cout(pcout[22]), .a(net210842), .b(
        s3[22]), .c(c3[21]) );
  mul_csa32_612 sc4_21_ ( .sum(psum[21]), .cout(pcout[21]), .a(net210841), .b(
        s3[21]), .c(c3[20]) );
  mul_csa32_611 sc4_20_ ( .sum(psum[20]), .cout(pcout[20]), .a(net210840), .b(
        s3[20]), .c(c3[19]) );
  mul_csa32_610 sc4_96_ ( .sum(psum[96]), .cout(pcout[96]), .a(net210839), .b(
        s2[96]), .c(c2[95]) );
  mul_csa32_609 sc4_95_ ( .sum(psum[95]), .cout(pcout[95]), .a(net210838), .b(
        s2[95]), .c(c2[94]) );
  mul_csa32_608 sc4_94_ ( .sum(psum[94]), .cout(pcout[94]), .a(net210837), .b(
        s2[94]), .c(c2[93]) );
  mul_csa32_607 sc4_93_ ( .sum(psum[93]), .cout(pcout[93]), .a(net210836), .b(
        s2[93]), .c(c2[92]) );
  mul_csa32_606 sc4_92_ ( .sum(psum[92]), .cout(pcout[92]), .a(net210835), .b(
        s2[92]), .c(c2[91]) );
  mul_csa32_605 sc4_91_ ( .sum(psum[91]), .cout(pcout[91]), .a(net210834), .b(
        s2[91]), .c(c2[90]) );
  mul_csa32_604 sc4_90_ ( .sum(psum[90]), .cout(pcout[90]), .a(net210833), .b(
        s2[90]), .c(c2[89]) );
  mul_csa32_603 sc4_89_ ( .sum(psum[89]), .cout(pcout[89]), .a(net210832), .b(
        s2[89]), .c(c2[88]) );
  mul_csa32_602 sc4_88_ ( .sum(psum[88]), .cout(pcout[88]), .a(net210831), .b(
        s2[88]), .c(c2[87]) );
  mul_csa32_601 sc4_87_ ( .sum(psum[87]), .cout(pcout[87]), .a(net210830), .b(
        s2[87]), .c(c2[86]) );
  mul_csa32_600 sc4_86_ ( .sum(psum[86]), .cout(pcout[86]), .a(net210829), .b(
        s2[86]), .c(c2[85]) );
  mul_csa32_599 sc4_85_ ( .sum(psum[85]), .cout(pcout[85]), .a(net210828), .b(
        s2[85]), .c(c2[84]) );
  mul_csa32_598 sc4_84_ ( .sum(psum[84]), .cout(pcout[84]), .a(net210827), .b(
        s2[84]), .c(c2[83]) );
  mul_csa32_597 sc4_81_ ( .sum(psum[81]), .cout(pcout[81]), .a(net210826), .b(
        s3[81]), .c(c3[80]) );
  mul_csa32_596 sc4_80_ ( .sum(psum[80]), .cout(pcout[80]), .a(net210825), .b(
        s3[80]), .c(c3[79]) );
  mul_csa32_595 sc4_79_ ( .sum(psum[79]), .cout(pcout[79]), .a(net210824), .b(
        s3[79]), .c(c3[78]) );
  mul_csa32_594 sc4_78_ ( .sum(psum[78]), .cout(pcout[78]), .a(net210823), .b(
        s3[78]), .c(c3[77]) );
  mul_csa32_593 sc4_77_ ( .sum(psum[77]), .cout(pcout[77]), .a(net210822), .b(
        s3[77]), .c(c3[76]) );
  mul_csa32_592 sc4_76_ ( .sum(psum[76]), .cout(pcout[76]), .a(net210821), .b(
        s3[76]), .c(c3[75]) );
  mul_csa32_591 sc4_75_ ( .sum(psum[75]), .cout(pcout[75]), .a(net210820), .b(
        s3[75]), .c(c3[74]) );
  mul_csa32_590 sc4_74_ ( .sum(psum[74]), .cout(pcout[74]), .a(net210819), .b(
        s3[74]), .c(c3[73]) );
  mul_csa32_589 sc4_73_ ( .sum(psum[73]), .cout(pcout[73]), .a(net210818), .b(
        s3[73]), .c(c3[72]) );
  mul_csa32_588 sc4_72_ ( .sum(psum[72]), .cout(pcout[72]), .a(net210817), .b(
        s3[72]), .c(c3[71]) );
  mul_csa32_587 sc4_71_ ( .sum(psum[71]), .cout(pcout[71]), .a(net210816), .b(
        s3[71]), .c(c3[70]) );
  mul_csa32_586 sc4_70_ ( .sum(psum[70]), .cout(pcout[70]), .a(net210815), .b(
        s3[70]), .c(c3[69]) );
  mul_csa32_585 sc4_69_ ( .sum(psum[69]), .cout(pcout[69]), .a(net210814), .b(
        s3[69]), .c(c3[68]) );
  mul_csa32_584 acc_4_ ( .sum(psum[4]), .cout(pcout[4]), .a(net210813), .b(
        s2[4]), .c(c2[3]) );
  mul_csa32_583 acc_3_ ( .sum(psum[3]), .cout(pcout[3]), .a(net210812), .b(
        s2[3]), .c(c2[2]) );
  mul_csa32_582 acc_2_ ( .sum(psum[2]), .cout(pcout[2]), .a(net210811), .b(
        s2[2]), .c(c2[1]) );
  mul_csa32_581 acc_1_ ( .sum(psum[1]), .a(net210809), .b(s2[1]), .c(net210810) );
  mul_csa32_580 sc3_97_ ( .sum(psum[97]), .cout(pcout[97]), .a(a1s[81]), .b(
        net210808), .c(c2[96]) );
  mul_csa32_579 sc1_19_ ( .sum(s1[19]), .cout(c1[19]), .a(ps[51]), .b(pc[50]), 
        .c(a1s[3]) );
  mul_csa32_578 sc1_18_ ( .sum(s1[18]), .cout(c1[18]), .a(ps[50]), .b(pc[49]), 
        .c(a1s[2]) );
  mul_csa32_577 sc1_17_ ( .sum(s1[17]), .cout(c1[17]), .a(ps[49]), .b(pc[48]), 
        .c(a1s[1]) );
  mul_csa32_576 sc1_16_ ( .sum(s1[16]), .cout(c1[16]), .a(ps[48]), .b(pc[47]), 
        .c(a1s[0]) );
  mul_csa32_575 sc1_15_ ( .sum(s1[15]), .cout(c1[15]), .a(ps[47]), .b(pc[46]), 
        .c(1'b0) );
  mul_csa32_574 sc4_83_ ( .sum(psum[83]), .cout(pcout[83]), .a(net210807), .b(
        s2[83]), .c(c2[82]) );
  mul_csa32_573 sc2_83_ ( .sum(s2[83]), .cout(c2[83]), .a(a1s[67]), .b(a1c[66]), .c(c1[82]) );
  mul_csa32_572 sc2_19_ ( .sum(s2[19]), .cout(c2[19]), .a(s1[19]), .b(a0s[19]), 
        .c(a0c[18]) );
  mul_csa32_571 sc2_18_ ( .sum(s2[18]), .cout(c2[18]), .a(s1[18]), .b(a0s[18]), 
        .c(a0c[17]) );
  mul_csa32_570 sc2_17_ ( .sum(s2[17]), .cout(c2[17]), .a(s1[17]), .b(a0s[17]), 
        .c(a0c[16]) );
  mul_csa32_569 sc2_16_ ( .sum(s2[16]), .cout(c2[16]), .a(s1[16]), .b(a0s[16]), 
        .c(a0c[15]) );
  mul_csa32_568 sc2_15_ ( .sum(s2[15]), .cout(c2[15]), .a(s1[15]), .b(a0s[15]), 
        .c(a0c[14]) );
  mul_csa32_567 sc1_81_ ( .sum(s1[81]), .cout(c1[81]), .a(a1s[65]), .b(a1c[64]), .c(net210806) );
  mul_csa32_566 sc1_80_ ( .sum(s1[80]), .cout(c1[80]), .a(a1s[64]), .b(a1c[63]), .c(a0s[80]) );
  mul_csa32_565 sc1_79_ ( .sum(s1[79]), .cout(c1[79]), .a(a1s[63]), .b(a1c[62]), .c(a0s[79]) );
  mul_csa32_564 sc1_78_ ( .sum(s1[78]), .cout(c1[78]), .a(a1s[62]), .b(a1c[61]), .c(a0s[78]) );
  mul_csa32_563 sc1_77_ ( .sum(s1[77]), .cout(c1[77]), .a(a1s[61]), .b(a1c[60]), .c(a0s[77]) );
  mul_csa32_562 sc1_76_ ( .sum(s1[76]), .cout(c1[76]), .a(a1s[60]), .b(a1c[59]), .c(a0s[76]) );
  mul_csa32_561 sc1_75_ ( .sum(s1[75]), .cout(c1[75]), .a(a1s[59]), .b(a1c[58]), .c(a0s[75]) );
  mul_csa32_560 sc1_74_ ( .sum(s1[74]), .cout(c1[74]), .a(a1s[58]), .b(a1c[57]), .c(a0s[74]) );
  mul_csa32_559 sc1_73_ ( .sum(s1[73]), .cout(c1[73]), .a(a1s[57]), .b(a1c[56]), .c(a0s[73]) );
  mul_csa32_558 sc1_72_ ( .sum(s1[72]), .cout(c1[72]), .a(a1s[56]), .b(a1c[55]), .c(a0s[72]) );
  mul_csa32_557 sc1_71_ ( .sum(s1[71]), .cout(c1[71]), .a(a1s[55]), .b(a1c[54]), .c(a0s[71]) );
  mul_csa32_556 sc1_70_ ( .sum(s1[70]), .cout(c1[70]), .a(a1s[54]), .b(a1c[53]), .c(a0s[70]) );
  mul_csa32_555 sc1_69_ ( .sum(s1[69]), .cout(c1[69]), .a(a1s[53]), .b(a1c[52]), .c(a0s[69]) );
  mul_csa32_554 sc1_68_ ( .sum(s1[68]), .cout(c1[68]), .a(a1s[52]), .b(a1c[51]), .c(a0s[68]) );
  mul_csa32_553 sc3_19_ ( .sum(s3[19]), .cout(c3[19]), .a(s2[19]), .b(c1[18]), 
        .c(c2[18]) );
  mul_csa32_552 sc3_18_ ( .sum(s3[18]), .cout(c3[18]), .a(s2[18]), .b(c1[17]), 
        .c(c2[17]) );
  mul_csa32_551 sc3_17_ ( .sum(s3[17]), .cout(c3[17]), .a(s2[17]), .b(c1[16]), 
        .c(c2[16]) );
  mul_csa32_550 sc3_16_ ( .sum(s3[16]), .cout(c3[16]), .a(s2[16]), .b(c1[15]), 
        .c(c2[15]) );
  mul_csa32_549 sc3_15_ ( .sum(s3[15]), .cout(c3[15]), .a(s2[15]), .b(c1[14]), 
        .c(c2[14]) );
  mul_csa32_548 sc1_82_ ( .sum(s1[82]), .cout(c1[82]), .a(a1s[66]), .b(a1c[65]), .c(net210805) );
  mul_csa32_547 acc_14_ ( .sum(psum[14]), .cout(pcout[14]), .a(net210804), .b(
        s2[14]), .c(c2[13]) );
  mul_csa32_546 acc_13_ ( .sum(psum[13]), .cout(pcout[13]), .a(net210803), .b(
        s2[13]), .c(c2[12]) );
  mul_csa32_545 acc_12_ ( .sum(psum[12]), .cout(pcout[12]), .a(net210802), .b(
        s2[12]), .c(c2[11]) );
  mul_csa32_544 acc_11_ ( .sum(psum[11]), .cout(pcout[11]), .a(net210801), .b(
        s2[11]), .c(c2[10]) );
  mul_csa32_543 acc_10_ ( .sum(psum[10]), .cout(pcout[10]), .a(net210800), .b(
        s2[10]), .c(c2[9]) );
  mul_csa32_542 acc_9_ ( .sum(psum[9]), .cout(pcout[9]), .a(net210799), .b(
        s2[9]), .c(c2[8]) );
  mul_csa32_541 acc_8_ ( .sum(psum[8]), .cout(pcout[8]), .a(net210798), .b(
        s2[8]), .c(c2[7]) );
  mul_csa32_540 acc_7_ ( .sum(psum[7]), .cout(pcout[7]), .a(net210797), .b(
        s2[7]), .c(c2[6]) );
  mul_csa32_539 acc_6_ ( .sum(psum[6]), .cout(pcout[6]), .a(net210796), .b(
        s2[6]), .c(c2[5]) );
  mul_csa32_538 acc_5_ ( .sum(psum[5]), .cout(pcout[5]), .a(net210795), .b(
        s2[5]), .c(c2[4]) );
  mul_csa32_537 sc2_67_ ( .sum(s2[67]), .cout(c2[67]), .a(a0s[67]), .b(c1[66]), 
        .c(a0c[66]) );
  mul_csa32_536 sc1_14_ ( .sum(s1[14]), .cout(c1[14]), .a(ps[46]), .b(pc[45]), 
        .c(a0s[14]) );
  mul_csa32_535 sc1_13_ ( .sum(s1[13]), .cout(c1[13]), .a(ps[45]), .b(pc[44]), 
        .c(a0s[13]) );
  mul_csa32_534 sc1_12_ ( .sum(s1[12]), .cout(c1[12]), .a(ps[44]), .b(pc[43]), 
        .c(a0s[12]) );
  mul_csa32_533 sc1_11_ ( .sum(s1[11]), .cout(c1[11]), .a(ps[43]), .b(pc[42]), 
        .c(a0s[11]) );
  mul_csa32_532 sc1_10_ ( .sum(s1[10]), .cout(c1[10]), .a(ps[42]), .b(pc[41]), 
        .c(a0s[10]) );
  mul_csa32_531 sc1_9_ ( .sum(s1[9]), .cout(c1[9]), .a(ps[41]), .b(pc[40]), 
        .c(a0s[9]) );
  mul_csa32_530 sc1_8_ ( .sum(s1[8]), .cout(c1[8]), .a(ps[40]), .b(pc[39]), 
        .c(a0s[8]) );
  mul_csa32_529 sc1_7_ ( .sum(s1[7]), .cout(c1[7]), .a(ps[39]), .b(pc[38]), 
        .c(a0s[7]) );
  mul_csa32_528 sc1_6_ ( .sum(s1[6]), .cout(c1[6]), .a(ps[38]), .b(pc[37]), 
        .c(a0s[6]) );
  mul_csa32_527 sc1_5_ ( .sum(s1[5]), .cout(c1[5]), .a(ps[37]), .b(pc[36]), 
        .c(a0s[5]) );
  mul_csa32_526 sc2_14_ ( .sum(s2[14]), .cout(c2[14]), .a(s1[14]), .b(c1[13]), 
        .c(a0c[13]) );
  mul_csa32_525 sc2_13_ ( .sum(s2[13]), .cout(c2[13]), .a(s1[13]), .b(c1[12]), 
        .c(a0c[12]) );
  mul_csa32_524 sc2_12_ ( .sum(s2[12]), .cout(c2[12]), .a(s1[12]), .b(c1[11]), 
        .c(a0c[11]) );
  mul_csa32_523 sc2_11_ ( .sum(s2[11]), .cout(c2[11]), .a(s1[11]), .b(c1[10]), 
        .c(a0c[10]) );
  mul_csa32_522 sc2_10_ ( .sum(s2[10]), .cout(c2[10]), .a(s1[10]), .b(c1[9]), 
        .c(a0c[9]) );
  mul_csa32_521 sc2_9_ ( .sum(s2[9]), .cout(c2[9]), .a(s1[9]), .b(c1[8]), .c(
        a0c[8]) );
  mul_csa32_520 sc2_8_ ( .sum(s2[8]), .cout(c2[8]), .a(s1[8]), .b(c1[7]), .c(
        a0c[7]) );
  mul_csa32_519 sc2_7_ ( .sum(s2[7]), .cout(c2[7]), .a(s1[7]), .b(c1[6]), .c(
        a0c[6]) );
  mul_csa32_518 sc2_6_ ( .sum(s2[6]), .cout(c2[6]), .a(s1[6]), .b(c1[5]), .c(
        a0c[5]) );
  mul_csa32_517 sc2_5_ ( .sum(s2[5]), .cout(c2[5]), .a(s1[5]), .b(c1[4]), .c(
        a0c[4]) );
  mul_csa32_516 sc2_82_ ( .sum(s2[82]), .cout(c2[82]), .a(s1[82]), .b(c1[81]), 
        .c(c2[81]) );
  mul_csa32_515 sc1_4_ ( .sum(s1[4]), .cout(c1[4]), .a(ps[36]), .b(pc[35]), 
        .c(a0s[4]) );
  mul_csa32_514 sc1_3_ ( .sum(s1[3]), .cout(c1[3]), .a(ps[35]), .b(pc[34]), 
        .c(a0s[3]) );
  mul_csa32_513 sc1_2_ ( .sum(s1[2]), .cout(c1[2]), .a(ps[34]), .b(pc[33]), 
        .c(a0s[2]) );
  mul_csa32_512 sc1_1_ ( .sum(s1[1]), .cout(c1[1]), .a(ps[33]), .b(pc[32]), 
        .c(a0s[1]) );
  mul_csa32_511 sc2_66_ ( .sum(s2[66]), .cout(c2[66]), .a(a1c[49]), .b(a0s[66]), .c(a0c[65]) );
  mul_csa32_510 sc2_65_ ( .sum(s2[65]), .cout(c2[65]), .a(a1c[48]), .b(a0s[65]), .c(a0c[64]) );
  mul_csa32_509 sc2_64_ ( .sum(s2[64]), .cout(c2[64]), .a(a1c[47]), .b(a0s[64]), .c(a0c[63]) );
  mul_csa32_508 sc2_63_ ( .sum(s2[63]), .cout(c2[63]), .a(a1c[46]), .b(a0s[63]), .c(a0c[62]) );
  mul_csa32_507 sc2_62_ ( .sum(s2[62]), .cout(c2[62]), .a(a1c[45]), .b(a0s[62]), .c(a0c[61]) );
  mul_csa32_506 sc2_61_ ( .sum(s2[61]), .cout(c2[61]), .a(a1c[44]), .b(a0s[61]), .c(a0c[60]) );
  mul_csa32_505 sc2_60_ ( .sum(s2[60]), .cout(c2[60]), .a(a1c[43]), .b(a0s[60]), .c(a0c[59]) );
  mul_csa32_504 sc2_59_ ( .sum(s2[59]), .cout(c2[59]), .a(a1c[42]), .b(a0s[59]), .c(a0c[58]) );
  mul_csa32_503 sc2_58_ ( .sum(s2[58]), .cout(c2[58]), .a(a1c[41]), .b(a0s[58]), .c(a0c[57]) );
  mul_csa32_502 sc2_57_ ( .sum(s2[57]), .cout(c2[57]), .a(a1c[40]), .b(a0s[57]), .c(a0c[56]) );
  mul_csa32_501 sc2_56_ ( .sum(s2[56]), .cout(c2[56]), .a(a1c[39]), .b(a0s[56]), .c(a0c[55]) );
  mul_csa32_500 sc2_55_ ( .sum(s2[55]), .cout(c2[55]), .a(a1c[38]), .b(a0s[55]), .c(a0c[54]) );
  mul_csa32_499 sc2_54_ ( .sum(s2[54]), .cout(c2[54]), .a(a1c[37]), .b(a0s[54]), .c(a0c[53]) );
  mul_csa32_498 sc2_53_ ( .sum(s2[53]), .cout(c2[53]), .a(a1c[36]), .b(a0s[53]), .c(a0c[52]) );
  mul_csa32_497 sc2_52_ ( .sum(s2[52]), .cout(c2[52]), .a(a1c[35]), .b(a0s[52]), .c(a0c[51]) );
  mul_csa32_496 sc2_51_ ( .sum(s2[51]), .cout(c2[51]), .a(a1c[34]), .b(a0s[51]), .c(a0c[50]) );
  mul_csa32_495 sc2_50_ ( .sum(s2[50]), .cout(c2[50]), .a(a1c[33]), .b(a0s[50]), .c(a0c[49]) );
  mul_csa32_494 sc2_49_ ( .sum(s2[49]), .cout(c2[49]), .a(a1c[32]), .b(a0s[49]), .c(a0c[48]) );
  mul_csa32_493 sc2_48_ ( .sum(s2[48]), .cout(c2[48]), .a(a1c[31]), .b(a0s[48]), .c(a0c[47]) );
  mul_csa32_492 sc2_47_ ( .sum(s2[47]), .cout(c2[47]), .a(a1c[30]), .b(a0s[47]), .c(a0c[46]) );
  mul_csa32_491 sc2_46_ ( .sum(s2[46]), .cout(c2[46]), .a(a1c[29]), .b(a0s[46]), .c(a0c[45]) );
  mul_csa32_490 sc2_45_ ( .sum(s2[45]), .cout(c2[45]), .a(a1c[28]), .b(a0s[45]), .c(a0c[44]) );
  mul_csa32_489 sc2_44_ ( .sum(s2[44]), .cout(c2[44]), .a(a1c[27]), .b(a0s[44]), .c(a0c[43]) );
  mul_csa32_488 sc2_43_ ( .sum(s2[43]), .cout(c2[43]), .a(a1c[26]), .b(a0s[43]), .c(a0c[42]) );
  mul_csa32_487 sc2_42_ ( .sum(s2[42]), .cout(c2[42]), .a(a1c[25]), .b(a0s[42]), .c(a0c[41]) );
  mul_csa32_486 sc2_41_ ( .sum(s2[41]), .cout(c2[41]), .a(a1c[24]), .b(a0s[41]), .c(a0c[40]) );
  mul_csa32_485 sc2_40_ ( .sum(s2[40]), .cout(c2[40]), .a(a1c[23]), .b(a0s[40]), .c(a0c[39]) );
  mul_csa32_484 sc2_39_ ( .sum(s2[39]), .cout(c2[39]), .a(a1c[22]), .b(a0s[39]), .c(a0c[38]) );
  mul_csa32_483 sc2_38_ ( .sum(s2[38]), .cout(c2[38]), .a(a1c[21]), .b(a0s[38]), .c(a0c[37]) );
  mul_csa32_482 sc2_37_ ( .sum(s2[37]), .cout(c2[37]), .a(a1c[20]), .b(a0s[37]), .c(a0c[36]) );
  mul_csa32_481 sc2_36_ ( .sum(s2[36]), .cout(c2[36]), .a(a1c[19]), .b(a0s[36]), .c(a0c[35]) );
  mul_csa32_480 sc2_35_ ( .sum(s2[35]), .cout(c2[35]), .a(a1c[18]), .b(a0s[35]), .c(a0c[34]) );
  mul_csa32_479 sc2_34_ ( .sum(s2[34]), .cout(c2[34]), .a(a1c[17]), .b(a0s[34]), .c(a0c[33]) );
  mul_csa32_478 sc2_33_ ( .sum(s2[33]), .cout(c2[33]), .a(a1c[16]), .b(a0s[33]), .c(a0c[32]) );
  mul_csa32_477 sc2_32_ ( .sum(s2[32]), .cout(c2[32]), .a(a1c[15]), .b(a0s[32]), .c(a0c[31]) );
  mul_csa32_476 sc2_31_ ( .sum(s2[31]), .cout(c2[31]), .a(a1c[14]), .b(a0s[31]), .c(a0c[30]) );
  mul_csa32_475 sc2_30_ ( .sum(s2[30]), .cout(c2[30]), .a(a1c[13]), .b(a0s[30]), .c(a0c[29]) );
  mul_csa32_474 sc2_29_ ( .sum(s2[29]), .cout(c2[29]), .a(a1c[12]), .b(a0s[29]), .c(a0c[28]) );
  mul_csa32_473 sc2_28_ ( .sum(s2[28]), .cout(c2[28]), .a(a1c[11]), .b(a0s[28]), .c(a0c[27]) );
  mul_csa32_472 sc2_27_ ( .sum(s2[27]), .cout(c2[27]), .a(a1c[10]), .b(a0s[27]), .c(a0c[26]) );
  mul_csa32_471 sc2_26_ ( .sum(s2[26]), .cout(c2[26]), .a(a1c[9]), .b(a0s[26]), 
        .c(a0c[25]) );
  mul_csa32_470 sc2_25_ ( .sum(s2[25]), .cout(c2[25]), .a(a1c[8]), .b(a0s[25]), 
        .c(a0c[24]) );
  mul_csa32_469 sc2_24_ ( .sum(s2[24]), .cout(c2[24]), .a(a1c[7]), .b(a0s[24]), 
        .c(a0c[23]) );
  mul_csa32_468 sc2_23_ ( .sum(s2[23]), .cout(c2[23]), .a(a1c[6]), .b(a0s[23]), 
        .c(a0c[22]) );
  mul_csa32_467 sc2_22_ ( .sum(s2[22]), .cout(c2[22]), .a(a1c[5]), .b(a0s[22]), 
        .c(a0c[21]) );
  mul_csa32_466 sc2_21_ ( .sum(s2[21]), .cout(c2[21]), .a(a1c[4]), .b(a0s[21]), 
        .c(a0c[20]) );
  mul_csa32_465 sc2_20_ ( .sum(s2[20]), .cout(c2[20]), .a(1'b0), .b(a0s[20]), 
        .c(a0c[19]) );
  mul_csa32_464 sc1_66_ ( .sum(s1[66]), .cout(c1[66]), .a(ps[98]), .b(pc[97]), 
        .c(a1s[50]) );
  mul_csa32_463 sc1_65_ ( .sum(s1[65]), .cout(c1[65]), .a(ps[97]), .b(pc[96]), 
        .c(a1s[49]) );
  mul_csa32_462 sc1_64_ ( .sum(s1[64]), .cout(c1[64]), .a(ps[96]), .b(pc[95]), 
        .c(a1s[48]) );
  mul_csa32_461 sc1_63_ ( .sum(s1[63]), .cout(c1[63]), .a(ps[95]), .b(pc[94]), 
        .c(a1s[47]) );
  mul_csa32_460 sc1_62_ ( .sum(s1[62]), .cout(c1[62]), .a(ps[94]), .b(pc[93]), 
        .c(a1s[46]) );
  mul_csa32_459 sc1_61_ ( .sum(s1[61]), .cout(c1[61]), .a(ps[93]), .b(pc[92]), 
        .c(a1s[45]) );
  mul_csa32_458 sc1_60_ ( .sum(s1[60]), .cout(c1[60]), .a(ps[92]), .b(pc[91]), 
        .c(a1s[44]) );
  mul_csa32_457 sc1_59_ ( .sum(s1[59]), .cout(c1[59]), .a(ps[91]), .b(pc[90]), 
        .c(a1s[43]) );
  mul_csa32_456 sc1_58_ ( .sum(s1[58]), .cout(c1[58]), .a(ps[90]), .b(pc[89]), 
        .c(a1s[42]) );
  mul_csa32_455 sc1_57_ ( .sum(s1[57]), .cout(c1[57]), .a(ps[89]), .b(pc[88]), 
        .c(a1s[41]) );
  mul_csa32_454 sc1_56_ ( .sum(s1[56]), .cout(c1[56]), .a(ps[88]), .b(pc[87]), 
        .c(a1s[40]) );
  mul_csa32_453 sc1_55_ ( .sum(s1[55]), .cout(c1[55]), .a(ps[87]), .b(pc[86]), 
        .c(a1s[39]) );
  mul_csa32_452 sc1_54_ ( .sum(s1[54]), .cout(c1[54]), .a(ps[86]), .b(pc[85]), 
        .c(a1s[38]) );
  mul_csa32_451 sc1_53_ ( .sum(s1[53]), .cout(c1[53]), .a(ps[85]), .b(pc[84]), 
        .c(a1s[37]) );
  mul_csa32_450 sc1_52_ ( .sum(s1[52]), .cout(c1[52]), .a(ps[84]), .b(pc[83]), 
        .c(a1s[36]) );
  mul_csa32_449 sc1_51_ ( .sum(s1[51]), .cout(c1[51]), .a(ps[83]), .b(pc[82]), 
        .c(a1s[35]) );
  mul_csa32_448 sc1_50_ ( .sum(s1[50]), .cout(c1[50]), .a(ps[82]), .b(pc[81]), 
        .c(a1s[34]) );
  mul_csa32_447 sc1_49_ ( .sum(s1[49]), .cout(c1[49]), .a(ps[81]), .b(pc[80]), 
        .c(a1s[33]) );
  mul_csa32_446 sc1_48_ ( .sum(s1[48]), .cout(c1[48]), .a(ps[80]), .b(pc[79]), 
        .c(a1s[32]) );
  mul_csa32_445 sc1_47_ ( .sum(s1[47]), .cout(c1[47]), .a(ps[79]), .b(pc[78]), 
        .c(a1s[31]) );
  mul_csa32_444 sc1_46_ ( .sum(s1[46]), .cout(c1[46]), .a(ps[78]), .b(pc[77]), 
        .c(a1s[30]) );
  mul_csa32_443 sc1_45_ ( .sum(s1[45]), .cout(c1[45]), .a(ps[77]), .b(pc[76]), 
        .c(a1s[29]) );
  mul_csa32_442 sc1_44_ ( .sum(s1[44]), .cout(c1[44]), .a(ps[76]), .b(pc[75]), 
        .c(a1s[28]) );
  mul_csa32_441 sc1_43_ ( .sum(s1[43]), .cout(c1[43]), .a(ps[75]), .b(pc[74]), 
        .c(a1s[27]) );
  mul_csa32_440 sc1_42_ ( .sum(s1[42]), .cout(c1[42]), .a(ps[74]), .b(pc[73]), 
        .c(a1s[26]) );
  mul_csa32_439 sc1_41_ ( .sum(s1[41]), .cout(c1[41]), .a(ps[73]), .b(pc[72]), 
        .c(a1s[25]) );
  mul_csa32_438 sc1_40_ ( .sum(s1[40]), .cout(c1[40]), .a(ps[72]), .b(pc[71]), 
        .c(a1s[24]) );
  mul_csa32_437 sc1_39_ ( .sum(s1[39]), .cout(c1[39]), .a(ps[71]), .b(pc[70]), 
        .c(a1s[23]) );
  mul_csa32_436 sc1_38_ ( .sum(s1[38]), .cout(c1[38]), .a(ps[70]), .b(pc[69]), 
        .c(a1s[22]) );
  mul_csa32_435 sc1_37_ ( .sum(s1[37]), .cout(c1[37]), .a(ps[69]), .b(pc[68]), 
        .c(a1s[21]) );
  mul_csa32_434 sc1_36_ ( .sum(s1[36]), .cout(c1[36]), .a(ps[68]), .b(pc[67]), 
        .c(a1s[20]) );
  mul_csa32_433 sc1_35_ ( .sum(s1[35]), .cout(c1[35]), .a(ps[67]), .b(pc[66]), 
        .c(a1s[19]) );
  mul_csa32_432 sc1_34_ ( .sum(s1[34]), .cout(c1[34]), .a(ps[66]), .b(pc[65]), 
        .c(a1s[18]) );
  mul_csa32_431 sc1_33_ ( .sum(s1[33]), .cout(c1[33]), .a(ps[65]), .b(pc[64]), 
        .c(a1s[17]) );
  mul_csa32_430 sc1_32_ ( .sum(s1[32]), .cout(c1[32]), .a(ps[64]), .b(pc[63]), 
        .c(a1s[16]) );
  mul_csa32_429 sc1_31_ ( .sum(s1[31]), .cout(c1[31]), .a(ps[63]), .b(pc[62]), 
        .c(a1s[15]) );
  mul_csa32_428 sc1_30_ ( .sum(s1[30]), .cout(c1[30]), .a(ps[62]), .b(pc[61]), 
        .c(a1s[14]) );
  mul_csa32_427 sc1_29_ ( .sum(s1[29]), .cout(c1[29]), .a(ps[61]), .b(pc[60]), 
        .c(a1s[13]) );
  mul_csa32_426 sc1_28_ ( .sum(s1[28]), .cout(c1[28]), .a(ps[60]), .b(pc[59]), 
        .c(a1s[12]) );
  mul_csa32_425 sc1_27_ ( .sum(s1[27]), .cout(c1[27]), .a(ps[59]), .b(pc[58]), 
        .c(a1s[11]) );
  mul_csa32_424 sc1_26_ ( .sum(s1[26]), .cout(c1[26]), .a(ps[58]), .b(pc[57]), 
        .c(a1s[10]) );
  mul_csa32_423 sc1_25_ ( .sum(s1[25]), .cout(c1[25]), .a(ps[57]), .b(pc[56]), 
        .c(a1s[9]) );
  mul_csa32_422 sc1_24_ ( .sum(s1[24]), .cout(c1[24]), .a(ps[56]), .b(pc[55]), 
        .c(a1s[8]) );
  mul_csa32_421 sc1_23_ ( .sum(s1[23]), .cout(c1[23]), .a(ps[55]), .b(pc[54]), 
        .c(a1s[7]) );
  mul_csa32_420 sc1_22_ ( .sum(s1[22]), .cout(c1[22]), .a(ps[54]), .b(pc[53]), 
        .c(a1s[6]) );
  mul_csa32_419 sc1_21_ ( .sum(s1[21]), .cout(c1[21]), .a(ps[53]), .b(pc[52]), 
        .c(a1s[5]) );
  mul_csa32_418 sc1_20_ ( .sum(s1[20]), .cout(c1[20]), .a(ps[52]), .b(pc[51]), 
        .c(a1s[4]) );
  mul_csa32_417 sc2_81_ ( .sum(s2[81]), .cout(c2[81]), .a(s1[81]), .b(c1[80]), 
        .c(net210794) );
  mul_csa32_416 sc2_80_ ( .sum(s2[80]), .cout(c2[80]), .a(s1[80]), .b(c1[79]), 
        .c(a0c[79]) );
  mul_csa32_415 sc2_79_ ( .sum(s2[79]), .cout(c2[79]), .a(s1[79]), .b(c1[78]), 
        .c(a0c[78]) );
  mul_csa32_414 sc2_78_ ( .sum(s2[78]), .cout(c2[78]), .a(s1[78]), .b(c1[77]), 
        .c(a0c[77]) );
  mul_csa32_413 sc2_77_ ( .sum(s2[77]), .cout(c2[77]), .a(s1[77]), .b(c1[76]), 
        .c(a0c[76]) );
  mul_csa32_412 sc2_76_ ( .sum(s2[76]), .cout(c2[76]), .a(s1[76]), .b(c1[75]), 
        .c(a0c[75]) );
  mul_csa32_411 sc2_75_ ( .sum(s2[75]), .cout(c2[75]), .a(s1[75]), .b(c1[74]), 
        .c(a0c[74]) );
  mul_csa32_410 sc2_74_ ( .sum(s2[74]), .cout(c2[74]), .a(s1[74]), .b(c1[73]), 
        .c(a0c[73]) );
  mul_csa32_409 sc2_73_ ( .sum(s2[73]), .cout(c2[73]), .a(s1[73]), .b(c1[72]), 
        .c(a0c[72]) );
  mul_csa32_408 sc2_72_ ( .sum(s2[72]), .cout(c2[72]), .a(s1[72]), .b(c1[71]), 
        .c(a0c[71]) );
  mul_csa32_407 sc2_71_ ( .sum(s2[71]), .cout(c2[71]), .a(s1[71]), .b(c1[70]), 
        .c(a0c[70]) );
  mul_csa32_406 sc2_70_ ( .sum(s2[70]), .cout(c2[70]), .a(s1[70]), .b(c1[69]), 
        .c(a0c[69]) );
  mul_csa32_405 sc2_69_ ( .sum(s2[69]), .cout(c2[69]), .a(s1[69]), .b(c1[68]), 
        .c(a0c[68]) );
  mul_csa32_404 sc2_68_ ( .sum(s2[68]), .cout(c2[68]), .a(s1[68]), .b(c1[67]), 
        .c(a0c[67]) );
  mul_csa32_403 acc_19_ ( .sum(psum[19]), .cout(pcout[19]), .a(net210793), .b(
        s3[19]), .c(c3[18]) );
  mul_csa32_402 acc_18_ ( .sum(psum[18]), .cout(pcout[18]), .a(net210792), .b(
        s3[18]), .c(c3[17]) );
  mul_csa32_401 acc_17_ ( .sum(psum[17]), .cout(pcout[17]), .a(net210791), .b(
        s3[17]), .c(c3[16]) );
  mul_csa32_400 acc_16_ ( .sum(psum[16]), .cout(pcout[16]), .a(net210790), .b(
        s3[16]), .c(c3[15]) );
  mul_csa32_399 acc_15_ ( .sum(psum[15]), .a(net210789), .b(s3[15]), .c(1'b0)
         );
  mul_csa32_398 sc1_0_ ( .sum(s1[0]), .cout(c1[0]), .a(ps[32]), .b(pc[31]), 
        .c(a0s[0]) );
  mul_csa32_397 sc1_67_ ( .sum(s1[67]), .cout(c1[67]), .a(a1s[51]), .b(
        net210788), .c(a1c[50]) );
  mul_ha_47 acc_0_ ( .sum(psum[0]), .a(net210787), .b(s2[0]) );
  mul_ha_45 sc2_96_ ( .cout(c2[96]), .sum(s2[96]), .a(a1s[80]), .b(a1c[79]) );
  mul_ha_44 sc2_95_ ( .cout(c2[95]), .sum(s2[95]), .a(a1s[79]), .b(a1c[78]) );
  mul_ha_43 sc2_94_ ( .cout(c2[94]), .sum(s2[94]), .a(a1s[78]), .b(a1c[77]) );
  mul_ha_42 sc2_93_ ( .cout(c2[93]), .sum(s2[93]), .a(a1s[77]), .b(a1c[76]) );
  mul_ha_41 sc2_92_ ( .cout(c2[92]), .sum(s2[92]), .a(a1s[76]), .b(a1c[75]) );
  mul_ha_40 sc2_91_ ( .cout(c2[91]), .sum(s2[91]), .a(a1s[75]), .b(a1c[74]) );
  mul_ha_39 sc2_90_ ( .cout(c2[90]), .sum(s2[90]), .a(a1s[74]), .b(a1c[73]) );
  mul_ha_38 sc2_89_ ( .cout(c2[89]), .sum(s2[89]), .a(a1s[73]), .b(a1c[72]) );
  mul_ha_37 sc2_88_ ( .cout(c2[88]), .sum(s2[88]), .a(a1s[72]), .b(a1c[71]) );
  mul_ha_36 sc2_87_ ( .cout(c2[87]), .sum(s2[87]), .a(a1s[71]), .b(a1c[70]) );
  mul_ha_35 sc2_86_ ( .cout(c2[86]), .sum(s2[86]), .a(a1s[70]), .b(a1c[69]) );
  mul_ha_34 sc2_85_ ( .cout(c2[85]), .sum(s2[85]), .a(a1s[69]), .b(a1c[68]) );
  mul_ha_33 sc2_84_ ( .cout(c2[84]), .sum(s2[84]), .a(a1s[68]), .b(a1c[67]) );
  mul_ha_32 sc3_81_ ( .cout(c3[81]), .sum(s3[81]), .a(s2[81]), .b(c2[80]) );
  mul_ha_31 sc3_80_ ( .cout(c3[80]), .sum(s3[80]), .a(s2[80]), .b(c2[79]) );
  mul_ha_30 sc3_79_ ( .cout(c3[79]), .sum(s3[79]), .a(s2[79]), .b(c2[78]) );
  mul_ha_29 sc3_78_ ( .cout(c3[78]), .sum(s3[78]), .a(s2[78]), .b(c2[77]) );
  mul_ha_28 sc3_77_ ( .cout(c3[77]), .sum(s3[77]), .a(s2[77]), .b(c2[76]) );
  mul_ha_27 sc3_76_ ( .cout(c3[76]), .sum(s3[76]), .a(s2[76]), .b(c2[75]) );
  mul_ha_26 sc3_75_ ( .cout(c3[75]), .sum(s3[75]), .a(s2[75]), .b(c2[74]) );
  mul_ha_25 sc3_74_ ( .cout(c3[74]), .sum(s3[74]), .a(s2[74]), .b(c2[73]) );
  mul_ha_24 sc3_73_ ( .cout(c3[73]), .sum(s3[73]), .a(s2[73]), .b(c2[72]) );
  mul_ha_23 sc3_72_ ( .cout(c3[72]), .sum(s3[72]), .a(s2[72]), .b(c2[71]) );
  mul_ha_22 sc3_71_ ( .cout(c3[71]), .sum(s3[71]), .a(s2[71]), .b(c2[70]) );
  mul_ha_21 sc3_70_ ( .cout(c3[70]), .sum(s3[70]), .a(s2[70]), .b(c2[69]) );
  mul_ha_20 sc3_69_ ( .cout(c3[69]), .sum(s3[69]), .a(s2[69]), .b(c2[68]) );
  mul_ha_18 sc2_4_ ( .cout(c2[4]), .sum(s2[4]), .a(s1[4]), .b(c1[3]) );
  mul_ha_17 sc2_3_ ( .cout(c2[3]), .sum(s2[3]), .a(s1[3]), .b(c1[2]) );
  mul_ha_16 sc2_2_ ( .cout(c2[2]), .sum(s2[2]), .a(s1[2]), .b(c1[1]) );
  mul_ha_15 sc2_1_ ( .cout(c2[1]), .sum(s2[1]), .a(s1[1]), .b(c1[0]) );
  mul_ha_14 sc2_0_ ( .sum(s2[0]), .a(s1[0]), .b(net210786) );
endmodule


module dp_mux2es_SIZE97 ( dout, in0, in1, sel );
  output [96:0] dout;
  input [96:0] in0;
  input [96:0] in1;
  input sel;

  assign dout[72] = in0[72];
  assign dout[71] = in0[71];
  assign dout[70] = in0[70];
  assign dout[69] = in0[69];
  assign dout[68] = in0[68];
  assign dout[67] = in0[67];
  assign dout[66] = in0[66];
  assign dout[65] = in0[65];
  assign dout[64] = in0[64];
  assign dout[63] = in0[63];
  assign dout[62] = in0[62];
  assign dout[61] = in0[61];
  assign dout[60] = in0[60];
  assign dout[59] = in0[59];
  assign dout[58] = in0[58];
  assign dout[57] = in0[57];
  assign dout[56] = in0[56];
  assign dout[55] = in0[55];
  assign dout[54] = in0[54];
  assign dout[53] = in0[53];
  assign dout[52] = in0[52];
  assign dout[51] = in0[51];
  assign dout[50] = in0[50];
  assign dout[49] = in0[49];
  assign dout[48] = in0[48];
  assign dout[47] = in0[47];
  assign dout[46] = in0[46];
  assign dout[45] = in0[45];
  assign dout[44] = in0[44];
  assign dout[43] = in0[43];
  assign dout[42] = in0[42];
  assign dout[41] = in0[41];
  assign dout[40] = in0[40];
  assign dout[39] = in0[39];
  assign dout[38] = in0[38];
  assign dout[37] = in0[37];
  assign dout[36] = in0[36];
  assign dout[35] = in0[35];
  assign dout[34] = in0[34];
  assign dout[33] = in0[33];
  assign dout[32] = in0[32];
  assign dout[31] = in0[31];
  assign dout[30] = in0[30];
  assign dout[29] = in0[29];
  assign dout[28] = in0[28];
  assign dout[27] = in0[27];
  assign dout[26] = in0[26];
  assign dout[25] = in0[25];
  assign dout[24] = in0[24];
  assign dout[23] = in0[23];
  assign dout[22] = in0[22];
  assign dout[21] = in0[21];
  assign dout[20] = in0[20];
  assign dout[19] = in0[19];
  assign dout[18] = in0[18];
  assign dout[17] = in0[17];
  assign dout[16] = in0[16];
  assign dout[14] = in0[14];
  assign dout[13] = in0[13];
  assign dout[12] = in0[12];
  assign dout[11] = in0[11];
  assign dout[10] = in0[10];
  assign dout[9] = in0[9];
  assign dout[8] = in0[8];
  assign dout[7] = in0[7];
  assign dout[6] = in0[6];
  assign dout[5] = in0[5];
  assign dout[4] = in0[4];
  assign dout[3] = in0[3];
  assign dout[2] = in0[2];

endmodule


module dp_mux2es_SIZE98 ( dout, in0, in1, sel );
  output [97:0] dout;
  input [97:0] in0;
  input [97:0] in1;
  input sel;

  assign dout[73] = in0[73];
  assign dout[72] = in0[72];
  assign dout[71] = in0[71];
  assign dout[70] = in0[70];
  assign dout[69] = in0[69];
  assign dout[68] = in0[68];
  assign dout[67] = in0[67];
  assign dout[66] = in0[66];
  assign dout[65] = in0[65];
  assign dout[64] = in0[64];
  assign dout[63] = in0[63];
  assign dout[62] = in0[62];
  assign dout[61] = in0[61];
  assign dout[60] = in0[60];
  assign dout[59] = in0[59];
  assign dout[58] = in0[58];
  assign dout[57] = in0[57];
  assign dout[56] = in0[56];
  assign dout[55] = in0[55];
  assign dout[54] = in0[54];
  assign dout[53] = in0[53];
  assign dout[52] = in0[52];
  assign dout[51] = in0[51];
  assign dout[50] = in0[50];
  assign dout[49] = in0[49];
  assign dout[48] = in0[48];
  assign dout[47] = in0[47];
  assign dout[46] = in0[46];
  assign dout[45] = in0[45];
  assign dout[44] = in0[44];
  assign dout[43] = in0[43];
  assign dout[42] = in0[42];
  assign dout[41] = in0[41];
  assign dout[40] = in0[40];
  assign dout[39] = in0[39];
  assign dout[38] = in0[38];
  assign dout[37] = in0[37];
  assign dout[36] = in0[36];
  assign dout[35] = in0[35];
  assign dout[34] = in0[34];
  assign dout[33] = in0[33];
  assign dout[32] = in0[32];
  assign dout[31] = in0[31];
  assign dout[30] = in0[30];
  assign dout[29] = in0[29];
  assign dout[28] = in0[28];
  assign dout[27] = in0[27];
  assign dout[26] = in0[26];
  assign dout[25] = in0[25];
  assign dout[24] = in0[24];
  assign dout[23] = in0[23];
  assign dout[22] = in0[22];
  assign dout[21] = in0[21];
  assign dout[20] = in0[20];
  assign dout[19] = in0[19];
  assign dout[18] = in0[18];
  assign dout[17] = in0[17];
  assign dout[16] = in0[16];
  assign dout[15] = in0[15];
  assign dout[14] = in0[14];
  assign dout[13] = in0[13];
  assign dout[12] = in0[12];
  assign dout[11] = in0[11];
  assign dout[10] = in0[10];
  assign dout[9] = in0[9];
  assign dout[8] = in0[8];
  assign dout[7] = in0[7];
  assign dout[6] = in0[6];
  assign dout[5] = in0[5];
  assign dout[4] = in0[4];
  assign dout[3] = in0[3];
  assign dout[2] = in0[2];
  assign dout[1] = in0[1];
  assign dout[0] = in0[0];

endmodule


module mul_ppgen_187 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_188 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_189 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_190 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_191 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_192 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_2 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_csa32_63 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_64 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_65 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  OR2X1_RVT U1 ( .A1(a), .A2(c), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(a), .A2(c), .Y(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(cout), .Y(sum) );
endmodule


module mul_csa32_66 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ppgensign_1 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_2 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_3 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_1 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net42, net47, p2_l_67, net073, p1_l_65, net38, net0118, p2_l_66,
         net078, p2_l_65, net8, p2_l_64, net15, p1_l_64, net43, net48, net35;

  mul_ppgensign_3 p0_64_ ( .p_l(net42), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_2 p2_68_ ( .p_l(sum[5]), .z(net073), .b(b2), .pm1_l(p2_l_67)
         );
  mul_ppgensign_1 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ha_2 sc1_68_ ( .cout(cout[4]), .sum(sum[4]), .a(1'b1), .b(net073) );
  mul_ppgen_192 p2_67_ ( .p_l(p2_l_67), .z(net078), .a(am1), .b(b2), .pm1_l(
        p2_l_66) );
  mul_ppgen_191 p2_66_ ( .p_l(p2_l_66), .z(net8), .a(am2), .b(b2), .pm1_l(
        p2_l_65) );
  mul_ppgen_190 p2_65_ ( .p_l(p2_l_65), .z(net15), .a(am3), .b(b2), .pm1_l(
        p2_l_64) );
  mul_ppgen_189 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_188 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_ppgen_187 p2_64_ ( .p_l(p2_l_64), .z(net35), .a(am4), .b(b2), .pm1_l(
        p2m1_l) );
  mul_csa32_66 sc1_67_ ( .sum(sum[3]), .cout(cout[3]), .a(net0118), .b(1'b0), 
        .c(net078) );
  mul_csa32_65 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(1'b1), 
        .c(net8) );
  mul_csa32_64 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net15) );
  mul_csa32_63 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net35) );
endmodule


module mul_ppgen_1 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_2 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_3 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_4 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_5 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_6 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_1 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_1 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_2 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_1 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_2 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_1 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_2 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_1 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_2 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_1 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_1 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_6 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_5 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_4 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(p0_l_1)
         );
  mul_ppgen_3 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(p0_l_0)
         );
  mul_ppgen_2 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_1 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_7 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_8 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_9 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_csa32_3 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_1 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043, net210263;

  mul_csa32_3 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_9 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(net210263)
         );
  mul_ppgen_8 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_7 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_10 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_11 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_12 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_4 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_2 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_4 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_12 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_11 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_10 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_13 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_14 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_15 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_5 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_3 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_5 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_15 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_14 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_13 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_16 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_17 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_18 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_6 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_4 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_6 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_18 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_17 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_16 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_19 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_20 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_21 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_7 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_5 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_7 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_21 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_20 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_19 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_22 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_23 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_24 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_8 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_6 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_8 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_24 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_23 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_22 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_25 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_26 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_27 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_9 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_7 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_9 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_27 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_26 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_25 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_28 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_29 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_30 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_10 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_8 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_10 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_30 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_29 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_28 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_31 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_32 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_33 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_11 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_9 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_11 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_33 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_32 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_31 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_34 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_35 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_36 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_12 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_10 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_12 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_36 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_35 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_34 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_37 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_38 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_39 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_13 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_11 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_13 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_39 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_38 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_37 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_40 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_41 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_42 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_14 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_12 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_14 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_42 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_41 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_40 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_43 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_44 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_45 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_15 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_13 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_15 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_45 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_44 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_43 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_46 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_47 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_48 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_16 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_14 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_16 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_48 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_47 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_46 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_49 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_50 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_51 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_17 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_15 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_17 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_51 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_50 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_49 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_52 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_53 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_54 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_18 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_16 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_18 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_54 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_53 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_52 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_55 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_56 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_57 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_19 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_17 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_19 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_57 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_56 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_55 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_58 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_59 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_60 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_20 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_18 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_20 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_60 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_59 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_58 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_61 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_62 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_63 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_21 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_19 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_21 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_63 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_62 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_61 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_64 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_65 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_66 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_22 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_20 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_22 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_66 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_65 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_64 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_67 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_68 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_69 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_23 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_21 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_23 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_69 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_68 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_67 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_70 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_71 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_72 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_24 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_22 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_24 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_72 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_71 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_70 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_73 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_74 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_75 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_25 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_23 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_25 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_75 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_74 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_73 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_76 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_77 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_78 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_26 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_24 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_26 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_78 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_77 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_76 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_79 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_80 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_81 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_27 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_25 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_27 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_81 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_80 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_79 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_82 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_83 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_84 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_28 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_26 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_28 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_84 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_83 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_82 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_85 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_86 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_87 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_29 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_27 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_29 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_87 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_86 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_85 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_88 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_89 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_90 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_30 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_28 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_30 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_90 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_89 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_88 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_91 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_92 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_93 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_31 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_29 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_31 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_93 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_92 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_91 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_94 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_95 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_96 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_32 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_30 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_32 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_96 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_95 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_94 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_97 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_98 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_99 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_33 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_31 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_33 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_99 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen_98 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen_97 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_100 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_101 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_102 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_34 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_32 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_34 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_102 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_101 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_100 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_103 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_104 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_105 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_35 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_33 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_35 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_105 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_104 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_103 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_106 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_107 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_108 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_36 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_34 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_36 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_108 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_107 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_106 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_109 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_110 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_111 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_37 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_35 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_37 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_111 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_110 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_109 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_112 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_113 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_114 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_38 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_36 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_38 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_114 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_113 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_112 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_115 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_116 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_117 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_39 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_37 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_39 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_117 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_116 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_115 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_118 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_119 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_120 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_40 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_38 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_40 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_120 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_119 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_118 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_121 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_122 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_123 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_41 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_39 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_41 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_123 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_122 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_121 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_124 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_125 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_126 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_42 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_40 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_42 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_126 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_125 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_124 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_127 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_128 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_129 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_43 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_41 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_43 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_129 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_128 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_127 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_130 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_131 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_132 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_44 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_42 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_44 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_132 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_131 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_130 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_133 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_134 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_135 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_45 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_43 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_45 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_135 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_134 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_133 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_136 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_137 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_138 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_46 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_44 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_46 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_138 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_137 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_136 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_139 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_140 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_141 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_47 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_45 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_47 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_141 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_140 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_139 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_142 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_143 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_144 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_48 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_46 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_48 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_144 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_143 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_142 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_145 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_146 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_147 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_49 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_47 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_49 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_147 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_146 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_145 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_148 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_149 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_150 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_50 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_48 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_50 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_150 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_149 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_148 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_151 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_152 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_153 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_51 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_49 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_51 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_153 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_152 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_151 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_154 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_155 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_156 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_52 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_50 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_52 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_156 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_155 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_154 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_157 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_158 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_159 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_53 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_51 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_53 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_159 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_158 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_157 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_160 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_161 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_162 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_54 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_52 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_54 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_162 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_161 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_160 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_163 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_164 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_165 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_55 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_53 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_55 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_165 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_164 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_163 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_166 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_167 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_168 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_56 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_54 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_56 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_168 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_167 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_166 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_169 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_170 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_171 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_57 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_55 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_57 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_171 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_170 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_169 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_172 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_173 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_174 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_58 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_56 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_58 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_174 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_173 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_172 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_175 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_176 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_177 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_59 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_57 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_59 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_177 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_176 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_175 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_178 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_179 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_180 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_60 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_58 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_60 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_180 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_179 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_178 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_181 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_182 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_183 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_61 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_59 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_61 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_183 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_182 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_181 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_184 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_185 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_186 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_62 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_60 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_62 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_186 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_185 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_184 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_1 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210526, net210527;
  wire   [63:4] p2_l;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;

  mul_ppgen3sign_1 I2 ( .cout(cout[68:64]), .sum(sum[69:64]), .am1(a[63]), 
        .am2(a[62]), .am3(a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2(b2), 
        .bot(net210526), .head(net210527), .p0m1_l(p0_l[63]), .p1m1_l(p1_l[63]), .p2m1_l(p2_l[63]) );
  mul_ppgen3_60 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .p2_l(p2_l[63]), .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[62]), .p1m1_l(p1_l[62]), 
        .p2m1_l(p2_l[62]) );
  mul_ppgen3_59 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .p2_l(p2_l[62]), .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[61]), .p1m1_l(p1_l[61]), 
        .p2m1_l(p2_l[61]) );
  mul_ppgen3_58 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .p2_l(p2_l[61]), .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[60]), .p1m1_l(p1_l[60]), 
        .p2m1_l(p2_l[60]) );
  mul_ppgen3_57 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .p2_l(p2_l[60]), .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[59]), .p1m1_l(p1_l[59]), 
        .p2m1_l(p2_l[59]) );
  mul_ppgen3_56 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .p2_l(p2_l[59]), .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[58]), .p1m1_l(p1_l[58]), 
        .p2m1_l(p2_l[58]) );
  mul_ppgen3_55 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .p2_l(p2_l[58]), .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[57]), .p1m1_l(p1_l[57]), 
        .p2m1_l(p2_l[57]) );
  mul_ppgen3_54 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .p2_l(p2_l[57]), .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[56]), .p1m1_l(p1_l[56]), 
        .p2m1_l(p2_l[56]) );
  mul_ppgen3_53 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .p2_l(p2_l[56]), .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[55]), .p1m1_l(p1_l[55]), 
        .p2m1_l(p2_l[55]) );
  mul_ppgen3_52 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .p2_l(p2_l[55]), .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[54]), .p1m1_l(p1_l[54]), 
        .p2m1_l(p2_l[54]) );
  mul_ppgen3_51 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .p2_l(p2_l[54]), .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[53]), .p1m1_l(p1_l[53]), 
        .p2m1_l(p2_l[53]) );
  mul_ppgen3_50 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .p2_l(p2_l[53]), .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[52]), .p1m1_l(p1_l[52]), 
        .p2m1_l(p2_l[52]) );
  mul_ppgen3_49 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .p2_l(p2_l[52]), .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[51]), .p1m1_l(p1_l[51]), 
        .p2m1_l(p2_l[51]) );
  mul_ppgen3_48 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .p2_l(p2_l[51]), .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[50]), .p1m1_l(p1_l[50]), 
        .p2m1_l(p2_l[50]) );
  mul_ppgen3_47 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .p2_l(p2_l[50]), .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[49]), .p1m1_l(p1_l[49]), 
        .p2m1_l(p2_l[49]) );
  mul_ppgen3_46 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .p2_l(p2_l[49]), .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[48]), .p1m1_l(p1_l[48]), 
        .p2m1_l(p2_l[48]) );
  mul_ppgen3_45 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .p2_l(p2_l[48]), .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[47]), .p1m1_l(p1_l[47]), 
        .p2m1_l(p2_l[47]) );
  mul_ppgen3_44 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .p2_l(p2_l[47]), .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[46]), .p1m1_l(p1_l[46]), 
        .p2m1_l(p2_l[46]) );
  mul_ppgen3_43 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .p2_l(p2_l[46]), .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[45]), .p1m1_l(p1_l[45]), 
        .p2m1_l(p2_l[45]) );
  mul_ppgen3_42 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .p2_l(p2_l[45]), .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[44]), .p1m1_l(p1_l[44]), 
        .p2m1_l(p2_l[44]) );
  mul_ppgen3_41 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .p2_l(p2_l[44]), .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[43]), .p1m1_l(p1_l[43]), 
        .p2m1_l(p2_l[43]) );
  mul_ppgen3_40 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .p2_l(p2_l[43]), .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[42]), .p1m1_l(p1_l[42]), 
        .p2m1_l(p2_l[42]) );
  mul_ppgen3_39 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .p2_l(p2_l[42]), .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[41]), .p1m1_l(p1_l[41]), 
        .p2m1_l(p2_l[41]) );
  mul_ppgen3_38 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .p2_l(p2_l[41]), .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[40]), .p1m1_l(p1_l[40]), 
        .p2m1_l(p2_l[40]) );
  mul_ppgen3_37 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .p2_l(p2_l[40]), .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[39]), .p1m1_l(p1_l[39]), 
        .p2m1_l(p2_l[39]) );
  mul_ppgen3_36 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .p2_l(p2_l[39]), .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[38]), .p1m1_l(p1_l[38]), 
        .p2m1_l(p2_l[38]) );
  mul_ppgen3_35 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .p2_l(p2_l[38]), .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[37]), .p1m1_l(p1_l[37]), 
        .p2m1_l(p2_l[37]) );
  mul_ppgen3_34 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .p2_l(p2_l[37]), .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[36]), .p1m1_l(p1_l[36]), 
        .p2m1_l(p2_l[36]) );
  mul_ppgen3_33 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .p2_l(p2_l[36]), .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[35]), .p1m1_l(p1_l[35]), 
        .p2m1_l(p2_l[35]) );
  mul_ppgen3_32 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .p2_l(p2_l[35]), .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[34]), .p1m1_l(p1_l[34]), 
        .p2m1_l(p2_l[34]) );
  mul_ppgen3_31 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .p2_l(p2_l[34]), .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[33]), .p1m1_l(p1_l[33]), 
        .p2m1_l(p2_l[33]) );
  mul_ppgen3_30 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .p2_l(p2_l[33]), .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[32]), .p1m1_l(p1_l[32]), 
        .p2m1_l(p2_l[32]) );
  mul_ppgen3_29 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .p2_l(p2_l[32]), .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[31]), .p1m1_l(p1_l[31]), 
        .p2m1_l(p2_l[31]) );
  mul_ppgen3_28 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .p2_l(p2_l[31]), .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[30]), .p1m1_l(p1_l[30]), 
        .p2m1_l(p2_l[30]) );
  mul_ppgen3_27 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .p2_l(p2_l[30]), .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[29]), .p1m1_l(p1_l[29]), 
        .p2m1_l(p2_l[29]) );
  mul_ppgen3_26 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .p2_l(p2_l[29]), .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[28]), .p1m1_l(p1_l[28]), 
        .p2m1_l(p2_l[28]) );
  mul_ppgen3_25 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .p2_l(p2_l[28]), .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[27]), .p1m1_l(p1_l[27]), 
        .p2m1_l(p2_l[27]) );
  mul_ppgen3_24 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .p2_l(p2_l[27]), .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[26]), .p1m1_l(p1_l[26]), 
        .p2m1_l(p2_l[26]) );
  mul_ppgen3_23 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .p2_l(p2_l[26]), .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[25]), .p1m1_l(p1_l[25]), 
        .p2m1_l(p2_l[25]) );
  mul_ppgen3_22 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .p2_l(p2_l[25]), .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[24]), .p1m1_l(p1_l[24]), 
        .p2m1_l(p2_l[24]) );
  mul_ppgen3_21 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .p2_l(p2_l[24]), .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[23]), .p1m1_l(p1_l[23]), 
        .p2m1_l(p2_l[23]) );
  mul_ppgen3_20 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .p2_l(p2_l[23]), .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[22]), .p1m1_l(p1_l[22]), 
        .p2m1_l(p2_l[22]) );
  mul_ppgen3_19 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .p2_l(p2_l[22]), .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[21]), .p1m1_l(p1_l[21]), 
        .p2m1_l(p2_l[21]) );
  mul_ppgen3_18 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .p2_l(p2_l[21]), .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[20]), .p1m1_l(p1_l[20]), 
        .p2m1_l(p2_l[20]) );
  mul_ppgen3_17 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .p2_l(p2_l[20]), .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[19]), .p1m1_l(p1_l[19]), 
        .p2m1_l(p2_l[19]) );
  mul_ppgen3_16 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .p2_l(p2_l[19]), .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[18]), .p1m1_l(p1_l[18]), 
        .p2m1_l(p2_l[18]) );
  mul_ppgen3_15 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .p2_l(p2_l[18]), .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[17]), .p1m1_l(p1_l[17]), 
        .p2m1_l(p2_l[17]) );
  mul_ppgen3_14 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .p2_l(p2_l[17]), .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[16]), .p1m1_l(p1_l[16]), 
        .p2m1_l(p2_l[16]) );
  mul_ppgen3_13 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .p2_l(p2_l[16]), .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[15]), .p1m1_l(p1_l[15]), 
        .p2m1_l(p2_l[15]) );
  mul_ppgen3_12 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .p2_l(p2_l[15]), .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[14]), .p1m1_l(p1_l[14]), 
        .p2m1_l(p2_l[14]) );
  mul_ppgen3_11 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .p2_l(p2_l[14]), .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[13]), .p1m1_l(p1_l[13]), 
        .p2m1_l(p2_l[13]) );
  mul_ppgen3_10 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .p2_l(p2_l[13]), .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[12]), .p1m1_l(p1_l[12]), 
        .p2m1_l(p2_l[12]) );
  mul_ppgen3_9 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .p2_l(p2_l[12]), .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[11]), .p1m1_l(p1_l[11]), 
        .p2m1_l(p2_l[11]) );
  mul_ppgen3_8 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .p2_l(p2_l[11]), .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[10]), .p1m1_l(p1_l[10]), 
        .p2m1_l(p2_l[10]) );
  mul_ppgen3_7 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .p2_l(p2_l[10]), .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[9]), .p1m1_l(p1_l[9]), 
        .p2m1_l(p2_l[9]) );
  mul_ppgen3_6 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), .p2_l(
        p2_l[9]), .sum(sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), .p2m1_l(p2_l[8])
         );
  mul_ppgen3_5 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), .p2_l(
        p2_l[8]), .sum(sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), .p2m1_l(p2_l[7])
         );
  mul_ppgen3_4 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), .p2_l(
        p2_l[7]), .sum(sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), .p2m1_l(p2_l[6])
         );
  mul_ppgen3_3 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), .p2_l(
        p2_l[6]), .sum(sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), .p2m1_l(p2_l[5])
         );
  mul_ppgen3_2 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), .p2_l(
        p2_l[5]), .sum(sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), .p2m1_l(p2_l[4])
         );
  mul_ppgen3_1 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), .p2_l(
        p2_l[4]), .sum(sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), .p2m1_l(1'b1) );
  mul_ppgen3lsb4_1 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ppgen_379 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_380 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_381 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_382 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_383 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_384 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_4 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_csa32_129 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_130 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_131 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  OR2X1_RVT U1 ( .A1(a), .A2(c), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(a), .A2(c), .Y(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(cout), .Y(sum) );
endmodule


module mul_csa32_132 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(c), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ppgensign_4 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_5 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_6 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_2 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net42, net47, p2_l_67, net073, p1_l_65, net38, net0118, p2_l_66,
         net078, p2_l_65, net8, p2_l_64, net15, p1_l_64, net43, net48, net35;

  mul_ppgensign_6 p0_64_ ( .p_l(net42), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_5 p2_68_ ( .p_l(sum[5]), .z(net073), .b(b2), .pm1_l(p2_l_67)
         );
  mul_ppgensign_4 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ha_4 sc1_68_ ( .cout(cout[4]), .sum(sum[4]), .a(1'b1), .b(net073) );
  mul_ppgen_384 p2_67_ ( .p_l(p2_l_67), .z(net078), .a(am1), .b(b2), .pm1_l(
        p2_l_66) );
  mul_ppgen_383 p2_66_ ( .p_l(p2_l_66), .z(net8), .a(am2), .b(b2), .pm1_l(
        p2_l_65) );
  mul_ppgen_382 p2_65_ ( .p_l(p2_l_65), .z(net15), .a(am3), .b(b2), .pm1_l(
        p2_l_64) );
  mul_ppgen_381 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_380 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_ppgen_379 p2_64_ ( .p_l(p2_l_64), .z(net35), .a(am4), .b(b2), .pm1_l(
        p2m1_l) );
  mul_csa32_132 sc1_67_ ( .sum(sum[3]), .cout(cout[3]), .a(net0118), .b(1'b0), 
        .c(net078) );
  mul_csa32_131 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(1'b1), 
        .c(net8) );
  mul_csa32_130 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net15) );
  mul_csa32_129 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net35) );
endmodule


module mul_ppgen_193 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_194 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_195 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_196 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_197 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_198 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_3 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_3 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_4 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_67 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_68 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_2 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_4 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_3 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_68 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_67 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_3 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_198 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_197 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_196 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(
        p0_l_1) );
  mul_ppgen_195 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(
        p0_l_0) );
  mul_ppgen_194 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_193 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_199 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_200 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_201 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_csa32_69 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_61 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043, net210262;

  mul_csa32_69 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_201 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(net210262) );
  mul_ppgen_200 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_199 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_202 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_203 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_204 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_70 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_62 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_70 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_204 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_203 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_202 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_205 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_206 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_207 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_71 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_63 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_71 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_207 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_206 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_205 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_208 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_209 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_210 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_72 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_64 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_72 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_210 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_209 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_208 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_211 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_212 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_213 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_73 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_65 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_73 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_213 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_212 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_211 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_214 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_215 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_216 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_74 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_66 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_74 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_216 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_215 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_214 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_217 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_218 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_219 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_75 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_67 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_75 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_219 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_218 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_217 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_220 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_221 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_222 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_76 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_68 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_76 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_222 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_221 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_220 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_223 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_224 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_225 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_77 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_69 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_77 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_225 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_224 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_223 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_226 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_227 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_228 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_78 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_70 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_78 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_228 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_227 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_226 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_229 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_230 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_231 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_79 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_71 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_79 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_231 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_230 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_229 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_232 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_233 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_234 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_80 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_72 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_80 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_234 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_233 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_232 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_235 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_236 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_237 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_81 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_73 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_81 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_237 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_236 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_235 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_238 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_239 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_240 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_82 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_74 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_82 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_240 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_239 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_238 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_241 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_242 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_243 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_83 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_75 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_83 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_243 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_242 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_241 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_244 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_245 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_246 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_84 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_76 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_84 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_246 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_245 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_244 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_247 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_248 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_249 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_85 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_77 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_85 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_249 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_248 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_247 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_250 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_251 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_252 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_86 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_78 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_86 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_252 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_251 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_250 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_253 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_254 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_255 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_87 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_79 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_87 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_255 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_254 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_253 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_256 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_257 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_258 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_88 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_80 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_88 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_258 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_257 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_256 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_259 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_260 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_261 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_89 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_81 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_89 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_261 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_260 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_259 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_262 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_263 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_264 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_90 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_82 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_90 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_264 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_263 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_262 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_265 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_266 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_267 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_91 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_83 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_91 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_267 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_266 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_265 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_268 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_269 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_270 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_92 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_84 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_92 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_270 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_269 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_268 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_271 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_272 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_273 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_93 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_85 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_93 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_273 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_272 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_271 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_274 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_275 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_276 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_94 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_86 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_94 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_276 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_275 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_274 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_277 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_278 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_279 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_95 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_87 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_95 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_279 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_278 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_277 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_280 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_281 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_282 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_96 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_88 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_96 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_282 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_281 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_280 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_283 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_284 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_285 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_97 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_89 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_97 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_285 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_284 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_283 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_286 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_287 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_288 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_98 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_90 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_98 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_288 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_287 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_286 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_289 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_290 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_291 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_99 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_91 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_99 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043)
         );
  mul_ppgen_291 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_290 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_289 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_292 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_293 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_294 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_100 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_92 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_100 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_294 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_293 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_292 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_295 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_296 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_297 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_101 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_93 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_101 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_297 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_296 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_295 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_298 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_299 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_300 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_102 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_94 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_102 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_300 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_299 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_298 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_301 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_302 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_303 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_103 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_95 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_103 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_303 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_302 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_301 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_304 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_305 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_306 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_104 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_96 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_104 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_306 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_305 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_304 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_307 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_308 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_309 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_105 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_97 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_105 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_309 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_308 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_307 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_310 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_311 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_312 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_106 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_98 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_106 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_312 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_311 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_310 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_313 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_314 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_315 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_107 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_99 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_107 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_315 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_314 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_313 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_316 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_317 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_318 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_108 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_100 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_108 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_318 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_317 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_316 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_319 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_320 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_321 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_109 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_101 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_109 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_321 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_320 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_319 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_322 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_323 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_324 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_110 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_102 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_110 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_324 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_323 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_322 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_325 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_326 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_327 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_111 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_103 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_111 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_327 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_326 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_325 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_328 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_329 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_330 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_112 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_104 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_112 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_330 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_329 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_328 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_331 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_332 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_333 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_113 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_105 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_113 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_333 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_332 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_331 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_334 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_335 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_336 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_114 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_106 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_114 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_336 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_335 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_334 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_337 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_338 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_339 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_115 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_107 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_115 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_339 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_338 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_337 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_340 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_341 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_342 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_116 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_108 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_116 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_342 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_341 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_340 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_343 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_344 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_345 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_117 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_109 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_117 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_345 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_344 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_343 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_346 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_347 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_348 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_118 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_110 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_118 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_348 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_347 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_346 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_349 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_350 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_351 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_119 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_111 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_119 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_351 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_350 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_349 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_352 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_353 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_354 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_120 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_112 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_120 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_354 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_353 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_352 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_355 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_356 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_357 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_121 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_113 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_121 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_357 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_356 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_355 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_358 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_359 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_360 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_122 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_114 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_122 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_360 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_359 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_358 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_361 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_362 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_363 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_123 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_115 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_123 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_363 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_362 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_361 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_364 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_365 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_366 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_124 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_116 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_124 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_366 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_365 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_364 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_367 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_368 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_369 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_125 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_117 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_125 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_369 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_368 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_367 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_370 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_371 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_372 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_126 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_118 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_126 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_372 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_371 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_370 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_373 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_374 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_375 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_127 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_119 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_127 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_375 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_374 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_373 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_376 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_377 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_378 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_128 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3_120 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32_128 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen_378 p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_ppgen_377 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_376 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_2 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210524, net210525;
  wire   [63:4] p2_l;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;

  mul_ppgen3sign_2 I2 ( .cout(cout[68:64]), .sum(sum[69:64]), .am1(a[63]), 
        .am2(a[62]), .am3(a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2(b2), 
        .bot(net210524), .head(net210525), .p0m1_l(p0_l[63]), .p1m1_l(p1_l[63]), .p2m1_l(p2_l[63]) );
  mul_ppgen3_120 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .p2_l(p2_l[63]), .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[62]), .p1m1_l(p1_l[62]), 
        .p2m1_l(p2_l[62]) );
  mul_ppgen3_119 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .p2_l(p2_l[62]), .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[61]), .p1m1_l(p1_l[61]), 
        .p2m1_l(p2_l[61]) );
  mul_ppgen3_118 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .p2_l(p2_l[61]), .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[60]), .p1m1_l(p1_l[60]), 
        .p2m1_l(p2_l[60]) );
  mul_ppgen3_117 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .p2_l(p2_l[60]), .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[59]), .p1m1_l(p1_l[59]), 
        .p2m1_l(p2_l[59]) );
  mul_ppgen3_116 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .p2_l(p2_l[59]), .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[58]), .p1m1_l(p1_l[58]), 
        .p2m1_l(p2_l[58]) );
  mul_ppgen3_115 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .p2_l(p2_l[58]), .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[57]), .p1m1_l(p1_l[57]), 
        .p2m1_l(p2_l[57]) );
  mul_ppgen3_114 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .p2_l(p2_l[57]), .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[56]), .p1m1_l(p1_l[56]), 
        .p2m1_l(p2_l[56]) );
  mul_ppgen3_113 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .p2_l(p2_l[56]), .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[55]), .p1m1_l(p1_l[55]), 
        .p2m1_l(p2_l[55]) );
  mul_ppgen3_112 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .p2_l(p2_l[55]), .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[54]), .p1m1_l(p1_l[54]), 
        .p2m1_l(p2_l[54]) );
  mul_ppgen3_111 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .p2_l(p2_l[54]), .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[53]), .p1m1_l(p1_l[53]), 
        .p2m1_l(p2_l[53]) );
  mul_ppgen3_110 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .p2_l(p2_l[53]), .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[52]), .p1m1_l(p1_l[52]), 
        .p2m1_l(p2_l[52]) );
  mul_ppgen3_109 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .p2_l(p2_l[52]), .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[51]), .p1m1_l(p1_l[51]), 
        .p2m1_l(p2_l[51]) );
  mul_ppgen3_108 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .p2_l(p2_l[51]), .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[50]), .p1m1_l(p1_l[50]), 
        .p2m1_l(p2_l[50]) );
  mul_ppgen3_107 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .p2_l(p2_l[50]), .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[49]), .p1m1_l(p1_l[49]), 
        .p2m1_l(p2_l[49]) );
  mul_ppgen3_106 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .p2_l(p2_l[49]), .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[48]), .p1m1_l(p1_l[48]), 
        .p2m1_l(p2_l[48]) );
  mul_ppgen3_105 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .p2_l(p2_l[48]), .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[47]), .p1m1_l(p1_l[47]), 
        .p2m1_l(p2_l[47]) );
  mul_ppgen3_104 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .p2_l(p2_l[47]), .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[46]), .p1m1_l(p1_l[46]), 
        .p2m1_l(p2_l[46]) );
  mul_ppgen3_103 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .p2_l(p2_l[46]), .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[45]), .p1m1_l(p1_l[45]), 
        .p2m1_l(p2_l[45]) );
  mul_ppgen3_102 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .p2_l(p2_l[45]), .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[44]), .p1m1_l(p1_l[44]), 
        .p2m1_l(p2_l[44]) );
  mul_ppgen3_101 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .p2_l(p2_l[44]), .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[43]), .p1m1_l(p1_l[43]), 
        .p2m1_l(p2_l[43]) );
  mul_ppgen3_100 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .p2_l(p2_l[43]), .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[42]), .p1m1_l(p1_l[42]), 
        .p2m1_l(p2_l[42]) );
  mul_ppgen3_99 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .p2_l(p2_l[42]), .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[41]), .p1m1_l(p1_l[41]), 
        .p2m1_l(p2_l[41]) );
  mul_ppgen3_98 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .p2_l(p2_l[41]), .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[40]), .p1m1_l(p1_l[40]), 
        .p2m1_l(p2_l[40]) );
  mul_ppgen3_97 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .p2_l(p2_l[40]), .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[39]), .p1m1_l(p1_l[39]), 
        .p2m1_l(p2_l[39]) );
  mul_ppgen3_96 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .p2_l(p2_l[39]), .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[38]), .p1m1_l(p1_l[38]), 
        .p2m1_l(p2_l[38]) );
  mul_ppgen3_95 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .p2_l(p2_l[38]), .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[37]), .p1m1_l(p1_l[37]), 
        .p2m1_l(p2_l[37]) );
  mul_ppgen3_94 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .p2_l(p2_l[37]), .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[36]), .p1m1_l(p1_l[36]), 
        .p2m1_l(p2_l[36]) );
  mul_ppgen3_93 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .p2_l(p2_l[36]), .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[35]), .p1m1_l(p1_l[35]), 
        .p2m1_l(p2_l[35]) );
  mul_ppgen3_92 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .p2_l(p2_l[35]), .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[34]), .p1m1_l(p1_l[34]), 
        .p2m1_l(p2_l[34]) );
  mul_ppgen3_91 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .p2_l(p2_l[34]), .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[33]), .p1m1_l(p1_l[33]), 
        .p2m1_l(p2_l[33]) );
  mul_ppgen3_90 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .p2_l(p2_l[33]), .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[32]), .p1m1_l(p1_l[32]), 
        .p2m1_l(p2_l[32]) );
  mul_ppgen3_89 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .p2_l(p2_l[32]), .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[31]), .p1m1_l(p1_l[31]), 
        .p2m1_l(p2_l[31]) );
  mul_ppgen3_88 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .p2_l(p2_l[31]), .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[30]), .p1m1_l(p1_l[30]), 
        .p2m1_l(p2_l[30]) );
  mul_ppgen3_87 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .p2_l(p2_l[30]), .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[29]), .p1m1_l(p1_l[29]), 
        .p2m1_l(p2_l[29]) );
  mul_ppgen3_86 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .p2_l(p2_l[29]), .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[28]), .p1m1_l(p1_l[28]), 
        .p2m1_l(p2_l[28]) );
  mul_ppgen3_85 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .p2_l(p2_l[28]), .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[27]), .p1m1_l(p1_l[27]), 
        .p2m1_l(p2_l[27]) );
  mul_ppgen3_84 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .p2_l(p2_l[27]), .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[26]), .p1m1_l(p1_l[26]), 
        .p2m1_l(p2_l[26]) );
  mul_ppgen3_83 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .p2_l(p2_l[26]), .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[25]), .p1m1_l(p1_l[25]), 
        .p2m1_l(p2_l[25]) );
  mul_ppgen3_82 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .p2_l(p2_l[25]), .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[24]), .p1m1_l(p1_l[24]), 
        .p2m1_l(p2_l[24]) );
  mul_ppgen3_81 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .p2_l(p2_l[24]), .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[23]), .p1m1_l(p1_l[23]), 
        .p2m1_l(p2_l[23]) );
  mul_ppgen3_80 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .p2_l(p2_l[23]), .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[22]), .p1m1_l(p1_l[22]), 
        .p2m1_l(p2_l[22]) );
  mul_ppgen3_79 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .p2_l(p2_l[22]), .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[21]), .p1m1_l(p1_l[21]), 
        .p2m1_l(p2_l[21]) );
  mul_ppgen3_78 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .p2_l(p2_l[21]), .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[20]), .p1m1_l(p1_l[20]), 
        .p2m1_l(p2_l[20]) );
  mul_ppgen3_77 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .p2_l(p2_l[20]), .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[19]), .p1m1_l(p1_l[19]), 
        .p2m1_l(p2_l[19]) );
  mul_ppgen3_76 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .p2_l(p2_l[19]), .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[18]), .p1m1_l(p1_l[18]), 
        .p2m1_l(p2_l[18]) );
  mul_ppgen3_75 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .p2_l(p2_l[18]), .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[17]), .p1m1_l(p1_l[17]), 
        .p2m1_l(p2_l[17]) );
  mul_ppgen3_74 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .p2_l(p2_l[17]), .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[16]), .p1m1_l(p1_l[16]), 
        .p2m1_l(p2_l[16]) );
  mul_ppgen3_73 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .p2_l(p2_l[16]), .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[15]), .p1m1_l(p1_l[15]), 
        .p2m1_l(p2_l[15]) );
  mul_ppgen3_72 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .p2_l(p2_l[15]), .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[14]), .p1m1_l(p1_l[14]), 
        .p2m1_l(p2_l[14]) );
  mul_ppgen3_71 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .p2_l(p2_l[14]), .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[13]), .p1m1_l(p1_l[13]), 
        .p2m1_l(p2_l[13]) );
  mul_ppgen3_70 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .p2_l(p2_l[13]), .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[12]), .p1m1_l(p1_l[12]), 
        .p2m1_l(p2_l[12]) );
  mul_ppgen3_69 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .p2_l(p2_l[12]), .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[11]), .p1m1_l(p1_l[11]), 
        .p2m1_l(p2_l[11]) );
  mul_ppgen3_68 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .p2_l(p2_l[11]), .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[10]), .p1m1_l(p1_l[10]), 
        .p2m1_l(p2_l[10]) );
  mul_ppgen3_67 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .p2_l(p2_l[10]), .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[9]), .p1m1_l(p1_l[9]), 
        .p2m1_l(p2_l[9]) );
  mul_ppgen3_66 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), .p2_l(
        p2_l[9]), .sum(sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), .p2m1_l(p2_l[8])
         );
  mul_ppgen3_65 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), .p2_l(
        p2_l[8]), .sum(sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), .p2m1_l(p2_l[7])
         );
  mul_ppgen3_64 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), .p2_l(
        p2_l[7]), .sum(sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), .p2m1_l(p2_l[6])
         );
  mul_ppgen3_63 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), .p2_l(
        p2_l[6]), .sum(sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), .p2m1_l(p2_l[5])
         );
  mul_ppgen3_62 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), .p2_l(
        p2_l[5]), .sum(sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), .p2m1_l(p2_l[4])
         );
  mul_ppgen3_61 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), .p2_l(
        p2_l[4]), .sum(sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), .p2m1_l(1'b1) );
  mul_ppgen3lsb4_2 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ppgen_572 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_573 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_195 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_196 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_csa32_197 ( sum, cout, a, b, c_BAR );
  input a, b, c_BAR;
  output sum, cout;
  wire   a;
  assign cout = a;

  INVX1_RVT U1 ( .A(a), .Y(sum) );
endmodule


module mul_csa32_198 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   a;
  assign sum = a;

endmodule


module mul_ppgensign_7 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgensign_9 ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   n1;

  INVX0_RVT U1 ( .A(b[0]), .Y(n1) );
  NAND2X0_RVT U2 ( .A1(b[2]), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U3 ( .A1(b[0]), .A2(pm1_l), .A3(n1), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen3sign_3 ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   bot, net42, net47, p1_l_65, net38, net0118, p1_l_64, net43, net48,
         net210273, net210274, net210275, net210276;
  assign sum[5] = bot;

  mul_ppgensign_9 p0_64_ ( .p_l(net42), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign_7 p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65)
         );
  mul_ppgen_573 p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(
        p1_l_64) );
  mul_ppgen_572 p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(
        p1m1_l) );
  mul_csa32_198 sc1_67_ ( .sum(sum[3]), .a(net0118), .b(1'b0), .c(net210276)
         );
  mul_csa32_197 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(1'b1), 
        .c_BAR(net210275) );
  mul_csa32_196 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), 
        .c(net210274) );
  mul_csa32_195 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), 
        .c(net210273) );
endmodule


module mul_ppgen_385 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_386 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1;

  HADDX1_RVT U1 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U2 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  NOR2X0_RVT U3 ( .A1(b[0]), .A2(p_l), .Y(z) );
endmodule


module mul_ppgen_387 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_388 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_389 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_390 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ha_5 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_5 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_6 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
  AND3X1_RVT U3 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
endmodule


module mul_csa32_133 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_134 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_ppgen3lsb4_3 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0;

  mul_negen_6 p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen_5 p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32_134 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32_133 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha_5 sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen_390 p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2)
         );
  mul_ppgen_389 p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2)
         );
  mul_ppgen_388 p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(
        p0_l_1) );
  mul_ppgen_387 p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(
        p0_l_0) );
  mul_ppgen_386 p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1)
         );
  mul_ppgen_385 p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1)
         );
  AO21X1_RVT U3 ( .A1(p0_0), .A2(b0n_0), .A3(b0n_1), .Y(b0n) );
  HADDX1_RVT U4 ( .A0(b0n_0), .B0(p0_0), .SO(sum[0]) );
endmodule


module mul_ppgen_391 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_392 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_135 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_121 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210261;

  mul_csa32_135 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210261) );
  mul_ppgen_392 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_391 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_394 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_395 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_136 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_122 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210260;

  mul_csa32_136 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210260) );
  mul_ppgen_395 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_394 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_397 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_398 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_137 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_123 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210259;

  mul_csa32_137 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210259) );
  mul_ppgen_398 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_397 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_400 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_401 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_138 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_124 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210258;

  mul_csa32_138 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210258) );
  mul_ppgen_401 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_400 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_403 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_404 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_139 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_125 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210257;

  mul_csa32_139 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210257) );
  mul_ppgen_404 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_403 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_406 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_407 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_140 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_126 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210256;

  mul_csa32_140 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210256) );
  mul_ppgen_407 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_406 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_409 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_410 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_141 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_127 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210255;

  mul_csa32_141 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210255) );
  mul_ppgen_410 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_409 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_412 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_413 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_142 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_128 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210254;

  mul_csa32_142 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210254) );
  mul_ppgen_413 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_412 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_415 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_416 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_143 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_129 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210253;

  mul_csa32_143 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210253) );
  mul_ppgen_416 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_415 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_418 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_419 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_144 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_130 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210252;

  mul_csa32_144 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210252) );
  mul_ppgen_419 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_418 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_421 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_422 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_145 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_131 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210251;

  mul_csa32_145 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210251) );
  mul_ppgen_422 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_421 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_424 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_425 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_146 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_132 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210250;

  mul_csa32_146 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210250) );
  mul_ppgen_425 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_424 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_427 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_428 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_147 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_133 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210249;

  mul_csa32_147 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210249) );
  mul_ppgen_428 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_427 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_430 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_431 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_148 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_134 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210248;

  mul_csa32_148 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210248) );
  mul_ppgen_431 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_430 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_433 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_434 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_149 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_135 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210247;

  mul_csa32_149 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210247) );
  mul_ppgen_434 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_433 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_436 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_437 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_150 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_136 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210246;

  mul_csa32_150 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210246) );
  mul_ppgen_437 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_436 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_439 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_440 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_151 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_137 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210245;

  mul_csa32_151 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210245) );
  mul_ppgen_440 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_439 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_442 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_443 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_152 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_138 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210244;

  mul_csa32_152 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210244) );
  mul_ppgen_443 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_442 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_445 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_446 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_153 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_139 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210243;

  mul_csa32_153 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210243) );
  mul_ppgen_446 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_445 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_448 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_449 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_154 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_140 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210242;

  mul_csa32_154 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210242) );
  mul_ppgen_449 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_448 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_451 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_452 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_155 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_141 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210241;

  mul_csa32_155 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210241) );
  mul_ppgen_452 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_451 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_454 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_455 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_156 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_142 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210240;

  mul_csa32_156 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210240) );
  mul_ppgen_455 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_454 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_457 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_458 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_157 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_143 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210239;

  mul_csa32_157 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210239) );
  mul_ppgen_458 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_457 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_460 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_461 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_158 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_144 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210238;

  mul_csa32_158 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210238) );
  mul_ppgen_461 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_460 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_463 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_464 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_159 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_145 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210237;

  mul_csa32_159 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210237) );
  mul_ppgen_464 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_463 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_466 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_467 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_160 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_146 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210236;

  mul_csa32_160 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210236) );
  mul_ppgen_467 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_466 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_469 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_470 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_161 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_147 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210235;

  mul_csa32_161 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210235) );
  mul_ppgen_470 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_469 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_472 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_473 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_162 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_148 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210234;

  mul_csa32_162 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210234) );
  mul_ppgen_473 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_472 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_475 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_476 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_163 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_149 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210233;

  mul_csa32_163 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210233) );
  mul_ppgen_476 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_475 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_478 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_479 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_164 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_150 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210232;

  mul_csa32_164 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210232) );
  mul_ppgen_479 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_478 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_481 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_482 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_165 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_151 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210231;

  mul_csa32_165 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210231) );
  mul_ppgen_482 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_481 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_484 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_485 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_166 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_152 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210230;

  mul_csa32_166 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210230) );
  mul_ppgen_485 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_484 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_487 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_488 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_167 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_153 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210229;

  mul_csa32_167 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210229) );
  mul_ppgen_488 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_487 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_490 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_491 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_168 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_154 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210228;

  mul_csa32_168 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210228) );
  mul_ppgen_491 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_490 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_493 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_494 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_169 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_155 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210227;

  mul_csa32_169 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210227) );
  mul_ppgen_494 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_493 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_496 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_497 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_170 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_156 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210226;

  mul_csa32_170 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210226) );
  mul_ppgen_497 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_496 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_499 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_500 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_171 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_157 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210225;

  mul_csa32_171 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210225) );
  mul_ppgen_500 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_499 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_502 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_503 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_172 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_158 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210224;

  mul_csa32_172 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210224) );
  mul_ppgen_503 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_502 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_505 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_506 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_173 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_159 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210223;

  mul_csa32_173 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210223) );
  mul_ppgen_506 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_505 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_508 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_509 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_174 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_160 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210222;

  mul_csa32_174 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210222) );
  mul_ppgen_509 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_508 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_511 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_512 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_175 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_161 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210221;

  mul_csa32_175 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210221) );
  mul_ppgen_512 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_511 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_514 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_515 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_176 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_162 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210220;

  mul_csa32_176 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210220) );
  mul_ppgen_515 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_514 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_517 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_518 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_177 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_163 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210219;

  mul_csa32_177 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210219) );
  mul_ppgen_518 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_517 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_520 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_521 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_178 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_164 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210218;

  mul_csa32_178 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210218) );
  mul_ppgen_521 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_520 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_523 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_524 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_179 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_165 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210217;

  mul_csa32_179 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210217) );
  mul_ppgen_524 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_523 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_526 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_527 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_180 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_166 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210216;

  mul_csa32_180 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210216) );
  mul_ppgen_527 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_526 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_529 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_530 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_181 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_167 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210215;

  mul_csa32_181 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210215) );
  mul_ppgen_530 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_529 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_532 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_533 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_182 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_168 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210214;

  mul_csa32_182 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210214) );
  mul_ppgen_533 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_532 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_535 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_536 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_183 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_169 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210213;

  mul_csa32_183 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210213) );
  mul_ppgen_536 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_535 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_538 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_539 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_184 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_170 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210212;

  mul_csa32_184 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210212) );
  mul_ppgen_539 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_538 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_541 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_542 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_185 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_171 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210211;

  mul_csa32_185 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210211) );
  mul_ppgen_542 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_541 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_544 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_545 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_186 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_172 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210210;

  mul_csa32_186 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210210) );
  mul_ppgen_545 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_544 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_547 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_548 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_187 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_173 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210209;

  mul_csa32_187 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210209) );
  mul_ppgen_548 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_547 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_550 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_551 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_188 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_174 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210208;

  mul_csa32_188 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210208) );
  mul_ppgen_551 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_550 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_553 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_554 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_189 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_175 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210207;

  mul_csa32_189 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210207) );
  mul_ppgen_554 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_553 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_556 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_557 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_190 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_176 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210206;

  mul_csa32_190 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210206) );
  mul_ppgen_557 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_556 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_559 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_560 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_191 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_177 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210205;

  mul_csa32_191 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210205) );
  mul_ppgen_560 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_559 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_562 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_563 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_192 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_178 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210204;

  mul_csa32_192 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210204) );
  mul_ppgen_563 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_562 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_565 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_566 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_193 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_179 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210203;

  mul_csa32_193 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210203) );
  mul_ppgen_566 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_565 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen_568 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_ppgen_569 ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  HADDX1_RVT U2 ( .A0(a), .B0(b[2]), .SO(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(b[1]), .Y(p_l) );
  AOI22X1_RVT U4 ( .A1(b[0]), .A2(pm1_l), .A3(n2), .A4(p_l), .Y(z) );
endmodule


module mul_csa32_194 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(a), .A2(b), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(a), .A2(b), .A3(n1), .Y(sum) );
endmodule


module mul_ppgen3_180 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net210202;

  mul_csa32_194 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(
        net210202) );
  mul_ppgen_569 p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen_568 p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgenrow3_3 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;
  wire   net210280, net210281, net210282, net210283, net210284, net210285,
         net210286, net210287, net210288, net210289, net210290, net210291,
         net210292, net210293, net210294, net210295, net210296, net210297,
         net210298, net210299, net210300, net210301, net210302, net210303,
         net210304, net210305, net210306, net210307, net210308, net210309,
         net210310, net210311, net210312, net210313, net210314, net210315,
         net210316, net210317, net210318, net210319, net210320, net210321,
         net210322, net210323, net210324, net210325, net210326, net210327,
         net210328, net210329, net210330, net210331, net210332, net210333,
         net210334, net210335, net210336, net210337, net210338, net210339,
         net210340, net210341, net210342, net210343, net210344, net210345,
         net210346, net210347, net210348, net210349, net210350, net210351,
         net210352, net210353, net210354, net210355, net210356, net210357,
         net210358, net210359, net210360, net210361, net210362, net210363,
         net210364, net210365, net210366, net210367, net210368, net210369,
         net210370, net210371, net210372, net210373, net210374, net210375,
         net210376, net210377, net210378, net210379, net210380, net210381,
         net210382, net210383, net210384, net210385, net210386, net210387,
         net210388, net210389, net210390, net210391, net210392, net210393,
         net210394, net210395, net210396, net210397, net210398, net210399,
         net210400, net210401, net210402, net210403, net210404, net210405,
         net210406, net210407, net210408, net210409, net210410, net210411,
         net210412, net210413, net210414, net210415, net210416, net210417,
         net210418, net210419, net210420, net210421, net210422, net210423,
         net210424, net210425, net210426, net210427, net210428, net210429,
         net210430, net210431, net210432, net210433, net210434, net210435,
         net210436, net210437, net210438, net210439, net210440, net210441,
         net210442, net210443, net210444, net210445, net210446, net210447,
         net210448, net210449, net210450, net210451, net210452, net210453,
         net210454, net210455, net210456, net210457, net210458, net210459,
         net210460, net210461, net210462, net210463, net210464, net210465,
         net210466, net210467, net210468, net210469, net210470, net210471,
         net210472, net210473, net210474, net210475, net210476, net210477,
         net210478, net210479, net210480, net210481, net210482, net210483,
         net210484, net210485, net210486, net210487, net210488, net210489,
         net210490, net210491, net210492, net210493, net210494, net210495,
         net210496, net210497, net210498, net210499, net210500, net210501,
         net210502, net210503, net210504, net210505, net210506, net210507,
         net210508, net210509, net210510, net210511, net210512, net210513,
         net210514, net210515, net210516, net210517, net210518, net210519,
         net210520, net210521, net210522, net210523;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  mul_ppgen3sign_3 I2 ( .cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, cout[66:64]}), .sum({sum[69], 
        SYNOPSYS_UNCONNECTED__2, sum[67:64]}), .am1(a[63]), .am2(a[62]), .am3(
        a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2({net210519, net210520, 
        net210521}), .bot(bot), .head(net210522), .p0m1_l(p0_l[63]), .p1m1_l(
        p1_l[63]), .p2m1_l(net210523) );
  mul_ppgen3_180 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), .b0(b0), .b1(b1), 
        .b2({net210515, net210516, net210517}), .p0m1_l(p0_l[62]), .p1m1_l(
        p1_l[62]), .p2m1_l(net210518) );
  mul_ppgen3_179 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), .b0(b0), .b1(b1), 
        .b2({net210511, net210512, net210513}), .p0m1_l(p0_l[61]), .p1m1_l(
        p1_l[61]), .p2m1_l(net210514) );
  mul_ppgen3_178 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), .b0(b0), .b1(b1), 
        .b2({net210507, net210508, net210509}), .p0m1_l(p0_l[60]), .p1m1_l(
        p1_l[60]), .p2m1_l(net210510) );
  mul_ppgen3_177 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), .b0(b0), .b1(b1), 
        .b2({net210503, net210504, net210505}), .p0m1_l(p0_l[59]), .p1m1_l(
        p1_l[59]), .p2m1_l(net210506) );
  mul_ppgen3_176 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), .b0(b0), .b1(b1), 
        .b2({net210499, net210500, net210501}), .p0m1_l(p0_l[58]), .p1m1_l(
        p1_l[58]), .p2m1_l(net210502) );
  mul_ppgen3_175 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), .b0(b0), .b1(b1), 
        .b2({net210495, net210496, net210497}), .p0m1_l(p0_l[57]), .p1m1_l(
        p1_l[57]), .p2m1_l(net210498) );
  mul_ppgen3_174 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), .b0(b0), .b1(b1), 
        .b2({net210491, net210492, net210493}), .p0m1_l(p0_l[56]), .p1m1_l(
        p1_l[56]), .p2m1_l(net210494) );
  mul_ppgen3_173 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), .b0(b0), .b1(b1), 
        .b2({net210487, net210488, net210489}), .p0m1_l(p0_l[55]), .p1m1_l(
        p1_l[55]), .p2m1_l(net210490) );
  mul_ppgen3_172 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), .b0(b0), .b1(b1), 
        .b2({net210483, net210484, net210485}), .p0m1_l(p0_l[54]), .p1m1_l(
        p1_l[54]), .p2m1_l(net210486) );
  mul_ppgen3_171 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), .b0(b0), .b1(b1), 
        .b2({net210479, net210480, net210481}), .p0m1_l(p0_l[53]), .p1m1_l(
        p1_l[53]), .p2m1_l(net210482) );
  mul_ppgen3_170 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), .b0(b0), .b1(b1), 
        .b2({net210475, net210476, net210477}), .p0m1_l(p0_l[52]), .p1m1_l(
        p1_l[52]), .p2m1_l(net210478) );
  mul_ppgen3_169 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), .b0(b0), .b1(b1), 
        .b2({net210471, net210472, net210473}), .p0m1_l(p0_l[51]), .p1m1_l(
        p1_l[51]), .p2m1_l(net210474) );
  mul_ppgen3_168 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), .b0(b0), .b1(b1), 
        .b2({net210467, net210468, net210469}), .p0m1_l(p0_l[50]), .p1m1_l(
        p1_l[50]), .p2m1_l(net210470) );
  mul_ppgen3_167 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), .b0(b0), .b1(b1), 
        .b2({net210463, net210464, net210465}), .p0m1_l(p0_l[49]), .p1m1_l(
        p1_l[49]), .p2m1_l(net210466) );
  mul_ppgen3_166 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), .b0(b0), .b1(b1), 
        .b2({net210459, net210460, net210461}), .p0m1_l(p0_l[48]), .p1m1_l(
        p1_l[48]), .p2m1_l(net210462) );
  mul_ppgen3_165 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), .b0(b0), .b1(b1), 
        .b2({net210455, net210456, net210457}), .p0m1_l(p0_l[47]), .p1m1_l(
        p1_l[47]), .p2m1_l(net210458) );
  mul_ppgen3_164 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), .b0(b0), .b1(b1), 
        .b2({net210451, net210452, net210453}), .p0m1_l(p0_l[46]), .p1m1_l(
        p1_l[46]), .p2m1_l(net210454) );
  mul_ppgen3_163 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), .b0(b0), .b1(b1), 
        .b2({net210447, net210448, net210449}), .p0m1_l(p0_l[45]), .p1m1_l(
        p1_l[45]), .p2m1_l(net210450) );
  mul_ppgen3_162 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), .b0(b0), .b1(b1), 
        .b2({net210443, net210444, net210445}), .p0m1_l(p0_l[44]), .p1m1_l(
        p1_l[44]), .p2m1_l(net210446) );
  mul_ppgen3_161 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), .b0(b0), .b1(b1), 
        .b2({net210439, net210440, net210441}), .p0m1_l(p0_l[43]), .p1m1_l(
        p1_l[43]), .p2m1_l(net210442) );
  mul_ppgen3_160 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), .b0(b0), .b1(b1), 
        .b2({net210435, net210436, net210437}), .p0m1_l(p0_l[42]), .p1m1_l(
        p1_l[42]), .p2m1_l(net210438) );
  mul_ppgen3_159 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), .b0(b0), .b1(b1), 
        .b2({net210431, net210432, net210433}), .p0m1_l(p0_l[41]), .p1m1_l(
        p1_l[41]), .p2m1_l(net210434) );
  mul_ppgen3_158 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), .b0(b0), .b1(b1), 
        .b2({net210427, net210428, net210429}), .p0m1_l(p0_l[40]), .p1m1_l(
        p1_l[40]), .p2m1_l(net210430) );
  mul_ppgen3_157 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), .b0(b0), .b1(b1), 
        .b2({net210423, net210424, net210425}), .p0m1_l(p0_l[39]), .p1m1_l(
        p1_l[39]), .p2m1_l(net210426) );
  mul_ppgen3_156 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), .b0(b0), .b1(b1), 
        .b2({net210419, net210420, net210421}), .p0m1_l(p0_l[38]), .p1m1_l(
        p1_l[38]), .p2m1_l(net210422) );
  mul_ppgen3_155 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), .b0(b0), .b1(b1), 
        .b2({net210415, net210416, net210417}), .p0m1_l(p0_l[37]), .p1m1_l(
        p1_l[37]), .p2m1_l(net210418) );
  mul_ppgen3_154 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), .b0(b0), .b1(b1), 
        .b2({net210411, net210412, net210413}), .p0m1_l(p0_l[36]), .p1m1_l(
        p1_l[36]), .p2m1_l(net210414) );
  mul_ppgen3_153 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), .b0(b0), .b1(b1), 
        .b2({net210407, net210408, net210409}), .p0m1_l(p0_l[35]), .p1m1_l(
        p1_l[35]), .p2m1_l(net210410) );
  mul_ppgen3_152 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), .b0(b0), .b1(b1), 
        .b2({net210403, net210404, net210405}), .p0m1_l(p0_l[34]), .p1m1_l(
        p1_l[34]), .p2m1_l(net210406) );
  mul_ppgen3_151 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), .b0(b0), .b1(b1), 
        .b2({net210399, net210400, net210401}), .p0m1_l(p0_l[33]), .p1m1_l(
        p1_l[33]), .p2m1_l(net210402) );
  mul_ppgen3_150 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), .b0(b0), .b1(b1), 
        .b2({net210395, net210396, net210397}), .p0m1_l(p0_l[32]), .p1m1_l(
        p1_l[32]), .p2m1_l(net210398) );
  mul_ppgen3_149 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), .b0(b0), .b1(b1), 
        .b2({net210391, net210392, net210393}), .p0m1_l(p0_l[31]), .p1m1_l(
        p1_l[31]), .p2m1_l(net210394) );
  mul_ppgen3_148 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), .b0(b0), .b1(b1), 
        .b2({net210387, net210388, net210389}), .p0m1_l(p0_l[30]), .p1m1_l(
        p1_l[30]), .p2m1_l(net210390) );
  mul_ppgen3_147 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), .b0(b0), .b1(b1), 
        .b2({net210383, net210384, net210385}), .p0m1_l(p0_l[29]), .p1m1_l(
        p1_l[29]), .p2m1_l(net210386) );
  mul_ppgen3_146 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), .b0(b0), .b1(b1), 
        .b2({net210379, net210380, net210381}), .p0m1_l(p0_l[28]), .p1m1_l(
        p1_l[28]), .p2m1_l(net210382) );
  mul_ppgen3_145 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), .b0(b0), .b1(b1), 
        .b2({net210375, net210376, net210377}), .p0m1_l(p0_l[27]), .p1m1_l(
        p1_l[27]), .p2m1_l(net210378) );
  mul_ppgen3_144 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), .b0(b0), .b1(b1), 
        .b2({net210371, net210372, net210373}), .p0m1_l(p0_l[26]), .p1m1_l(
        p1_l[26]), .p2m1_l(net210374) );
  mul_ppgen3_143 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), .b0(b0), .b1(b1), 
        .b2({net210367, net210368, net210369}), .p0m1_l(p0_l[25]), .p1m1_l(
        p1_l[25]), .p2m1_l(net210370) );
  mul_ppgen3_142 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), .b0(b0), .b1(b1), 
        .b2({net210363, net210364, net210365}), .p0m1_l(p0_l[24]), .p1m1_l(
        p1_l[24]), .p2m1_l(net210366) );
  mul_ppgen3_141 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), .b0(b0), .b1(b1), 
        .b2({net210359, net210360, net210361}), .p0m1_l(p0_l[23]), .p1m1_l(
        p1_l[23]), .p2m1_l(net210362) );
  mul_ppgen3_140 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), .b0(b0), .b1(b1), 
        .b2({net210355, net210356, net210357}), .p0m1_l(p0_l[22]), .p1m1_l(
        p1_l[22]), .p2m1_l(net210358) );
  mul_ppgen3_139 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), .b0(b0), .b1(b1), 
        .b2({net210351, net210352, net210353}), .p0m1_l(p0_l[21]), .p1m1_l(
        p1_l[21]), .p2m1_l(net210354) );
  mul_ppgen3_138 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), .b0(b0), .b1(b1), 
        .b2({net210347, net210348, net210349}), .p0m1_l(p0_l[20]), .p1m1_l(
        p1_l[20]), .p2m1_l(net210350) );
  mul_ppgen3_137 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), .b0(b0), .b1(b1), 
        .b2({net210343, net210344, net210345}), .p0m1_l(p0_l[19]), .p1m1_l(
        p1_l[19]), .p2m1_l(net210346) );
  mul_ppgen3_136 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), .b0(b0), .b1(b1), 
        .b2({net210339, net210340, net210341}), .p0m1_l(p0_l[18]), .p1m1_l(
        p1_l[18]), .p2m1_l(net210342) );
  mul_ppgen3_135 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), .b0(b0), .b1(b1), 
        .b2({net210335, net210336, net210337}), .p0m1_l(p0_l[17]), .p1m1_l(
        p1_l[17]), .p2m1_l(net210338) );
  mul_ppgen3_134 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), .b0(b0), .b1(b1), 
        .b2({net210331, net210332, net210333}), .p0m1_l(p0_l[16]), .p1m1_l(
        p1_l[16]), .p2m1_l(net210334) );
  mul_ppgen3_133 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), .b0(b0), .b1(b1), 
        .b2({net210327, net210328, net210329}), .p0m1_l(p0_l[15]), .p1m1_l(
        p1_l[15]), .p2m1_l(net210330) );
  mul_ppgen3_132 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), .b0(b0), .b1(b1), 
        .b2({net210323, net210324, net210325}), .p0m1_l(p0_l[14]), .p1m1_l(
        p1_l[14]), .p2m1_l(net210326) );
  mul_ppgen3_131 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), .b0(b0), .b1(b1), 
        .b2({net210319, net210320, net210321}), .p0m1_l(p0_l[13]), .p1m1_l(
        p1_l[13]), .p2m1_l(net210322) );
  mul_ppgen3_130 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), .b0(b0), .b1(b1), 
        .b2({net210315, net210316, net210317}), .p0m1_l(p0_l[12]), .p1m1_l(
        p1_l[12]), .p2m1_l(net210318) );
  mul_ppgen3_129 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), .b0(b0), .b1(b1), 
        .b2({net210311, net210312, net210313}), .p0m1_l(p0_l[11]), .p1m1_l(
        p1_l[11]), .p2m1_l(net210314) );
  mul_ppgen3_128 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), .b0(b0), .b1(b1), 
        .b2({net210307, net210308, net210309}), .p0m1_l(p0_l[10]), .p1m1_l(
        p1_l[10]), .p2m1_l(net210310) );
  mul_ppgen3_127 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), .b0(b0), .b1(b1), 
        .b2({net210303, net210304, net210305}), .p0m1_l(p0_l[9]), .p1m1_l(
        p1_l[9]), .p2m1_l(net210306) );
  mul_ppgen3_126 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), .sum(
        sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), .b1(b1), .b2({
        net210299, net210300, net210301}), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), 
        .p2m1_l(net210302) );
  mul_ppgen3_125 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), .sum(
        sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), .b1(b1), .b2({
        net210295, net210296, net210297}), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), 
        .p2m1_l(net210298) );
  mul_ppgen3_124 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), .sum(
        sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), .b1(b1), .b2({
        net210291, net210292, net210293}), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), 
        .p2m1_l(net210294) );
  mul_ppgen3_123 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), .sum(
        sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), .b1(b1), .b2({
        net210287, net210288, net210289}), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), 
        .p2m1_l(net210290) );
  mul_ppgen3_122 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), .sum(
        sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), .b1(b1), .b2({
        net210283, net210284, net210285}), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), 
        .p2m1_l(net210286) );
  mul_ppgen3_121 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), .sum(
        sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), .b1(b1), .b2({
        net210280, net210281, net210282}), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), 
        .p2m1_l(1'b1) );
  mul_ppgen3lsb4_3 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), 
        .sum(sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_ha_48 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_49 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_50 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_51 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_52 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   b;
  assign cout = b;

  INVX1_RVT U1 ( .A(b), .Y(sum) );
endmodule


module mul_ha_53 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_54 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_56 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   a;
  assign sum = a;

endmodule


module mul_ha_57 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_58 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_59 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_60 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  INVX0_RVT U1 ( .A(n1), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_ha_61 ( cout, sum, a, b );
  input a, b;
  output cout, sum;
  wire   n1;

  NAND2X0_RVT U1 ( .A1(b), .A2(a), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(b), .A2(a), .A3(n1), .Y(sum) );
endmodule


module mul_negen_13 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_negen_14 ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   n2;

  INVX0_RVT U1 ( .A(b[0]), .Y(n2) );
  AND3X1_RVT U2 ( .A1(b[2]), .A2(b[1]), .A3(n2), .Y(n0) );
  AND3X1_RVT U3 ( .A1(b[1]), .A2(b[2]), .A3(b[0]), .Y(n1) );
endmodule


module mul_csa32_661 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_662 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_663 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_664 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_665 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_666 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_667 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_668 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_669 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_670 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_671 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_672 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_673 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_674 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_675 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_676 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_677 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_678 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_679 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_680 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_681 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_682 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_683 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_684 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_685 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_686 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_687 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_688 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_689 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_690 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_691 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_692 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_693 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_694 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_695 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_696 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_697 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_698 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_699 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_700 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_701 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_702 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_703 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_704 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_705 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_706 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_707 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_708 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_709 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_710 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_711 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_712 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_713 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_714 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_715 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_716 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_717 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_718 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_719 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_720 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_721 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_722 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_723 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_724 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_725 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_726 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_727 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_728 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_729 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_730 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_731 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_732 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_733 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   n1;

  OR2X1_RVT U1 ( .A1(b), .A2(a), .Y(cout) );
  NAND2X0_RVT U2 ( .A1(b), .A2(a), .Y(n1) );
  NAND2X0_RVT U3 ( .A1(n1), .A2(cout), .Y(sum) );
endmodule


module mul_csa32_734 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_735 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_736 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_737 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_738 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_739 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_740 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_741 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_742 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_743 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_744 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_745 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_746 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_747 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_748 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_749 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_750 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_751 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_752 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_753 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_754 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_755 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_756 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_757 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_758 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_759 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_760 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_761 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_762 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_763 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_764 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_765 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_766 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_767 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_768 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_769 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_770 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_771 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_772 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_773 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_774 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_775 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_776 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_777 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_778 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_779 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_780 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_781 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_782 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_783 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_784 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_785 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_786 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_787 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_788 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_789 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_790 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_791 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_792 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_793 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa32_794 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;


  FADDX1_RVT U1 ( .A(c), .B(a), .CI(b), .CO(cout), .S(sum) );
endmodule


module mul_csa42_50 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  INVX0_RVT U1 ( .A(n1), .Y(carry) );
  NAND2X0_RVT U2 ( .A1(n2), .A2(b), .Y(n1) );
  OA21X1_RVT U3 ( .A1(n2), .A2(b), .A3(n1), .Y(sum) );
  FADDX1_RVT U4 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n2) );
endmodule


module mul_csa42_51 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_52 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_53 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_54 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_55 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_56 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_57 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_58 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_59 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_60 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_61 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_62 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_63 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_64 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_65 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_66 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_67 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_68 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_69 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_70 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_71 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_72 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_73 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_74 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_75 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_76 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_77 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_78 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_79 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_80 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_81 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_82 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_83 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_84 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_85 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_86 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_87 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_88 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_89 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_90 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_91 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_92 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_93 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_94 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_95 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_96 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_97 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_98 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_99 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_100 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_101 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_102 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_103 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_104 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_105 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_106 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_107 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_108 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_109 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_csa42_110 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;


  FADDX1_RVT U1 ( .A(c), .B(b), .CI(cin), .CO(carry), .S(sum) );
endmodule


module mul_csa42_111 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_112 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_113 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_114 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1, n2;

  NAND2X0_RVT U1 ( .A1(c), .A2(d), .Y(n1) );
  INVX1_RVT U2 ( .A(n1), .Y(cout) );
  OA21X1_RVT U3 ( .A1(c), .A2(d), .A3(n1), .Y(n2) );
  FADDX1_RVT U4 ( .A(b), .B(cin), .CI(n2), .CO(carry), .S(sum) );
endmodule


module mul_csa42_115 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   n1;

  FADDX1_RVT U1 ( .A(b), .B(cin), .CI(n1), .CO(carry), .S(sum) );
  FADDX1_RVT U2 ( .A(c), .B(d), .CI(a), .CO(cout), .S(n1) );
endmodule


module mul_array1_1 ( cout, sum, a, b0, b1, b2, b3, b4, b5, b6, b7, b8, bot, 
        head );
  output [81:4] cout;
  output [81:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input [2:0] b3;
  input [2:0] b4;
  input [2:0] b5;
  input [2:0] b6;
  input [2:0] b7;
  input [2:0] b8;
  input bot, head;
  wire   net210528, net210529, net210530, net210531, net210532;
  wire   [1:0] b5n;
  wire   [1:0] b2n;
  wire   [76:10] s_2;
  wire   [75:11] co;
  wire   [70:2] c_1;
  wire   [76:10] c_2;
  wire   [69:0] s1;
  wire   [70:4] s_1;
  wire   [68:1] c1;
  wire   [68:1] c2;
  wire   [69:0] s2;
  wire   [68:1] c0;
  wire   [69:2] s0;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  mul_negen_14 p1n ( .n0(b5n[0]), .n1(b5n[1]), .b(b5) );
  mul_negen_13 p0n ( .n0(b2n[0]), .n1(b2n[1]), .b(b2) );
  mul_csa42_115 sc3_71_ ( .sum(sum[71]), .carry(cout[71]), .cout(co[71]), .a(
        c_1[70]), .b(c_2[70]), .c(s_2[71]), .d(s1[65]), .cin(co[70]) );
  mul_csa42_114 sc3_75_ ( .sum(sum[75]), .carry(cout[75]), .cout(co[75]), .a(
        1'b0), .b(c_2[74]), .c(s_2[75]), .d(s1[69]), .cin(co[74]) );
  mul_csa42_113 sc3_74_ ( .sum(sum[74]), .carry(cout[74]), .cout(co[74]), .a(
        1'b0), .b(c_2[73]), .c(s_2[74]), .d(s1[68]), .cin(co[73]) );
  mul_csa42_112 sc3_73_ ( .sum(sum[73]), .carry(cout[73]), .cout(co[73]), .a(
        1'b0), .b(c_2[72]), .c(s_2[73]), .d(s1[67]), .cin(co[72]) );
  mul_csa42_111 sc3_72_ ( .sum(sum[72]), .carry(cout[72]), .cout(co[72]), .a(
        1'b0), .b(c_2[71]), .c(s_2[72]), .d(s1[66]), .cin(co[71]) );
  mul_csa42_110 sc3_76_ ( .sum(sum[76]), .carry(cout[76]), .a(1'b0), .b(
        c_2[75]), .c(s_2[76]), .d(1'b0), .cin(co[75]) );
  mul_csa42_109 sc3_70_ ( .sum(sum[70]), .carry(cout[70]), .cout(co[70]), .a(
        c_1[69]), .b(c_2[69]), .c(s_2[70]), .d(s_1[70]), .cin(co[69]) );
  mul_csa42_108 sc3_69_ ( .sum(sum[69]), .carry(cout[69]), .cout(co[69]), .a(
        c_1[68]), .b(c_2[68]), .c(s_2[69]), .d(s_1[69]), .cin(co[68]) );
  mul_csa42_107 sc3_68_ ( .sum(sum[68]), .carry(cout[68]), .cout(co[68]), .a(
        c_1[67]), .b(c_2[67]), .c(s_2[68]), .d(s_1[68]), .cin(co[67]) );
  mul_csa42_106 sc3_67_ ( .sum(sum[67]), .carry(cout[67]), .cout(co[67]), .a(
        c_1[66]), .b(c_2[66]), .c(s_2[67]), .d(s_1[67]), .cin(co[66]) );
  mul_csa42_105 sc3_66_ ( .sum(sum[66]), .carry(cout[66]), .cout(co[66]), .a(
        c_1[65]), .b(c_2[65]), .c(s_2[66]), .d(s_1[66]), .cin(co[65]) );
  mul_csa42_104 sc3_65_ ( .sum(sum[65]), .carry(cout[65]), .cout(co[65]), .a(
        c_1[64]), .b(c_2[64]), .c(s_2[65]), .d(s_1[65]), .cin(co[64]) );
  mul_csa42_103 sc3_64_ ( .sum(sum[64]), .carry(cout[64]), .cout(co[64]), .a(
        c_1[63]), .b(c_2[63]), .c(s_2[64]), .d(s_1[64]), .cin(co[63]) );
  mul_csa42_102 sc3_63_ ( .sum(sum[63]), .carry(cout[63]), .cout(co[63]), .a(
        c_1[62]), .b(c_2[62]), .c(s_2[63]), .d(s_1[63]), .cin(co[62]) );
  mul_csa42_101 sc3_62_ ( .sum(sum[62]), .carry(cout[62]), .cout(co[62]), .a(
        c_1[61]), .b(c_2[61]), .c(s_2[62]), .d(s_1[62]), .cin(co[61]) );
  mul_csa42_100 sc3_61_ ( .sum(sum[61]), .carry(cout[61]), .cout(co[61]), .a(
        c_1[60]), .b(c_2[60]), .c(s_2[61]), .d(s_1[61]), .cin(co[60]) );
  mul_csa42_99 sc3_60_ ( .sum(sum[60]), .carry(cout[60]), .cout(co[60]), .a(
        c_1[59]), .b(c_2[59]), .c(s_2[60]), .d(s_1[60]), .cin(co[59]) );
  mul_csa42_98 sc3_59_ ( .sum(sum[59]), .carry(cout[59]), .cout(co[59]), .a(
        c_1[58]), .b(c_2[58]), .c(s_2[59]), .d(s_1[59]), .cin(co[58]) );
  mul_csa42_97 sc3_58_ ( .sum(sum[58]), .carry(cout[58]), .cout(co[58]), .a(
        c_1[57]), .b(c_2[57]), .c(s_2[58]), .d(s_1[58]), .cin(co[57]) );
  mul_csa42_96 sc3_57_ ( .sum(sum[57]), .carry(cout[57]), .cout(co[57]), .a(
        c_1[56]), .b(c_2[56]), .c(s_2[57]), .d(s_1[57]), .cin(co[56]) );
  mul_csa42_95 sc3_56_ ( .sum(sum[56]), .carry(cout[56]), .cout(co[56]), .a(
        c_1[55]), .b(c_2[55]), .c(s_2[56]), .d(s_1[56]), .cin(co[55]) );
  mul_csa42_94 sc3_55_ ( .sum(sum[55]), .carry(cout[55]), .cout(co[55]), .a(
        c_1[54]), .b(c_2[54]), .c(s_2[55]), .d(s_1[55]), .cin(co[54]) );
  mul_csa42_93 sc3_54_ ( .sum(sum[54]), .carry(cout[54]), .cout(co[54]), .a(
        c_1[53]), .b(c_2[53]), .c(s_2[54]), .d(s_1[54]), .cin(co[53]) );
  mul_csa42_92 sc3_53_ ( .sum(sum[53]), .carry(cout[53]), .cout(co[53]), .a(
        c_1[52]), .b(c_2[52]), .c(s_2[53]), .d(s_1[53]), .cin(co[52]) );
  mul_csa42_91 sc3_52_ ( .sum(sum[52]), .carry(cout[52]), .cout(co[52]), .a(
        c_1[51]), .b(c_2[51]), .c(s_2[52]), .d(s_1[52]), .cin(co[51]) );
  mul_csa42_90 sc3_51_ ( .sum(sum[51]), .carry(cout[51]), .cout(co[51]), .a(
        c_1[50]), .b(c_2[50]), .c(s_2[51]), .d(s_1[51]), .cin(co[50]) );
  mul_csa42_89 sc3_50_ ( .sum(sum[50]), .carry(cout[50]), .cout(co[50]), .a(
        c_1[49]), .b(c_2[49]), .c(s_2[50]), .d(s_1[50]), .cin(co[49]) );
  mul_csa42_88 sc3_49_ ( .sum(sum[49]), .carry(cout[49]), .cout(co[49]), .a(
        c_1[48]), .b(c_2[48]), .c(s_2[49]), .d(s_1[49]), .cin(co[48]) );
  mul_csa42_87 sc3_48_ ( .sum(sum[48]), .carry(cout[48]), .cout(co[48]), .a(
        c_1[47]), .b(c_2[47]), .c(s_2[48]), .d(s_1[48]), .cin(co[47]) );
  mul_csa42_86 sc3_47_ ( .sum(sum[47]), .carry(cout[47]), .cout(co[47]), .a(
        c_1[46]), .b(c_2[46]), .c(s_2[47]), .d(s_1[47]), .cin(co[46]) );
  mul_csa42_85 sc3_46_ ( .sum(sum[46]), .carry(cout[46]), .cout(co[46]), .a(
        c_1[45]), .b(c_2[45]), .c(s_2[46]), .d(s_1[46]), .cin(co[45]) );
  mul_csa42_84 sc3_45_ ( .sum(sum[45]), .carry(cout[45]), .cout(co[45]), .a(
        c_1[44]), .b(c_2[44]), .c(s_2[45]), .d(s_1[45]), .cin(co[44]) );
  mul_csa42_83 sc3_44_ ( .sum(sum[44]), .carry(cout[44]), .cout(co[44]), .a(
        c_1[43]), .b(c_2[43]), .c(s_2[44]), .d(s_1[44]), .cin(co[43]) );
  mul_csa42_82 sc3_43_ ( .sum(sum[43]), .carry(cout[43]), .cout(co[43]), .a(
        c_1[42]), .b(c_2[42]), .c(s_2[43]), .d(s_1[43]), .cin(co[42]) );
  mul_csa42_81 sc3_42_ ( .sum(sum[42]), .carry(cout[42]), .cout(co[42]), .a(
        c_1[41]), .b(c_2[41]), .c(s_2[42]), .d(s_1[42]), .cin(co[41]) );
  mul_csa42_80 sc3_41_ ( .sum(sum[41]), .carry(cout[41]), .cout(co[41]), .a(
        c_1[40]), .b(c_2[40]), .c(s_2[41]), .d(s_1[41]), .cin(co[40]) );
  mul_csa42_79 sc3_40_ ( .sum(sum[40]), .carry(cout[40]), .cout(co[40]), .a(
        c_1[39]), .b(c_2[39]), .c(s_2[40]), .d(s_1[40]), .cin(co[39]) );
  mul_csa42_78 sc3_39_ ( .sum(sum[39]), .carry(cout[39]), .cout(co[39]), .a(
        c_1[38]), .b(c_2[38]), .c(s_2[39]), .d(s_1[39]), .cin(co[38]) );
  mul_csa42_77 sc3_38_ ( .sum(sum[38]), .carry(cout[38]), .cout(co[38]), .a(
        c_1[37]), .b(c_2[37]), .c(s_2[38]), .d(s_1[38]), .cin(co[37]) );
  mul_csa42_76 sc3_37_ ( .sum(sum[37]), .carry(cout[37]), .cout(co[37]), .a(
        c_1[36]), .b(c_2[36]), .c(s_2[37]), .d(s_1[37]), .cin(co[36]) );
  mul_csa42_75 sc3_36_ ( .sum(sum[36]), .carry(cout[36]), .cout(co[36]), .a(
        c_1[35]), .b(c_2[35]), .c(s_2[36]), .d(s_1[36]), .cin(co[35]) );
  mul_csa42_74 sc3_35_ ( .sum(sum[35]), .carry(cout[35]), .cout(co[35]), .a(
        c_1[34]), .b(c_2[34]), .c(s_2[35]), .d(s_1[35]), .cin(co[34]) );
  mul_csa42_73 sc3_34_ ( .sum(sum[34]), .carry(cout[34]), .cout(co[34]), .a(
        c_1[33]), .b(c_2[33]), .c(s_2[34]), .d(s_1[34]), .cin(co[33]) );
  mul_csa42_72 sc3_33_ ( .sum(sum[33]), .carry(cout[33]), .cout(co[33]), .a(
        c_1[32]), .b(c_2[32]), .c(s_2[33]), .d(s_1[33]), .cin(co[32]) );
  mul_csa42_71 sc3_32_ ( .sum(sum[32]), .carry(cout[32]), .cout(co[32]), .a(
        c_1[31]), .b(c_2[31]), .c(s_2[32]), .d(s_1[32]), .cin(co[31]) );
  mul_csa42_70 sc3_31_ ( .sum(sum[31]), .carry(cout[31]), .cout(co[31]), .a(
        c_1[30]), .b(c_2[30]), .c(s_2[31]), .d(s_1[31]), .cin(co[30]) );
  mul_csa42_69 sc3_30_ ( .sum(sum[30]), .carry(cout[30]), .cout(co[30]), .a(
        c_1[29]), .b(c_2[29]), .c(s_2[30]), .d(s_1[30]), .cin(co[29]) );
  mul_csa42_68 sc3_29_ ( .sum(sum[29]), .carry(cout[29]), .cout(co[29]), .a(
        c_1[28]), .b(c_2[28]), .c(s_2[29]), .d(s_1[29]), .cin(co[28]) );
  mul_csa42_67 sc3_28_ ( .sum(sum[28]), .carry(cout[28]), .cout(co[28]), .a(
        c_1[27]), .b(c_2[27]), .c(s_2[28]), .d(s_1[28]), .cin(co[27]) );
  mul_csa42_66 sc3_27_ ( .sum(sum[27]), .carry(cout[27]), .cout(co[27]), .a(
        c_1[26]), .b(c_2[26]), .c(s_2[27]), .d(s_1[27]), .cin(co[26]) );
  mul_csa42_65 sc3_26_ ( .sum(sum[26]), .carry(cout[26]), .cout(co[26]), .a(
        c_1[25]), .b(c_2[25]), .c(s_2[26]), .d(s_1[26]), .cin(co[25]) );
  mul_csa42_64 sc3_25_ ( .sum(sum[25]), .carry(cout[25]), .cout(co[25]), .a(
        c_1[24]), .b(c_2[24]), .c(s_2[25]), .d(s_1[25]), .cin(co[24]) );
  mul_csa42_63 sc3_24_ ( .sum(sum[24]), .carry(cout[24]), .cout(co[24]), .a(
        c_1[23]), .b(c_2[23]), .c(s_2[24]), .d(s_1[24]), .cin(co[23]) );
  mul_csa42_62 sc3_23_ ( .sum(sum[23]), .carry(cout[23]), .cout(co[23]), .a(
        c_1[22]), .b(c_2[22]), .c(s_2[23]), .d(s_1[23]), .cin(co[22]) );
  mul_csa42_61 sc3_22_ ( .sum(sum[22]), .carry(cout[22]), .cout(co[22]), .a(
        c_1[21]), .b(c_2[21]), .c(s_2[22]), .d(s_1[22]), .cin(co[21]) );
  mul_csa42_60 sc3_21_ ( .sum(sum[21]), .carry(cout[21]), .cout(co[21]), .a(
        c_1[20]), .b(c_2[20]), .c(s_2[21]), .d(s_1[21]), .cin(co[20]) );
  mul_csa42_59 sc3_20_ ( .sum(sum[20]), .carry(cout[20]), .cout(co[20]), .a(
        c_1[19]), .b(c_2[19]), .c(s_2[20]), .d(s_1[20]), .cin(co[19]) );
  mul_csa42_58 sc3_19_ ( .sum(sum[19]), .carry(cout[19]), .cout(co[19]), .a(
        c_1[18]), .b(c_2[18]), .c(s_2[19]), .d(s_1[19]), .cin(co[18]) );
  mul_csa42_57 sc3_18_ ( .sum(sum[18]), .carry(cout[18]), .cout(co[18]), .a(
        c_1[17]), .b(c_2[17]), .c(s_2[18]), .d(s_1[18]), .cin(co[17]) );
  mul_csa42_56 sc3_17_ ( .sum(sum[17]), .carry(cout[17]), .cout(co[17]), .a(
        c_1[16]), .b(c_2[16]), .c(s_2[17]), .d(s_1[17]), .cin(co[16]) );
  mul_csa42_55 sc3_16_ ( .sum(sum[16]), .carry(cout[16]), .cout(co[16]), .a(
        c_1[15]), .b(c_2[15]), .c(s_2[16]), .d(s_1[16]), .cin(co[15]) );
  mul_csa42_54 sc3_15_ ( .sum(sum[15]), .carry(cout[15]), .cout(co[15]), .a(
        c_1[14]), .b(c_2[14]), .c(s_2[15]), .d(s_1[15]), .cin(co[14]) );
  mul_csa42_53 sc3_14_ ( .sum(sum[14]), .carry(cout[14]), .cout(co[14]), .a(
        c_1[13]), .b(c_2[13]), .c(s_2[14]), .d(s_1[14]), .cin(co[13]) );
  mul_csa42_52 sc3_13_ ( .sum(sum[13]), .carry(cout[13]), .cout(co[13]), .a(
        c_1[12]), .b(c_2[12]), .c(s_2[13]), .d(s_1[13]), .cin(co[12]) );
  mul_csa42_51 sc3_12_ ( .sum(sum[12]), .carry(cout[12]), .cout(co[12]), .a(
        c_1[11]), .b(c_2[11]), .c(s_2[12]), .d(s_1[12]), .cin(co[11]) );
  mul_csa42_50 sc3_11_ ( .sum(sum[11]), .carry(cout[11]), .cout(co[11]), .a(
        c_1[10]), .b(c_2[10]), .c(s_2[11]), .d(s_1[11]), .cin(1'b0) );
  mul_csa32_794 sc2_2_70_ ( .sum(s_2[70]), .cout(c_2[70]), .a(s2[58]), .b(
        c2[57]), .c(c1[63]) );
  mul_csa32_793 sc2_2_69_ ( .sum(s_2[69]), .cout(c_2[69]), .a(s2[57]), .b(
        c2[56]), .c(c1[62]) );
  mul_csa32_792 sc2_2_68_ ( .sum(s_2[68]), .cout(c_2[68]), .a(s2[56]), .b(
        c2[55]), .c(c1[61]) );
  mul_csa32_791 sc2_2_67_ ( .sum(s_2[67]), .cout(c_2[67]), .a(s2[55]), .b(
        c2[54]), .c(c1[60]) );
  mul_csa32_790 sc2_2_66_ ( .sum(s_2[66]), .cout(c_2[66]), .a(s2[54]), .b(
        c2[53]), .c(c1[59]) );
  mul_csa32_789 sc2_2_65_ ( .sum(s_2[65]), .cout(c_2[65]), .a(s2[53]), .b(
        c2[52]), .c(c1[58]) );
  mul_csa32_788 sc2_2_64_ ( .sum(s_2[64]), .cout(c_2[64]), .a(s2[52]), .b(
        c2[51]), .c(c1[57]) );
  mul_csa32_787 sc2_2_63_ ( .sum(s_2[63]), .cout(c_2[63]), .a(s2[51]), .b(
        c2[50]), .c(c1[56]) );
  mul_csa32_786 sc2_2_62_ ( .sum(s_2[62]), .cout(c_2[62]), .a(s2[50]), .b(
        c2[49]), .c(c1[55]) );
  mul_csa32_785 sc2_2_61_ ( .sum(s_2[61]), .cout(c_2[61]), .a(s2[49]), .b(
        c2[48]), .c(c1[54]) );
  mul_csa32_784 sc2_2_60_ ( .sum(s_2[60]), .cout(c_2[60]), .a(s2[48]), .b(
        c2[47]), .c(c1[53]) );
  mul_csa32_783 sc2_2_59_ ( .sum(s_2[59]), .cout(c_2[59]), .a(s2[47]), .b(
        c2[46]), .c(c1[52]) );
  mul_csa32_782 sc2_2_58_ ( .sum(s_2[58]), .cout(c_2[58]), .a(s2[46]), .b(
        c2[45]), .c(c1[51]) );
  mul_csa32_781 sc2_2_57_ ( .sum(s_2[57]), .cout(c_2[57]), .a(s2[45]), .b(
        c2[44]), .c(c1[50]) );
  mul_csa32_780 sc2_2_56_ ( .sum(s_2[56]), .cout(c_2[56]), .a(s2[44]), .b(
        c2[43]), .c(c1[49]) );
  mul_csa32_779 sc2_2_55_ ( .sum(s_2[55]), .cout(c_2[55]), .a(s2[43]), .b(
        c2[42]), .c(c1[48]) );
  mul_csa32_778 sc2_2_54_ ( .sum(s_2[54]), .cout(c_2[54]), .a(s2[42]), .b(
        c2[41]), .c(c1[47]) );
  mul_csa32_777 sc2_2_53_ ( .sum(s_2[53]), .cout(c_2[53]), .a(s2[41]), .b(
        c2[40]), .c(c1[46]) );
  mul_csa32_776 sc2_2_52_ ( .sum(s_2[52]), .cout(c_2[52]), .a(s2[40]), .b(
        c2[39]), .c(c1[45]) );
  mul_csa32_775 sc2_2_51_ ( .sum(s_2[51]), .cout(c_2[51]), .a(s2[39]), .b(
        c2[38]), .c(c1[44]) );
  mul_csa32_774 sc2_2_50_ ( .sum(s_2[50]), .cout(c_2[50]), .a(s2[38]), .b(
        c2[37]), .c(c1[43]) );
  mul_csa32_773 sc2_2_49_ ( .sum(s_2[49]), .cout(c_2[49]), .a(s2[37]), .b(
        c2[36]), .c(c1[42]) );
  mul_csa32_772 sc2_2_48_ ( .sum(s_2[48]), .cout(c_2[48]), .a(s2[36]), .b(
        c2[35]), .c(c1[41]) );
  mul_csa32_771 sc2_2_47_ ( .sum(s_2[47]), .cout(c_2[47]), .a(s2[35]), .b(
        c2[34]), .c(c1[40]) );
  mul_csa32_770 sc2_2_46_ ( .sum(s_2[46]), .cout(c_2[46]), .a(s2[34]), .b(
        c2[33]), .c(c1[39]) );
  mul_csa32_769 sc2_2_45_ ( .sum(s_2[45]), .cout(c_2[45]), .a(s2[33]), .b(
        c2[32]), .c(c1[38]) );
  mul_csa32_768 sc2_2_44_ ( .sum(s_2[44]), .cout(c_2[44]), .a(s2[32]), .b(
        c2[31]), .c(c1[37]) );
  mul_csa32_767 sc2_2_43_ ( .sum(s_2[43]), .cout(c_2[43]), .a(s2[31]), .b(
        c2[30]), .c(c1[36]) );
  mul_csa32_766 sc2_2_42_ ( .sum(s_2[42]), .cout(c_2[42]), .a(s2[30]), .b(
        c2[29]), .c(c1[35]) );
  mul_csa32_765 sc2_2_41_ ( .sum(s_2[41]), .cout(c_2[41]), .a(s2[29]), .b(
        c2[28]), .c(c1[34]) );
  mul_csa32_764 sc2_2_40_ ( .sum(s_2[40]), .cout(c_2[40]), .a(s2[28]), .b(
        c2[27]), .c(c1[33]) );
  mul_csa32_763 sc2_2_39_ ( .sum(s_2[39]), .cout(c_2[39]), .a(s2[27]), .b(
        c2[26]), .c(c1[32]) );
  mul_csa32_762 sc2_2_38_ ( .sum(s_2[38]), .cout(c_2[38]), .a(s2[26]), .b(
        c2[25]), .c(c1[31]) );
  mul_csa32_761 sc2_2_37_ ( .sum(s_2[37]), .cout(c_2[37]), .a(s2[25]), .b(
        c2[24]), .c(c1[30]) );
  mul_csa32_760 sc2_2_36_ ( .sum(s_2[36]), .cout(c_2[36]), .a(s2[24]), .b(
        c2[23]), .c(c1[29]) );
  mul_csa32_759 sc2_2_35_ ( .sum(s_2[35]), .cout(c_2[35]), .a(s2[23]), .b(
        c2[22]), .c(c1[28]) );
  mul_csa32_758 sc2_2_34_ ( .sum(s_2[34]), .cout(c_2[34]), .a(s2[22]), .b(
        c2[21]), .c(c1[27]) );
  mul_csa32_757 sc2_2_33_ ( .sum(s_2[33]), .cout(c_2[33]), .a(s2[21]), .b(
        c2[20]), .c(c1[26]) );
  mul_csa32_756 sc2_2_32_ ( .sum(s_2[32]), .cout(c_2[32]), .a(s2[20]), .b(
        c2[19]), .c(c1[25]) );
  mul_csa32_755 sc2_2_31_ ( .sum(s_2[31]), .cout(c_2[31]), .a(s2[19]), .b(
        c2[18]), .c(c1[24]) );
  mul_csa32_754 sc2_2_30_ ( .sum(s_2[30]), .cout(c_2[30]), .a(s2[18]), .b(
        c2[17]), .c(c1[23]) );
  mul_csa32_753 sc2_2_29_ ( .sum(s_2[29]), .cout(c_2[29]), .a(s2[17]), .b(
        c2[16]), .c(c1[22]) );
  mul_csa32_752 sc2_2_28_ ( .sum(s_2[28]), .cout(c_2[28]), .a(s2[16]), .b(
        c2[15]), .c(c1[21]) );
  mul_csa32_751 sc2_2_27_ ( .sum(s_2[27]), .cout(c_2[27]), .a(s2[15]), .b(
        c2[14]), .c(c1[20]) );
  mul_csa32_750 sc2_2_26_ ( .sum(s_2[26]), .cout(c_2[26]), .a(s2[14]), .b(
        c2[13]), .c(c1[19]) );
  mul_csa32_749 sc2_2_25_ ( .sum(s_2[25]), .cout(c_2[25]), .a(s2[13]), .b(
        c2[12]), .c(c1[18]) );
  mul_csa32_748 sc2_2_24_ ( .sum(s_2[24]), .cout(c_2[24]), .a(s2[12]), .b(
        c2[11]), .c(c1[17]) );
  mul_csa32_747 sc2_2_23_ ( .sum(s_2[23]), .cout(c_2[23]), .a(s2[11]), .b(
        c2[10]), .c(c1[16]) );
  mul_csa32_746 sc2_2_22_ ( .sum(s_2[22]), .cout(c_2[22]), .a(s2[10]), .b(
        c2[9]), .c(c1[15]) );
  mul_csa32_745 sc2_2_21_ ( .sum(s_2[21]), .cout(c_2[21]), .a(s2[9]), .b(c2[8]), .c(c1[14]) );
  mul_csa32_744 sc2_2_20_ ( .sum(s_2[20]), .cout(c_2[20]), .a(s2[8]), .b(c2[7]), .c(c1[13]) );
  mul_csa32_743 sc2_2_19_ ( .sum(s_2[19]), .cout(c_2[19]), .a(s2[7]), .b(c2[6]), .c(c1[12]) );
  mul_csa32_742 sc2_2_18_ ( .sum(s_2[18]), .cout(c_2[18]), .a(s2[6]), .b(c2[5]), .c(c1[11]) );
  mul_csa32_741 sc2_2_17_ ( .sum(s_2[17]), .cout(c_2[17]), .a(s2[5]), .b(c2[4]), .c(c1[10]) );
  mul_csa32_740 sc2_2_16_ ( .sum(s_2[16]), .cout(c_2[16]), .a(s2[4]), .b(c2[3]), .c(c1[9]) );
  mul_csa32_739 sc2_2_15_ ( .sum(s_2[15]), .cout(c_2[15]), .a(s2[3]), .b(c2[2]), .c(c1[8]) );
  mul_csa32_738 sc2_2_14_ ( .sum(s_2[14]), .cout(c_2[14]), .a(s2[2]), .b(c2[1]), .c(c1[7]) );
  mul_csa32_737 sc2_2_13_ ( .sum(s_2[13]), .cout(c_2[13]), .a(s2[1]), .b(s1[7]), .c(c1[6]) );
  mul_csa32_736 sc2_2_12_ ( .sum(s_2[12]), .cout(c_2[12]), .a(s2[0]), .b(s1[6]), .c(c1[5]) );
  mul_csa32_735 sc2_2_11_ ( .sum(s_2[11]), .cout(c_2[11]), .a(b5n[1]), .b(
        s1[5]), .c(c1[4]) );
  mul_csa32_734 sc2_2_10_ ( .sum(s_2[10]), .cout(c_2[10]), .a(b5n[0]), .b(
        s1[4]), .c(c1[3]) );
  mul_csa32_733 sc2_2_76_ ( .sum(s_2[76]), .cout(c_2[76]), .a(s2[64]), .b(
        c2[63]), .c(1'b1) );
  mul_csa32_732 sc2_2_77_ ( .sum(sum[77]), .cout(cout[77]), .a(s2[65]), .b(
        c2[64]), .c(c_2[76]) );
  mul_csa32_731 sc2_1_9_ ( .sum(s_1[9]), .cout(c_1[9]), .a(s0[9]), .b(c0[8]), 
        .c(s1[3]) );
  mul_csa32_730 sc2_1_8_ ( .sum(s_1[8]), .cout(c_1[8]), .a(s0[8]), .b(c0[7]), 
        .c(s1[2]) );
  mul_csa32_729 sc2_1_3_ ( .sum(sum[3]), .cout(c_1[3]), .a(s0[3]), .b(c0[2]), 
        .c(c_1[2]) );
  mul_csa32_728 sc3_10_ ( .sum(sum[10]), .cout(cout[10]), .a(c_1[9]), .b(
        s_1[10]), .c(s_2[10]) );
  mul_csa32_727 sc3_9_ ( .sum(sum[9]), .cout(cout[9]), .a(c_1[8]), .b(s_1[9]), 
        .c(c1[2]) );
  mul_csa32_726 sc3_8_ ( .sum(sum[8]), .cout(cout[8]), .a(c_1[7]), .b(s_1[8]), 
        .c(c1[1]) );
  mul_csa32_725 sc2_2_71_ ( .sum(s_2[71]), .cout(c_2[71]), .a(s2[59]), .b(
        c2[58]), .c(c1[64]) );
  mul_csa32_724 sc2_2_75_ ( .sum(s_2[75]), .cout(c_2[75]), .a(s2[63]), .b(
        c2[62]), .c(c1[68]) );
  mul_csa32_723 sc2_2_74_ ( .sum(s_2[74]), .cout(c_2[74]), .a(s2[62]), .b(
        c2[61]), .c(c1[67]) );
  mul_csa32_722 sc2_2_73_ ( .sum(s_2[73]), .cout(c_2[73]), .a(s2[61]), .b(
        c2[60]), .c(c1[66]) );
  mul_csa32_721 sc2_2_72_ ( .sum(s_2[72]), .cout(c_2[72]), .a(s2[60]), .b(
        c2[59]), .c(c1[65]) );
  mul_csa32_720 sc2_1_69_ ( .sum(s_1[69]), .cout(c_1[69]), .a(s0[69]), .b(
        c0[68]), .c(s1[63]) );
  mul_csa32_719 sc2_1_68_ ( .sum(s_1[68]), .cout(c_1[68]), .a(s0[68]), .b(
        c0[67]), .c(s1[62]) );
  mul_csa32_718 sc2_1_67_ ( .sum(s_1[67]), .cout(c_1[67]), .a(s0[67]), .b(
        c0[66]), .c(s1[61]) );
  mul_csa32_717 sc2_1_66_ ( .sum(s_1[66]), .cout(c_1[66]), .a(s0[66]), .b(
        c0[65]), .c(s1[60]) );
  mul_csa32_716 sc2_1_65_ ( .sum(s_1[65]), .cout(c_1[65]), .a(s0[65]), .b(
        c0[64]), .c(s1[59]) );
  mul_csa32_715 sc2_1_64_ ( .sum(s_1[64]), .cout(c_1[64]), .a(s0[64]), .b(
        c0[63]), .c(s1[58]) );
  mul_csa32_714 sc2_1_63_ ( .sum(s_1[63]), .cout(c_1[63]), .a(s0[63]), .b(
        c0[62]), .c(s1[57]) );
  mul_csa32_713 sc2_1_62_ ( .sum(s_1[62]), .cout(c_1[62]), .a(s0[62]), .b(
        c0[61]), .c(s1[56]) );
  mul_csa32_712 sc2_1_61_ ( .sum(s_1[61]), .cout(c_1[61]), .a(s0[61]), .b(
        c0[60]), .c(s1[55]) );
  mul_csa32_711 sc2_1_60_ ( .sum(s_1[60]), .cout(c_1[60]), .a(s0[60]), .b(
        c0[59]), .c(s1[54]) );
  mul_csa32_710 sc2_1_59_ ( .sum(s_1[59]), .cout(c_1[59]), .a(s0[59]), .b(
        c0[58]), .c(s1[53]) );
  mul_csa32_709 sc2_1_58_ ( .sum(s_1[58]), .cout(c_1[58]), .a(s0[58]), .b(
        c0[57]), .c(s1[52]) );
  mul_csa32_708 sc2_1_57_ ( .sum(s_1[57]), .cout(c_1[57]), .a(s0[57]), .b(
        c0[56]), .c(s1[51]) );
  mul_csa32_707 sc2_1_56_ ( .sum(s_1[56]), .cout(c_1[56]), .a(s0[56]), .b(
        c0[55]), .c(s1[50]) );
  mul_csa32_706 sc2_1_55_ ( .sum(s_1[55]), .cout(c_1[55]), .a(s0[55]), .b(
        c0[54]), .c(s1[49]) );
  mul_csa32_705 sc2_1_54_ ( .sum(s_1[54]), .cout(c_1[54]), .a(s0[54]), .b(
        c0[53]), .c(s1[48]) );
  mul_csa32_704 sc2_1_53_ ( .sum(s_1[53]), .cout(c_1[53]), .a(s0[53]), .b(
        c0[52]), .c(s1[47]) );
  mul_csa32_703 sc2_1_52_ ( .sum(s_1[52]), .cout(c_1[52]), .a(s0[52]), .b(
        c0[51]), .c(s1[46]) );
  mul_csa32_702 sc2_1_51_ ( .sum(s_1[51]), .cout(c_1[51]), .a(s0[51]), .b(
        c0[50]), .c(s1[45]) );
  mul_csa32_701 sc2_1_50_ ( .sum(s_1[50]), .cout(c_1[50]), .a(s0[50]), .b(
        c0[49]), .c(s1[44]) );
  mul_csa32_700 sc2_1_49_ ( .sum(s_1[49]), .cout(c_1[49]), .a(s0[49]), .b(
        c0[48]), .c(s1[43]) );
  mul_csa32_699 sc2_1_48_ ( .sum(s_1[48]), .cout(c_1[48]), .a(s0[48]), .b(
        c0[47]), .c(s1[42]) );
  mul_csa32_698 sc2_1_47_ ( .sum(s_1[47]), .cout(c_1[47]), .a(s0[47]), .b(
        c0[46]), .c(s1[41]) );
  mul_csa32_697 sc2_1_46_ ( .sum(s_1[46]), .cout(c_1[46]), .a(s0[46]), .b(
        c0[45]), .c(s1[40]) );
  mul_csa32_696 sc2_1_45_ ( .sum(s_1[45]), .cout(c_1[45]), .a(s0[45]), .b(
        c0[44]), .c(s1[39]) );
  mul_csa32_695 sc2_1_44_ ( .sum(s_1[44]), .cout(c_1[44]), .a(s0[44]), .b(
        c0[43]), .c(s1[38]) );
  mul_csa32_694 sc2_1_43_ ( .sum(s_1[43]), .cout(c_1[43]), .a(s0[43]), .b(
        c0[42]), .c(s1[37]) );
  mul_csa32_693 sc2_1_42_ ( .sum(s_1[42]), .cout(c_1[42]), .a(s0[42]), .b(
        c0[41]), .c(s1[36]) );
  mul_csa32_692 sc2_1_41_ ( .sum(s_1[41]), .cout(c_1[41]), .a(s0[41]), .b(
        c0[40]), .c(s1[35]) );
  mul_csa32_691 sc2_1_40_ ( .sum(s_1[40]), .cout(c_1[40]), .a(s0[40]), .b(
        c0[39]), .c(s1[34]) );
  mul_csa32_690 sc2_1_39_ ( .sum(s_1[39]), .cout(c_1[39]), .a(s0[39]), .b(
        c0[38]), .c(s1[33]) );
  mul_csa32_689 sc2_1_38_ ( .sum(s_1[38]), .cout(c_1[38]), .a(s0[38]), .b(
        c0[37]), .c(s1[32]) );
  mul_csa32_688 sc2_1_37_ ( .sum(s_1[37]), .cout(c_1[37]), .a(s0[37]), .b(
        c0[36]), .c(s1[31]) );
  mul_csa32_687 sc2_1_36_ ( .sum(s_1[36]), .cout(c_1[36]), .a(s0[36]), .b(
        c0[35]), .c(s1[30]) );
  mul_csa32_686 sc2_1_35_ ( .sum(s_1[35]), .cout(c_1[35]), .a(s0[35]), .b(
        c0[34]), .c(s1[29]) );
  mul_csa32_685 sc2_1_34_ ( .sum(s_1[34]), .cout(c_1[34]), .a(s0[34]), .b(
        c0[33]), .c(s1[28]) );
  mul_csa32_684 sc2_1_33_ ( .sum(s_1[33]), .cout(c_1[33]), .a(s0[33]), .b(
        c0[32]), .c(s1[27]) );
  mul_csa32_683 sc2_1_32_ ( .sum(s_1[32]), .cout(c_1[32]), .a(s0[32]), .b(
        c0[31]), .c(s1[26]) );
  mul_csa32_682 sc2_1_31_ ( .sum(s_1[31]), .cout(c_1[31]), .a(s0[31]), .b(
        c0[30]), .c(s1[25]) );
  mul_csa32_681 sc2_1_30_ ( .sum(s_1[30]), .cout(c_1[30]), .a(s0[30]), .b(
        c0[29]), .c(s1[24]) );
  mul_csa32_680 sc2_1_29_ ( .sum(s_1[29]), .cout(c_1[29]), .a(s0[29]), .b(
        c0[28]), .c(s1[23]) );
  mul_csa32_679 sc2_1_28_ ( .sum(s_1[28]), .cout(c_1[28]), .a(s0[28]), .b(
        c0[27]), .c(s1[22]) );
  mul_csa32_678 sc2_1_27_ ( .sum(s_1[27]), .cout(c_1[27]), .a(s0[27]), .b(
        c0[26]), .c(s1[21]) );
  mul_csa32_677 sc2_1_26_ ( .sum(s_1[26]), .cout(c_1[26]), .a(s0[26]), .b(
        c0[25]), .c(s1[20]) );
  mul_csa32_676 sc2_1_25_ ( .sum(s_1[25]), .cout(c_1[25]), .a(s0[25]), .b(
        c0[24]), .c(s1[19]) );
  mul_csa32_675 sc2_1_24_ ( .sum(s_1[24]), .cout(c_1[24]), .a(s0[24]), .b(
        c0[23]), .c(s1[18]) );
  mul_csa32_674 sc2_1_23_ ( .sum(s_1[23]), .cout(c_1[23]), .a(s0[23]), .b(
        c0[22]), .c(s1[17]) );
  mul_csa32_673 sc2_1_22_ ( .sum(s_1[22]), .cout(c_1[22]), .a(s0[22]), .b(
        c0[21]), .c(s1[16]) );
  mul_csa32_672 sc2_1_21_ ( .sum(s_1[21]), .cout(c_1[21]), .a(s0[21]), .b(
        c0[20]), .c(s1[15]) );
  mul_csa32_671 sc2_1_20_ ( .sum(s_1[20]), .cout(c_1[20]), .a(s0[20]), .b(
        c0[19]), .c(s1[14]) );
  mul_csa32_670 sc2_1_19_ ( .sum(s_1[19]), .cout(c_1[19]), .a(s0[19]), .b(
        c0[18]), .c(s1[13]) );
  mul_csa32_669 sc2_1_18_ ( .sum(s_1[18]), .cout(c_1[18]), .a(s0[18]), .b(
        c0[17]), .c(s1[12]) );
  mul_csa32_668 sc2_1_17_ ( .sum(s_1[17]), .cout(c_1[17]), .a(s0[17]), .b(
        c0[16]), .c(s1[11]) );
  mul_csa32_667 sc2_1_16_ ( .sum(s_1[16]), .cout(c_1[16]), .a(s0[16]), .b(
        c0[15]), .c(s1[10]) );
  mul_csa32_666 sc2_1_15_ ( .sum(s_1[15]), .cout(c_1[15]), .a(s0[15]), .b(
        c0[14]), .c(s1[9]) );
  mul_csa32_665 sc2_1_14_ ( .sum(s_1[14]), .cout(c_1[14]), .a(s0[14]), .b(
        c0[13]), .c(s1[8]) );
  mul_csa32_664 sc2_1_7_ ( .sum(s_1[7]), .cout(c_1[7]), .a(s0[7]), .b(c0[6]), 
        .c(s1[1]) );
  mul_csa32_663 sc2_1_6_ ( .sum(s_1[6]), .cout(c_1[6]), .a(s0[6]), .b(c0[5]), 
        .c(s1[0]) );
  mul_csa32_662 sc2_1_5_ ( .sum(s_1[5]), .cout(c_1[5]), .a(s0[5]), .b(c0[4]), 
        .c(b2n[1]) );
  mul_csa32_661 sc2_1_4_ ( .sum(s_1[4]), .cout(c_1[4]), .a(s0[4]), .b(c0[3]), 
        .c(b2n[0]) );
  mul_ha_61 sc2_1_10_ ( .cout(c_1[10]), .sum(s_1[10]), .a(s0[10]), .b(c0[9])
         );
  mul_ha_60 sc3_7_ ( .cout(cout[7]), .sum(sum[7]), .a(c_1[6]), .b(s_1[7]) );
  mul_ha_59 sc3_6_ ( .cout(cout[6]), .sum(sum[6]), .a(c_1[5]), .b(s_1[6]) );
  mul_ha_58 sc3_5_ ( .cout(cout[5]), .sum(sum[5]), .a(c_1[4]), .b(s_1[5]) );
  mul_ha_57 sc3_4_ ( .cout(cout[4]), .sum(sum[4]), .a(c_1[3]), .b(s_1[4]) );
  mul_ha_56 sc2_2_81_ ( .sum(sum[81]), .a(s2[69]), .b(net210532) );
  mul_ha_54 sc2_2_79_ ( .cout(cout[79]), .sum(sum[79]), .a(s2[67]), .b(c2[66])
         );
  mul_ha_53 sc2_2_78_ ( .cout(cout[78]), .sum(sum[78]), .a(s2[66]), .b(c2[65])
         );
  mul_ha_52 sc2_1_70_ ( .cout(c_1[70]), .sum(s_1[70]), .a(1'b1), .b(s1[64]) );
  mul_ha_51 sc2_1_2_ ( .cout(c_1[2]), .sum(sum[2]), .a(s0[2]), .b(c0[1]) );
  mul_ha_50 sc2_1_13_ ( .cout(c_1[13]), .sum(s_1[13]), .a(s0[13]), .b(c0[12])
         );
  mul_ha_49 sc2_1_12_ ( .cout(c_1[12]), .sum(s_1[12]), .a(s0[12]), .b(c0[11])
         );
  mul_ha_48 sc2_1_11_ ( .cout(c_1[11]), .sum(s_1[11]), .a(s0[11]), .b(c0[10])
         );
  mul_ppgenrow3_3 I2 ( .cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        c2[66:1]}), .sum({s2[69], SYNOPSYS_UNCONNECTED__2, s2[67:0]}), .a(a), 
        .b0(b6), .b1(b7), .b2({net210529, net210530, net210531}), .bot(bot), 
        .head(1'b0) );
  mul_ppgenrow3_2 I1 ( .cout(c1), .sum(s1), .a(a), .b0(b3), .b1(b4), .b2(b5), 
        .bot(1'b1), .head(1'b0) );
  mul_ppgenrow3_1 I0 ( .cout(c0), .sum({s0, sum[1:0]}), .a(a), .b0(b0), .b1(b1), .b2(b2), .bot(1'b1), .head(net210528) );
endmodule


module clken_buf_6 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module clken_buf_7 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module dffr_SIZE1_9 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dffr_SIZE1_8 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dffr_SIZE1_7 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dff_SIZE64_1 ( din, clk, se, si, \q[63]_BAR , \so[63]_BAR , \q[62]_BAR , 
        \so[62]_BAR , \q[61]_BAR , \so[61]_BAR , \q[60]_BAR , \so[60]_BAR , 
        \q[59]_BAR , \so[59]_BAR , \q[58]_BAR , \so[58]_BAR , \q[57]_BAR , 
        \so[57]_BAR , \q[56]_BAR , \so[56]_BAR , \q[55]_BAR , \so[55]_BAR , 
        \q[54]_BAR , \so[54]_BAR , \q[53]_BAR , \so[53]_BAR , \q[52]_BAR , 
        \so[52]_BAR , \q[51]_BAR , \so[51]_BAR , \q[50]_BAR , \so[50]_BAR , 
        \q[49]_BAR , \so[49]_BAR , \q[48]_BAR , \so[48]_BAR , \q[47]_BAR , 
        \so[47]_BAR , \q[46]_BAR , \so[46]_BAR , \q[45]_BAR , \so[45]_BAR , 
        \q[44]_BAR , \so[44]_BAR , \q[43]_BAR , \so[43]_BAR , \q[42]_BAR , 
        \so[42]_BAR , \q[41]_BAR , \so[41]_BAR , \q[40]_BAR , \so[40]_BAR , 
        \q[39]_BAR , \so[39]_BAR , \q[38]_BAR , \so[38]_BAR , \q[37]_BAR , 
        \so[37]_BAR , \q[36]_BAR , \so[36]_BAR , \q[35]_BAR , \so[35]_BAR , 
        \q[34]_BAR , \so[34]_BAR , \q[33]_BAR , \so[33]_BAR , \q[32]_BAR , 
        \so[32]_BAR , \q[31]_BAR , \so[31]_BAR , \q[30]_BAR , \so[30]_BAR , 
        \q[29]_BAR , \so[29]_BAR , \q[28]_BAR , \so[28]_BAR , \q[27]_BAR , 
        \so[27]_BAR , \q[26]_BAR , \so[26]_BAR , \q[25]_BAR , \so[25]_BAR , 
        \q[24]_BAR , \so[24]_BAR , \q[23]_BAR , \so[23]_BAR , \q[22]_BAR , 
        \so[22]_BAR , \q[21]_BAR , \so[21]_BAR , \q[20]_BAR , \so[20]_BAR , 
        \q[19]_BAR , \so[19]_BAR , \q[18]_BAR , \so[18]_BAR , \q[17]_BAR , 
        \so[17]_BAR , \q[16]_BAR , \so[16]_BAR , \q[15]_BAR , \so[15]_BAR , 
        \q[14]_BAR , \so[14]_BAR , \q[13]_BAR , \so[13]_BAR , \q[12]_BAR , 
        \so[12]_BAR , \q[11]_BAR , \so[11]_BAR , \q[10]_BAR , \so[10]_BAR , 
        \q[9]_BAR , \so[9]_BAR , \q[8]_BAR , \so[8]_BAR , \q[7]_BAR , 
        \so[7]_BAR , \q[6]_BAR , \so[6]_BAR , \q[5]_BAR , \so[5]_BAR , 
        \q[4]_BAR , \so[4]_BAR , \q[3]_BAR , \so[3]_BAR , \q[2]_BAR , 
        \so[2]_BAR , \q[1]_BAR , \so[1]_BAR , \q[0]_BAR , \so[0]_BAR  );
  input [63:0] din;
  input [63:0] si;
  input clk, se;
  output \q[63]_BAR , \so[63]_BAR , \q[62]_BAR , \so[62]_BAR , \q[61]_BAR ,
         \so[61]_BAR , \q[60]_BAR , \so[60]_BAR , \q[59]_BAR , \so[59]_BAR ,
         \q[58]_BAR , \so[58]_BAR , \q[57]_BAR , \so[57]_BAR , \q[56]_BAR ,
         \so[56]_BAR , \q[55]_BAR , \so[55]_BAR , \q[54]_BAR , \so[54]_BAR ,
         \q[53]_BAR , \so[53]_BAR , \q[52]_BAR , \so[52]_BAR , \q[51]_BAR ,
         \so[51]_BAR , \q[50]_BAR , \so[50]_BAR , \q[49]_BAR , \so[49]_BAR ,
         \q[48]_BAR , \so[48]_BAR , \q[47]_BAR , \so[47]_BAR , \q[46]_BAR ,
         \so[46]_BAR , \q[45]_BAR , \so[45]_BAR , \q[44]_BAR , \so[44]_BAR ,
         \q[43]_BAR , \so[43]_BAR , \q[42]_BAR , \so[42]_BAR , \q[41]_BAR ,
         \so[41]_BAR , \q[40]_BAR , \so[40]_BAR , \q[39]_BAR , \so[39]_BAR ,
         \q[38]_BAR , \so[38]_BAR , \q[37]_BAR , \so[37]_BAR , \q[36]_BAR ,
         \so[36]_BAR , \q[35]_BAR , \so[35]_BAR , \q[34]_BAR , \so[34]_BAR ,
         \q[33]_BAR , \so[33]_BAR , \q[32]_BAR , \so[32]_BAR , \q[31]_BAR ,
         \so[31]_BAR , \q[30]_BAR , \so[30]_BAR , \q[29]_BAR , \so[29]_BAR ,
         \q[28]_BAR , \so[28]_BAR , \q[27]_BAR , \so[27]_BAR , \q[26]_BAR ,
         \so[26]_BAR , \q[25]_BAR , \so[25]_BAR , \q[24]_BAR , \so[24]_BAR ,
         \q[23]_BAR , \so[23]_BAR , \q[22]_BAR , \so[22]_BAR , \q[21]_BAR ,
         \so[21]_BAR , \q[20]_BAR , \so[20]_BAR , \q[19]_BAR , \so[19]_BAR ,
         \q[18]_BAR , \so[18]_BAR , \q[17]_BAR , \so[17]_BAR , \q[16]_BAR ,
         \so[16]_BAR , \q[15]_BAR , \so[15]_BAR , \q[14]_BAR , \so[14]_BAR ,
         \q[13]_BAR , \so[13]_BAR , \q[12]_BAR , \so[12]_BAR , \q[11]_BAR ,
         \so[11]_BAR , \q[10]_BAR , \so[10]_BAR , \q[9]_BAR , \so[9]_BAR ,
         \q[8]_BAR , \so[8]_BAR , \q[7]_BAR , \so[7]_BAR , \q[6]_BAR ,
         \so[6]_BAR , \q[5]_BAR , \so[5]_BAR , \q[4]_BAR , \so[4]_BAR ,
         \q[3]_BAR , \so[3]_BAR , \q[2]_BAR , \so[2]_BAR , \q[1]_BAR ,
         \so[1]_BAR , \q[0]_BAR , \so[0]_BAR ;
  wire   n54, \so[0]_BAR , \so[1]_BAR , \so[2]_BAR , \so[3]_BAR , \so[4]_BAR ,
         \so[5]_BAR , \so[6]_BAR , \so[7]_BAR , \so[8]_BAR , \so[9]_BAR ,
         \so[10]_BAR , \so[11]_BAR , \so[12]_BAR , \so[13]_BAR , \so[14]_BAR ,
         \so[15]_BAR , \so[16]_BAR , \so[17]_BAR , \so[18]_BAR , \so[19]_BAR ,
         \so[20]_BAR , \so[21]_BAR , \so[22]_BAR , \so[23]_BAR , \so[24]_BAR ,
         \so[25]_BAR , \so[26]_BAR , \so[27]_BAR , \so[28]_BAR , \so[29]_BAR ,
         \so[30]_BAR , \so[31]_BAR , \so[32]_BAR , \so[33]_BAR , \so[34]_BAR ,
         \so[35]_BAR , \so[36]_BAR , \so[37]_BAR , \so[38]_BAR , \so[39]_BAR ,
         \so[40]_BAR , \so[41]_BAR , \so[42]_BAR , \so[43]_BAR , \so[44]_BAR ,
         \so[45]_BAR , \so[46]_BAR , \so[47]_BAR , \so[48]_BAR , \so[49]_BAR ,
         \so[50]_BAR , \so[51]_BAR , \so[52]_BAR , \q[53]_BAR ;
  assign \q[0]_BAR  = \so[0]_BAR ;
  assign \q[1]_BAR  = \so[1]_BAR ;
  assign \q[2]_BAR  = \so[2]_BAR ;
  assign \q[3]_BAR  = \so[3]_BAR ;
  assign \q[4]_BAR  = \so[4]_BAR ;
  assign \q[5]_BAR  = \so[5]_BAR ;
  assign \q[6]_BAR  = \so[6]_BAR ;
  assign \q[7]_BAR  = \so[7]_BAR ;
  assign \q[8]_BAR  = \so[8]_BAR ;
  assign \q[9]_BAR  = \so[9]_BAR ;
  assign \q[10]_BAR  = \so[10]_BAR ;
  assign \q[11]_BAR  = \so[11]_BAR ;
  assign \q[12]_BAR  = \so[12]_BAR ;
  assign \q[13]_BAR  = \so[13]_BAR ;
  assign \q[14]_BAR  = \so[14]_BAR ;
  assign \q[15]_BAR  = \so[15]_BAR ;
  assign \q[16]_BAR  = \so[16]_BAR ;
  assign \q[17]_BAR  = \so[17]_BAR ;
  assign \q[18]_BAR  = \so[18]_BAR ;
  assign \q[19]_BAR  = \so[19]_BAR ;
  assign \q[20]_BAR  = \so[20]_BAR ;
  assign \q[21]_BAR  = \so[21]_BAR ;
  assign \q[22]_BAR  = \so[22]_BAR ;
  assign \q[23]_BAR  = \so[23]_BAR ;
  assign \q[24]_BAR  = \so[24]_BAR ;
  assign \q[25]_BAR  = \so[25]_BAR ;
  assign \q[26]_BAR  = \so[26]_BAR ;
  assign \q[27]_BAR  = \so[27]_BAR ;
  assign \q[28]_BAR  = \so[28]_BAR ;
  assign \q[29]_BAR  = \so[29]_BAR ;
  assign \q[30]_BAR  = \so[30]_BAR ;
  assign \q[31]_BAR  = \so[31]_BAR ;
  assign \q[32]_BAR  = \so[32]_BAR ;
  assign \q[33]_BAR  = \so[33]_BAR ;
  assign \q[34]_BAR  = \so[34]_BAR ;
  assign \q[35]_BAR  = \so[35]_BAR ;
  assign \q[36]_BAR  = \so[36]_BAR ;
  assign \q[37]_BAR  = \so[37]_BAR ;
  assign \q[38]_BAR  = \so[38]_BAR ;
  assign \q[39]_BAR  = \so[39]_BAR ;
  assign \q[40]_BAR  = \so[40]_BAR ;
  assign \q[41]_BAR  = \so[41]_BAR ;
  assign \q[42]_BAR  = \so[42]_BAR ;
  assign \q[43]_BAR  = \so[43]_BAR ;
  assign \q[44]_BAR  = \so[44]_BAR ;
  assign \q[45]_BAR  = \so[45]_BAR ;
  assign \q[46]_BAR  = \so[46]_BAR ;
  assign \q[47]_BAR  = \so[47]_BAR ;
  assign \q[48]_BAR  = \so[48]_BAR ;
  assign \q[49]_BAR  = \so[49]_BAR ;
  assign \q[50]_BAR  = \so[50]_BAR ;
  assign \q[51]_BAR  = \so[51]_BAR ;
  assign \q[52]_BAR  = \so[52]_BAR ;
  assign \so[63]_BAR  = \q[53]_BAR ;
  assign \so[54]_BAR  = \q[53]_BAR ;
  assign \so[55]_BAR  = \q[53]_BAR ;
  assign \so[62]_BAR  = \q[53]_BAR ;
  assign \so[56]_BAR  = \q[53]_BAR ;
  assign \so[53]_BAR  = \q[53]_BAR ;
  assign \so[57]_BAR  = \q[53]_BAR ;
  assign \so[61]_BAR  = \q[53]_BAR ;
  assign \so[58]_BAR  = \q[53]_BAR ;
  assign \so[59]_BAR  = \q[53]_BAR ;
  assign \so[60]_BAR  = \q[53]_BAR ;
  assign \q[63]_BAR  = \q[53]_BAR ;
  assign \q[62]_BAR  = \q[53]_BAR ;
  assign \q[60]_BAR  = \q[53]_BAR ;
  assign \q[61]_BAR  = \q[53]_BAR ;
  assign \q[59]_BAR  = \q[53]_BAR ;
  assign \q[58]_BAR  = \q[53]_BAR ;
  assign \q[57]_BAR  = \q[53]_BAR ;
  assign \q[56]_BAR  = \q[53]_BAR ;
  assign \q[55]_BAR  = \q[53]_BAR ;
  assign \q[54]_BAR  = \q[53]_BAR ;

  DFFX1_RVT \q_reg[63]  ( .D(n54), .CLK(clk), .QN(\q[53]_BAR ) );
  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\so[0]_BAR ) );
  DFFSSRX1_RVT \q_reg[5]  ( .D(1'b0), .SETB(se), .RSTB(din[5]), .CLK(clk), 
        .QN(\so[5]_BAR ) );
  DFFSSRX1_RVT \q_reg[4]  ( .D(1'b0), .SETB(se), .RSTB(din[4]), .CLK(clk), 
        .QN(\so[4]_BAR ) );
  DFFSSRX1_RVT \q_reg[3]  ( .D(1'b0), .SETB(se), .RSTB(din[3]), .CLK(clk), 
        .QN(\so[3]_BAR ) );
  DFFSSRX1_RVT \q_reg[2]  ( .D(1'b0), .SETB(se), .RSTB(din[2]), .CLK(clk), 
        .QN(\so[2]_BAR ) );
  DFFSSRX1_RVT \q_reg[1]  ( .D(1'b0), .SETB(se), .RSTB(din[1]), .CLK(clk), 
        .QN(\so[1]_BAR ) );
  DFFSSRX1_RVT \q_reg[28]  ( .D(1'b0), .SETB(se), .RSTB(din[28]), .CLK(clk), 
        .QN(\so[28]_BAR ) );
  DFFSSRX1_RVT \q_reg[27]  ( .D(1'b0), .SETB(se), .RSTB(din[27]), .CLK(clk), 
        .QN(\so[27]_BAR ) );
  DFFSSRX1_RVT \q_reg[26]  ( .D(1'b0), .SETB(se), .RSTB(din[26]), .CLK(clk), 
        .QN(\so[26]_BAR ) );
  DFFSSRX1_RVT \q_reg[25]  ( .D(1'b0), .SETB(se), .RSTB(din[25]), .CLK(clk), 
        .QN(\so[25]_BAR ) );
  DFFSSRX1_RVT \q_reg[24]  ( .D(1'b0), .SETB(se), .RSTB(din[24]), .CLK(clk), 
        .QN(\so[24]_BAR ) );
  DFFSSRX1_RVT \q_reg[23]  ( .D(1'b0), .SETB(se), .RSTB(din[23]), .CLK(clk), 
        .QN(\so[23]_BAR ) );
  DFFSSRX1_RVT \q_reg[22]  ( .D(1'b0), .SETB(se), .RSTB(din[22]), .CLK(clk), 
        .QN(\so[22]_BAR ) );
  DFFSSRX1_RVT \q_reg[21]  ( .D(1'b0), .SETB(se), .RSTB(din[21]), .CLK(clk), 
        .QN(\so[21]_BAR ) );
  DFFSSRX1_RVT \q_reg[20]  ( .D(1'b0), .SETB(se), .RSTB(din[20]), .CLK(clk), 
        .QN(\so[20]_BAR ) );
  DFFSSRX1_RVT \q_reg[19]  ( .D(1'b0), .SETB(se), .RSTB(din[19]), .CLK(clk), 
        .QN(\so[19]_BAR ) );
  DFFSSRX1_RVT \q_reg[18]  ( .D(1'b0), .SETB(se), .RSTB(din[18]), .CLK(clk), 
        .QN(\so[18]_BAR ) );
  DFFSSRX1_RVT \q_reg[17]  ( .D(1'b0), .SETB(se), .RSTB(din[17]), .CLK(clk), 
        .QN(\so[17]_BAR ) );
  DFFSSRX1_RVT \q_reg[16]  ( .D(1'b0), .SETB(se), .RSTB(din[16]), .CLK(clk), 
        .QN(\so[16]_BAR ) );
  DFFSSRX1_RVT \q_reg[15]  ( .D(1'b0), .SETB(se), .RSTB(din[15]), .CLK(clk), 
        .QN(\so[15]_BAR ) );
  DFFSSRX1_RVT \q_reg[14]  ( .D(1'b0), .SETB(se), .RSTB(din[14]), .CLK(clk), 
        .QN(\so[14]_BAR ) );
  DFFSSRX1_RVT \q_reg[13]  ( .D(1'b0), .SETB(se), .RSTB(din[13]), .CLK(clk), 
        .QN(\so[13]_BAR ) );
  DFFSSRX1_RVT \q_reg[12]  ( .D(1'b0), .SETB(se), .RSTB(din[12]), .CLK(clk), 
        .QN(\so[12]_BAR ) );
  DFFSSRX1_RVT \q_reg[11]  ( .D(1'b0), .SETB(se), .RSTB(din[11]), .CLK(clk), 
        .QN(\so[11]_BAR ) );
  DFFSSRX1_RVT \q_reg[10]  ( .D(1'b0), .SETB(se), .RSTB(din[10]), .CLK(clk), 
        .QN(\so[10]_BAR ) );
  DFFSSRX1_RVT \q_reg[9]  ( .D(1'b0), .SETB(se), .RSTB(din[9]), .CLK(clk), 
        .QN(\so[9]_BAR ) );
  DFFSSRX1_RVT \q_reg[8]  ( .D(1'b0), .SETB(se), .RSTB(din[8]), .CLK(clk), 
        .QN(\so[8]_BAR ) );
  DFFSSRX1_RVT \q_reg[7]  ( .D(1'b0), .SETB(se), .RSTB(din[7]), .CLK(clk), 
        .QN(\so[7]_BAR ) );
  DFFSSRX1_RVT \q_reg[6]  ( .D(1'b0), .SETB(se), .RSTB(din[6]), .CLK(clk), 
        .QN(\so[6]_BAR ) );
  DFFSSRX1_RVT \q_reg[52]  ( .D(1'b0), .SETB(se), .RSTB(din[52]), .CLK(clk), 
        .QN(\so[52]_BAR ) );
  DFFSSRX1_RVT \q_reg[51]  ( .D(1'b0), .SETB(se), .RSTB(din[51]), .CLK(clk), 
        .QN(\so[51]_BAR ) );
  DFFSSRX1_RVT \q_reg[29]  ( .D(1'b0), .SETB(se), .RSTB(din[29]), .CLK(clk), 
        .QN(\so[29]_BAR ) );
  DFFSSRX1_RVT \q_reg[31]  ( .D(1'b0), .SETB(se), .RSTB(din[31]), .CLK(clk), 
        .QN(\so[31]_BAR ) );
  DFFSSRX1_RVT \q_reg[30]  ( .D(1'b0), .SETB(se), .RSTB(din[30]), .CLK(clk), 
        .QN(\so[30]_BAR ) );
  DFFSSRX1_RVT \q_reg[50]  ( .D(1'b0), .SETB(se), .RSTB(din[50]), .CLK(clk), 
        .QN(\so[50]_BAR ) );
  DFFSSRX1_RVT \q_reg[49]  ( .D(1'b0), .SETB(se), .RSTB(din[49]), .CLK(clk), 
        .QN(\so[49]_BAR ) );
  DFFSSRX1_RVT \q_reg[48]  ( .D(1'b0), .SETB(se), .RSTB(din[48]), .CLK(clk), 
        .QN(\so[48]_BAR ) );
  DFFSSRX1_RVT \q_reg[47]  ( .D(1'b0), .SETB(se), .RSTB(din[47]), .CLK(clk), 
        .QN(\so[47]_BAR ) );
  DFFSSRX1_RVT \q_reg[46]  ( .D(1'b0), .SETB(se), .RSTB(din[46]), .CLK(clk), 
        .QN(\so[46]_BAR ) );
  DFFSSRX1_RVT \q_reg[45]  ( .D(1'b0), .SETB(se), .RSTB(din[45]), .CLK(clk), 
        .QN(\so[45]_BAR ) );
  DFFSSRX1_RVT \q_reg[44]  ( .D(1'b0), .SETB(se), .RSTB(din[44]), .CLK(clk), 
        .QN(\so[44]_BAR ) );
  DFFSSRX1_RVT \q_reg[43]  ( .D(1'b0), .SETB(se), .RSTB(din[43]), .CLK(clk), 
        .QN(\so[43]_BAR ) );
  DFFSSRX1_RVT \q_reg[42]  ( .D(1'b0), .SETB(se), .RSTB(din[42]), .CLK(clk), 
        .QN(\so[42]_BAR ) );
  DFFSSRX1_RVT \q_reg[41]  ( .D(1'b0), .SETB(se), .RSTB(din[41]), .CLK(clk), 
        .QN(\so[41]_BAR ) );
  DFFSSRX1_RVT \q_reg[40]  ( .D(1'b0), .SETB(se), .RSTB(din[40]), .CLK(clk), 
        .QN(\so[40]_BAR ) );
  DFFSSRX1_RVT \q_reg[39]  ( .D(1'b0), .SETB(se), .RSTB(din[39]), .CLK(clk), 
        .QN(\so[39]_BAR ) );
  DFFSSRX1_RVT \q_reg[38]  ( .D(1'b0), .SETB(se), .RSTB(din[38]), .CLK(clk), 
        .QN(\so[38]_BAR ) );
  DFFSSRX1_RVT \q_reg[37]  ( .D(1'b0), .SETB(se), .RSTB(din[37]), .CLK(clk), 
        .QN(\so[37]_BAR ) );
  DFFSSRX1_RVT \q_reg[36]  ( .D(1'b0), .SETB(se), .RSTB(din[36]), .CLK(clk), 
        .QN(\so[36]_BAR ) );
  DFFSSRX1_RVT \q_reg[35]  ( .D(1'b0), .SETB(se), .RSTB(din[35]), .CLK(clk), 
        .QN(\so[35]_BAR ) );
  DFFSSRX1_RVT \q_reg[34]  ( .D(1'b0), .SETB(se), .RSTB(din[34]), .CLK(clk), 
        .QN(\so[34]_BAR ) );
  DFFSSRX1_RVT \q_reg[33]  ( .D(1'b0), .SETB(se), .RSTB(din[33]), .CLK(clk), 
        .QN(\so[33]_BAR ) );
  DFFSSRX1_RVT \q_reg[32]  ( .D(1'b0), .SETB(se), .RSTB(din[32]), .CLK(clk), 
        .QN(\so[32]_BAR ) );
  INVX1_RVT U56 ( .A(se), .Y(n54) );
endmodule


module dff_SIZE78_0 ( din, clk, q, se, si, so );
  input [77:0] din;
  output [77:0] q;
  input [77:0] si;
  output [77:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, n1;
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  AND2X1_RVT U3 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  INVX1_RVT U11 ( .A(se), .Y(n1) );
  AND2X1_RVT U12 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U13 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U14 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U15 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U16 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U41 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U42 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U61 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U62 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U63 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U64 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U65 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U66 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U67 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U68 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U69 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U70 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U71 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U72 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U73 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U74 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U75 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U76 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
  AND2X1_RVT U78 ( .A1(din[74]), .A2(n1), .Y(N77) );
  AND2X1_RVT U79 ( .A1(din[75]), .A2(n1), .Y(N78) );
endmodule


module dff_SIZE82_0 ( din, clk, q, se, si, so );
  input [81:0] din;
  output [81:0] q;
  input [81:0] si;
  output [81:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, n1;
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  DFFX1_RVT \q_reg[80]  ( .D(n1), .CLK(clk), .Q(q[80]) );
  DFFX1_RVT \q_reg[79]  ( .D(N82), .CLK(clk), .Q(q[79]) );
  DFFX1_RVT \q_reg[78]  ( .D(N81), .CLK(clk), .Q(q[78]) );
  DFFX1_RVT \q_reg[77]  ( .D(N80), .CLK(clk), .Q(q[77]) );
  DFFX1_RVT \q_reg[76]  ( .D(N79), .CLK(clk), .Q(q[76]) );
  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
  AND2X1_RVT U78 ( .A1(din[74]), .A2(n1), .Y(N77) );
  AND2X1_RVT U79 ( .A1(din[75]), .A2(n1), .Y(N78) );
  AND2X1_RVT U80 ( .A1(din[76]), .A2(n1), .Y(N79) );
  AND2X1_RVT U81 ( .A1(din[77]), .A2(n1), .Y(N80) );
  AND2X1_RVT U82 ( .A1(din[78]), .A2(n1), .Y(N81) );
  AND2X1_RVT U83 ( .A1(din[79]), .A2(n1), .Y(N82) );
endmodule


module dff_SIZE78_1 ( din, clk, q, se, si, so );
  input [77:0] din;
  output [77:0] q;
  input [77:0] si;
  output [77:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, n1;
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
  AND2X1_RVT U78 ( .A1(din[74]), .A2(n1), .Y(N77) );
  AND2X1_RVT U79 ( .A1(din[75]), .A2(n1), .Y(N78) );
endmodule


module dff_SIZE82_1 ( din, clk, q, se, si, so );
  input [81:0] din;
  output [81:0] q;
  input [81:0] si;
  output [81:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N84, n1;

  DFFX1_RVT \q_reg[81]  ( .D(N84), .CLK(clk), .Q(q[81]) );
  DFFX1_RVT \q_reg[80]  ( .D(n1), .CLK(clk), .Q(q[80]) );
  DFFX1_RVT \q_reg[79]  ( .D(N82), .CLK(clk), .Q(q[79]) );
  DFFX1_RVT \q_reg[78]  ( .D(N81), .CLK(clk), .Q(q[78]) );
  DFFX1_RVT \q_reg[77]  ( .D(N80), .CLK(clk), .Q(q[77]) );
  DFFX1_RVT \q_reg[76]  ( .D(N79), .CLK(clk), .Q(q[76]) );
  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
  AND2X1_RVT U78 ( .A1(din[74]), .A2(n1), .Y(N77) );
  AND2X1_RVT U79 ( .A1(din[75]), .A2(n1), .Y(N78) );
  AND2X1_RVT U80 ( .A1(din[76]), .A2(n1), .Y(N79) );
  AND2X1_RVT U81 ( .A1(din[77]), .A2(n1), .Y(N80) );
  AND2X1_RVT U82 ( .A1(din[78]), .A2(n1), .Y(N81) );
  AND2X1_RVT U83 ( .A1(din[79]), .A2(n1), .Y(N82) );
  AND2X1_RVT U84 ( .A1(din[81]), .A2(n1), .Y(N84) );
endmodule


module dff_SIZE97 ( din, clk, q, se, si, so );
  input [96:0] din;
  output [96:0] q;
  input [96:0] si;
  output [96:0] so;
  input clk, se;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, n1;
  assign q[72] = so[72];
  assign q[71] = so[71];
  assign q[70] = so[70];
  assign q[69] = so[69];
  assign q[68] = so[68];
  assign q[67] = so[67];
  assign q[66] = so[66];
  assign q[65] = so[65];
  assign q[64] = so[64];
  assign q[63] = so[63];
  assign q[62] = so[62];
  assign q[61] = so[61];
  assign q[60] = so[60];
  assign q[59] = so[59];
  assign q[58] = so[58];
  assign q[57] = so[57];
  assign q[56] = so[56];
  assign q[55] = so[55];
  assign q[54] = so[54];
  assign q[53] = so[53];
  assign q[52] = so[52];
  assign q[51] = so[51];
  assign q[50] = so[50];
  assign q[49] = so[49];
  assign q[48] = so[48];
  assign q[47] = so[47];
  assign q[46] = so[46];
  assign q[45] = so[45];
  assign q[44] = so[44];
  assign q[43] = so[43];
  assign q[42] = so[42];
  assign q[41] = so[41];
  assign q[40] = so[40];
  assign q[39] = so[39];
  assign q[38] = so[38];
  assign q[37] = so[37];
  assign q[36] = so[36];
  assign q[35] = so[35];
  assign q[34] = so[34];
  assign q[33] = so[33];
  assign q[32] = so[32];
  assign q[31] = so[31];
  assign q[30] = so[30];
  assign q[29] = so[29];
  assign q[28] = so[28];
  assign q[27] = so[27];
  assign q[26] = so[26];
  assign q[25] = so[25];
  assign q[24] = so[24];
  assign q[23] = so[23];
  assign q[22] = so[22];
  assign q[21] = so[21];
  assign q[20] = so[20];
  assign q[19] = so[19];
  assign q[18] = so[18];
  assign q[17] = so[17];
  assign q[16] = so[16];
  assign q[14] = so[14];
  assign q[13] = so[13];
  assign q[12] = so[12];
  assign q[11] = so[11];
  assign q[10] = so[10];
  assign q[9] = so[9];
  assign q[8] = so[8];
  assign q[7] = so[7];
  assign q[6] = so[6];
  assign q[5] = so[5];
  assign q[4] = so[4];
  assign q[3] = so[3];
  assign q[2] = so[2];

  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(so[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(so[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(so[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(so[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(so[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(so[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(so[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(so[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(so[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(so[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(so[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(so[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(so[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(so[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(so[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(so[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(so[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(so[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(so[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(so[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(so[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(so[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(so[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(so[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(so[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(so[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(so[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(so[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(so[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(so[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(so[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(so[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(so[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(so[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(so[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(so[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(so[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(so[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(so[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(so[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(so[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(so[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(so[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(so[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(so[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(so[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(so[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(so[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(so[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(so[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(so[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(so[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(so[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(so[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(so[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(so[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(so[16]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(so[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(so[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(so[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(so[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(so[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(so[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(so[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(so[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(so[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(so[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(so[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(so[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(so[2]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U16 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U17 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U18 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U19 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U20 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U21 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U22 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U23 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U24 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U25 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U26 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U27 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U28 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U29 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U30 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U31 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U32 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U33 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U34 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U35 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U36 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U37 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U38 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U39 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U40 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U41 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U42 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U43 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U44 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U45 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U46 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U47 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U48 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U49 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U50 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U51 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U52 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U53 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U54 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U55 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U56 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U57 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U58 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U59 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U60 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U61 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U62 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U63 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U64 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U65 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U66 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U67 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U68 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U69 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U70 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U71 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U72 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U73 ( .A1(din[72]), .A2(n1), .Y(N75) );
endmodule


module dff_SIZE98 ( din, clk, q, se, si, so );
  input [97:0] din;
  output [97:0] q;
  input [97:0] si;
  output [97:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, n1;

  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
endmodule


module dff_SIZE68 ( din, clk, q, se, si, so );
  input [67:0] din;
  output [67:0] q;
  input [67:0] si;
  output [67:0] so;
  input clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, n1;

  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U16 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U28 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U29 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U30 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U31 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U32 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U33 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U34 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U35 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U36 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U37 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U38 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U39 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U40 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U41 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U42 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U43 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U44 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U45 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U46 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U47 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U48 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U49 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U50 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U51 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U52 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U53 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U54 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U55 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U56 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U57 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U58 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U59 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U60 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U61 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U62 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U63 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U64 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U65 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U66 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U67 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U68 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U69 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U70 ( .A1(din[67]), .A2(n1), .Y(N70) );
endmodule


module dff_SIZE69 ( din, clk, q, se, si, so );
  input [68:0] din;
  output [68:0] q;
  input [68:0] si;
  output [68:0] so;
  input clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, n1;

  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U16 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U28 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U29 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U30 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U31 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U32 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U33 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U34 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U35 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U36 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U37 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U38 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U39 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U40 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U41 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U42 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U43 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U44 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U45 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U46 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U47 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U48 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U49 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U50 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U51 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U52 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U53 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U54 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U55 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U56 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U57 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U58 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U59 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U60 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U61 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U62 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U63 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U64 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U65 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U66 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U67 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U68 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U69 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U70 ( .A1(din[67]), .A2(n1), .Y(N70) );
endmodule


module dff_SIZE1_29 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE104 ( din, clk, q, se, si, so );
  input [103:0] din;
  output [103:0] q;
  input [103:0] si;
  output [103:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, n1;

  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[71]  ( .D(N74), .CLK(clk), .Q(q[71]) );
  DFFX1_RVT \q_reg[70]  ( .D(N73), .CLK(clk), .Q(q[70]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[64]  ( .D(N67), .CLK(clk), .Q(q[64]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[32]), .A2(n1), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[33]), .A2(n1), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[34]), .A2(n1), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[35]), .A2(n1), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[36]), .A2(n1), .Y(N39) );
  AND2X1_RVT U41 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U42 ( .A1(din[38]), .A2(n1), .Y(N41) );
  AND2X1_RVT U43 ( .A1(din[39]), .A2(n1), .Y(N42) );
  AND2X1_RVT U44 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U45 ( .A1(din[41]), .A2(n1), .Y(N44) );
  AND2X1_RVT U46 ( .A1(din[42]), .A2(n1), .Y(N45) );
  AND2X1_RVT U47 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U48 ( .A1(din[44]), .A2(n1), .Y(N47) );
  AND2X1_RVT U49 ( .A1(din[45]), .A2(n1), .Y(N48) );
  AND2X1_RVT U50 ( .A1(din[46]), .A2(n1), .Y(N49) );
  AND2X1_RVT U51 ( .A1(din[47]), .A2(n1), .Y(N50) );
  AND2X1_RVT U52 ( .A1(din[48]), .A2(n1), .Y(N51) );
  AND2X1_RVT U53 ( .A1(din[49]), .A2(n1), .Y(N52) );
  AND2X1_RVT U54 ( .A1(din[50]), .A2(n1), .Y(N53) );
  AND2X1_RVT U55 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U56 ( .A1(din[52]), .A2(n1), .Y(N55) );
  AND2X1_RVT U57 ( .A1(din[53]), .A2(n1), .Y(N56) );
  AND2X1_RVT U58 ( .A1(din[54]), .A2(n1), .Y(N57) );
  AND2X1_RVT U59 ( .A1(din[55]), .A2(n1), .Y(N58) );
  AND2X1_RVT U60 ( .A1(din[56]), .A2(n1), .Y(N59) );
  AND2X1_RVT U61 ( .A1(din[57]), .A2(n1), .Y(N60) );
  AND2X1_RVT U62 ( .A1(din[58]), .A2(n1), .Y(N61) );
  AND2X1_RVT U63 ( .A1(din[59]), .A2(n1), .Y(N62) );
  AND2X1_RVT U64 ( .A1(din[60]), .A2(n1), .Y(N63) );
  AND2X1_RVT U65 ( .A1(din[61]), .A2(n1), .Y(N64) );
  AND2X1_RVT U66 ( .A1(din[62]), .A2(n1), .Y(N65) );
  AND2X1_RVT U67 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U68 ( .A1(din[64]), .A2(n1), .Y(N67) );
  AND2X1_RVT U69 ( .A1(din[65]), .A2(n1), .Y(N68) );
  AND2X1_RVT U70 ( .A1(din[66]), .A2(n1), .Y(N69) );
  AND2X1_RVT U71 ( .A1(din[67]), .A2(n1), .Y(N70) );
  AND2X1_RVT U72 ( .A1(din[68]), .A2(n1), .Y(N71) );
  AND2X1_RVT U73 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U74 ( .A1(din[70]), .A2(n1), .Y(N73) );
  AND2X1_RVT U75 ( .A1(din[71]), .A2(n1), .Y(N74) );
  AND2X1_RVT U76 ( .A1(din[72]), .A2(n1), .Y(N75) );
  AND2X1_RVT U77 ( .A1(din[73]), .A2(n1), .Y(N76) );
endmodule


module dff_SIZE32_0 ( din, clk, q, se, si, so );
  input [31:0] din;
  output [31:0] q;
  input [31:0] si;
  output [31:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, n1;

  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n1), .Y(N15) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n1), .Y(N16) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n1), .Y(N17) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n1), .Y(N18) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n1), .Y(N19) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n1), .Y(N20) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n1), .Y(N21) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n1), .Y(N22) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n1), .Y(N23) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n1), .Y(N24) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n1), .Y(N25) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n1), .Y(N26) );
  AND2X1_RVT U28 ( .A1(din[24]), .A2(n1), .Y(N27) );
  AND2X1_RVT U29 ( .A1(din[25]), .A2(n1), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[26]), .A2(n1), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[27]), .A2(n1), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[28]), .A2(n1), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[29]), .A2(n1), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[30]), .A2(n1), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[31]), .A2(n1), .Y(N34) );
endmodule


module mul64 ( rs1_l, rs2, valid, areg, accreg, x2, out, rclk, si, so, se, 
        mul_rst_l, mul_step );
  input [63:0] rs1_l;
  input [63:0] rs2;
  input [96:0] areg;
  input [135:129] accreg;
  output [135:0] out;
  input valid, x2, rclk, si, se, mul_rst_l, mul_step;
  output so;
  wire   clk_enb0, cyc1, cyc2, cyc3, clk_enb1, add_cin, addin_cin, n76, n78,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n515, n516, net210935, net210936, net210937,
         net210938, net210939, net210940, net210941, net210942, net210943,
         net210944, net210945, net210946, net210947, net210948, net210949,
         net210950, net210951, net210952, net210953, net210954, net210955,
         net210956, net210957, net210958, net210959, net210960, net210961,
         net210962, net210963, net210964, net210965, net210966, net210967,
         net210968, net210969, net210970, net210971, net210972, net210973,
         net210974, net210975, net210976, net210977, net210978, net210979,
         net210980, net210981, net210982, net210983, net210984, net210985,
         net210986, net210987, net210988, net210989, net210990, net210991,
         net210992, net210993, net210994, net210995, net210996, net210997,
         net210998, net210999, net211000, net211001, net211002, net211003,
         net211004, net211005, net211006, net211007, net211008, net211009,
         net211010, net211011, net211012, net211013, net211014, net211015,
         net211016, net211017, net211018, net211019, net211020, net211021,
         net211022, net211023, net211024, net211025, net211026, net211027,
         net211028, net211029, net211030, net211031, net211032, net211033,
         net211034, net211035, net211036, net211037, net211038, net211039,
         net211040, net211041, net211042, net211043, net211044, net211045,
         net211046, net211047, net211048, net211049, net211050, net211051,
         net211052, net211053, net211054, net211055, net211056, net211057,
         net211058, net211059, net211060, net211061, net211062, net211063,
         net211064, net211065, net211066, net211067, net211068, net211069,
         net211070, net211071, net211072, net211073, net211074, net211075,
         net211076, net211077, net211078, net211079, net211080, net211081,
         net211082, net211083, net211084, net211085, net211086, net211087,
         net211088, net211089, net211090, net211091, net211092, net211093,
         net211094, net211095, net211096, net211097, net211098, net211099,
         net211100, net211101, net211102, net211103, net211104;
  wire   [63:0] op1_l;
  wire   [2:0] b0;
  wire   [2:0] b1;
  wire   [2:0] b2;
  wire   [2:0] b3;
  wire   [2:0] b4;
  wire   [2:0] b5;
  wire   [2:0] b6;
  wire   [2:0] b7;
  wire   [2:0] b8;
  wire   [2:0] b9;
  wire   [2:0] b10;
  wire   [2:0] b11;
  wire   [2:0] b12;
  wire   [2:0] b13;
  wire   [2:0] b14;
  wire   [2:0] b15;
  wire   [81:4] a0cout;
  wire   [81:0] a0sum;
  wire   [81:4] a0c;
  wire   [81:0] a0s;
  wire   [81:4] a1cout;
  wire   [81:0] a1sum;
  wire   [81:4] a1c;
  wire   [81:0] a1s;
  wire   [98:0] pcout;
  wire   [98:0] psum;
  wire   [98:30] pc;
  wire   [98:31] ps;
  wire   [96:0] ary2_cout;
  wire   [96:0] addin_cout;
  wire   [97:0] ary2_sum;
  wire   [97:0] addin_sum;
  wire   [98:31] psum_in;
  wire   [98:30] pcout_in;
  wire   [103:0] addout;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151;
  assign so = 1'b0;

  clken_buf_7 ckbuf_0 ( .clk(clk_enb0), .rclk(rclk), .enb_l(n515), .tmb_l(n516) );
  dffr_SIZE1_9 cyc1_dff ( .din(valid), .clk(clk_enb0), .rst(n78), .q(cyc1), 
        .se(se), .si(1'b0) );
  dffr_SIZE1_8 cyc2_dff ( .din(cyc1), .clk(clk_enb0), .rst(n78), .q(cyc2), 
        .se(se), .si(1'b0) );
  dffr_SIZE1_7 cyc3_dff ( .din(cyc2), .clk(clk_enb0), .rst(n78), .q(cyc3), 
        .se(se), .si(1'b0) );
  clken_buf_6 ckbuf_1 ( .clk(clk_enb1), .rclk(rclk), .enb_l(n76), .tmb_l(n516)
         );
  dff_SIZE64_1 ffrs1 ( .din({net211094, net211095, net211096, net211097, 
        net211098, net211099, net211100, net211101, net211102, net211103, 
        net211104, rs1_l[52:0]}), .clk(clk_enb1), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .\q[63]_BAR (op1_l[63]), .\q[62]_BAR (op1_l[62]), 
        .\q[61]_BAR (op1_l[61]), .\q[60]_BAR (op1_l[60]), .\q[59]_BAR (
        op1_l[59]), .\q[58]_BAR (op1_l[58]), .\q[57]_BAR (op1_l[57]), 
        .\q[56]_BAR (op1_l[56]), .\q[55]_BAR (op1_l[55]), .\q[54]_BAR (
        op1_l[54]), .\q[53]_BAR (op1_l[53]), .\q[52]_BAR (op1_l[52]), 
        .\q[51]_BAR (op1_l[51]), .\q[50]_BAR (op1_l[50]), .\q[49]_BAR (
        op1_l[49]), .\q[48]_BAR (op1_l[48]), .\q[47]_BAR (op1_l[47]), 
        .\q[46]_BAR (op1_l[46]), .\q[45]_BAR (op1_l[45]), .\q[44]_BAR (
        op1_l[44]), .\q[43]_BAR (op1_l[43]), .\q[42]_BAR (op1_l[42]), 
        .\q[41]_BAR (op1_l[41]), .\q[40]_BAR (op1_l[40]), .\q[39]_BAR (
        op1_l[39]), .\q[38]_BAR (op1_l[38]), .\q[37]_BAR (op1_l[37]), 
        .\q[36]_BAR (op1_l[36]), .\q[35]_BAR (op1_l[35]), .\q[34]_BAR (
        op1_l[34]), .\q[33]_BAR (op1_l[33]), .\q[32]_BAR (op1_l[32]), 
        .\q[31]_BAR (op1_l[31]), .\q[30]_BAR (op1_l[30]), .\q[29]_BAR (
        op1_l[29]), .\q[28]_BAR (op1_l[28]), .\q[27]_BAR (op1_l[27]), 
        .\q[26]_BAR (op1_l[26]), .\q[25]_BAR (op1_l[25]), .\q[24]_BAR (
        op1_l[24]), .\q[23]_BAR (op1_l[23]), .\q[22]_BAR (op1_l[22]), 
        .\q[21]_BAR (op1_l[21]), .\q[20]_BAR (op1_l[20]), .\q[19]_BAR (
        op1_l[19]), .\q[18]_BAR (op1_l[18]), .\q[17]_BAR (op1_l[17]), 
        .\q[16]_BAR (op1_l[16]), .\q[15]_BAR (op1_l[15]), .\q[14]_BAR (
        op1_l[14]), .\q[13]_BAR (op1_l[13]), .\q[12]_BAR (op1_l[12]), 
        .\q[11]_BAR (op1_l[11]), .\q[10]_BAR (op1_l[10]), .\q[9]_BAR (op1_l[9]), .\q[8]_BAR (op1_l[8]), .\q[7]_BAR (op1_l[7]), .\q[6]_BAR (op1_l[6]), 
        .\q[5]_BAR (op1_l[5]), .\q[4]_BAR (op1_l[4]), .\q[3]_BAR (op1_l[3]), 
        .\q[2]_BAR (op1_l[2]), .\q[1]_BAR (op1_l[1]), .\q[0]_BAR (op1_l[0]) );
  mul_booth booth ( .head(valid), .b_in({net211083, net211084, net211085, 
        net211086, net211087, net211088, net211089, net211090, net211091, 
        net211092, net211093, rs2[52:0]}), .b0(b0), .b1(b1), .b2(b2), .b3(b3), 
        .b4(b4), .b5(b5), .b6(b6), .b7(b7), .b8(b8), .b9(b9), .b10(b10), .b11(
        b11), .b12(b12), .b13(b13), .b14(b14), .b15(b15), .clk(rclk), .se(se), 
        .si(1'b0), .mul_step(mul_step), .tm_l(n516) );
  mul_array1_0 ary1_a0 ( .cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, a0cout[79:4]}), .sum({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, a0sum[79:0]}), .a({op1_l[59], op1_l[62:61], 
        op1_l[59], op1_l[59:0]}), .b0(b0), .b1(b1), .b2(b2), .b3(b3), .b4(b4), 
        .b5(b5), .b6(b6), .b7(b7), .b8({1'b0, 1'b0, 1'b0}), .bot(1'b0), .head(
        cyc1) );
  dff_SIZE78_0 a0cot_dff ( .din({net211081, net211082, a0cout[79:4]}), .clk(
        clk_enb0), .q({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        a0c[79:4]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE82_0 a0sum_dff ( .din({net211079, net211080, a0sum[79:0]}), .clk(
        clk_enb0), .q({SYNOPSYS_UNCONNECTED__6, a0s[80:0]}), .se(se), .si({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  mul_array1_1 ary1_a1 ( .cout({SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, a1cout[79:4]}), .sum({a1sum[81], 
        SYNOPSYS_UNCONNECTED__9, a1sum[79:0]}), .a({op1_l[63:62], op1_l[60], 
        op1_l[62:61], op1_l[58:54], op1_l[58], op1_l[52:0]}), .b0(b8), .b1(b9), 
        .b2(b10), .b3(b11), .b4(b12), .b5(b13), .b6(b14), .b7(b15), .b8({1'b0, 
        net211078, 1'b0}), .bot(cyc2), .head(1'b0) );
  dff_SIZE78_1 a1cot_dff ( .din({net211076, net211077, a1cout[79:4]}), .clk(
        clk_enb0), .q({SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        a1c[79:4]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE82_1 a1sum_dff ( .din({a1sum[81], net211075, a1sum[79:0]}), .clk(
        clk_enb0), .q(a1s), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  mul_array2 array2 ( .pcout({SYNOPSYS_UNCONNECTED__12, pcout[97:16], 
        SYNOPSYS_UNCONNECTED__13, pcout[14:2], SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15}), .psum({SYNOPSYS_UNCONNECTED__16, 
        psum[97:0]}), .a0c({net210970, net210971, a0c[79:4]}), .a0s({net210972, 
        a0s[80:0]}), .a1c({net210973, net210974, a1c[79:4]}), .a1s(a1s), 
        .areg({net210975, net210976, net210977, net210978, net210979, 
        net210980, net210981, net210982, net210983, net210984, net210985, 
        net210986, net210987, net210988, net210989, net210990, net210991, 
        net210992, net210993, net210994, net210995, net210996, net210997, 
        net210998, net210999, net211000, net211001, net211002, net211003, 
        net211004, net211005, net211006, net211007, net211008, net211009, 
        net211010, net211011, net211012, net211013, net211014, net211015, 
        net211016, net211017, net211018, net211019, net211020, net211021, 
        net211022, net211023, net211024, net211025, net211026, net211027, 
        net211028, net211029, net211030, net211031, net211032, net211033, 
        net211034, net211035, net211036, net211037, net211038, net211039, 
        net211040, net211041, net211042, net211043, net211044, net211045, 
        net211046, net211047, net211048, net211049, net211050, net211051, 
        net211052, net211053, net211054, net211055, net211056, net211057, 
        net211058, net211059, net211060, net211061, net211062, net211063, 
        net211064, net211065, net211066, net211067, net211068, net211069, 
        net211070, net211071}), .bot(cyc3), .pc({net211072, pc[97:31], 
        net211073}), .ps({ps[98:32], net211074}), .x2(1'b0) );
  dp_mux2es_SIZE97 ary2_cmux ( .dout({SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, ary2_cout[72:16], SYNOPSYS_UNCONNECTED__41, 
        ary2_cout[14:2], SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43}), 
        .in0({pcout[96:16], net210963, pcout[14:2], net210964, net210965}), 
        .in1({pcout[95:16], net210966, pcout[14:2], net210967, net210968, 
        net210969}), .sel(1'b0) );
  dff_SIZE97 a2cot_dff ( .din({net210936, net210937, net210938, net210939, 
        net210940, net210941, net210942, net210943, net210944, net210945, 
        net210946, net210947, net210948, net210949, net210950, net210951, 
        net210952, net210953, net210954, net210955, net210956, net210957, 
        net210958, net210959, ary2_cout[72:16], net210960, ary2_cout[14:2], 
        net210961, net210962}), .clk(clk_enb0), .q({SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, addin_cout[72:16], SYNOPSYS_UNCONNECTED__68, 
        addin_cout[14:2], SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70}), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dp_mux2es_SIZE98 ary2_smux ( .dout({SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, ary2_sum[73:0]}), .in0(psum[97:0]), .in1({
        psum[96:0], net210935}), .sel(1'b0) );
  dff_SIZE98 a2sum_dff ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, ary2_sum[73:0]}), .clk(clk_enb0), .q({
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, addin_sum[73:0]}), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE68 psum_dff ( .din({psum_in[98:32], 1'b0}), .clk(clk_enb0), .q({
        ps[98:32], SYNOPSYS_UNCONNECTED__119}), .se(se), .si({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE69 pcout_dff ( .din({1'b0, pcout_in[97:31], 1'b0}), .clk(clk_enb0), 
        .q({SYNOPSYS_UNCONNECTED__120, pc[97:31], SYNOPSYS_UNCONNECTED__121}), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE1_29 co31_dff ( .din(add_cin), .clk(clk_enb0), .q(addin_cin), .se(se), .si(1'b0) );
  dff_SIZE104 out_dff ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        addout[73:1], n1}), .clk(clk_enb0), .q({SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, out[105:32]}), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE32_0 pip_dff ( .din(out[63:32]), .clk(clk_enb0), .q(out[31:0]), .se(
        se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  INVX0_RVT U2 ( .A(n275), .Y(n278) );
  INVX0_RVT U3 ( .A(n181), .Y(n186) );
  INVX0_RVT U4 ( .A(n276), .Y(n277) );
  INVX0_RVT U5 ( .A(n136), .Y(n141) );
  INVX0_RVT U6 ( .A(n346), .Y(n347) );
  INVX0_RVT U7 ( .A(n325), .Y(n326) );
  INVX0_RVT U8 ( .A(n380), .Y(n383) );
  INVX0_RVT U9 ( .A(n381), .Y(n382) );
  INVX0_RVT U10 ( .A(n254), .Y(n255) );
  INVX0_RVT U11 ( .A(n253), .Y(n256) );
  INVX0_RVT U12 ( .A(n230), .Y(n235) );
  INVX0_RVT U13 ( .A(n210), .Y(n211) );
  INVX0_RVT U14 ( .A(n209), .Y(n212) );
  INVX0_RVT U15 ( .A(n301), .Y(n304) );
  INVX0_RVT U16 ( .A(n302), .Y(n303) );
  INVX0_RVT U17 ( .A(n180), .Y(n191) );
  INVX0_RVT U18 ( .A(n160), .Y(n161) );
  INVX0_RVT U19 ( .A(n159), .Y(n162) );
  INVX0_RVT U20 ( .A(n322), .Y(n327) );
  INVX0_RVT U21 ( .A(n480), .Y(n487) );
  INVX0_RVT U22 ( .A(n274), .Y(n283) );
  INVX0_RVT U23 ( .A(n345), .Y(n348) );
  INVX0_RVT U24 ( .A(n433), .Y(n434) );
  INVX0_RVT U25 ( .A(n432), .Y(n435) );
  INVX0_RVT U26 ( .A(n402), .Y(n408) );
  INVX0_RVT U27 ( .A(n176), .Y(n114) );
  INVX0_RVT U28 ( .A(n173), .Y(n113) );
  INVX0_RVT U29 ( .A(n196), .Y(n104) );
  INVX0_RVT U30 ( .A(n193), .Y(n103) );
  INVX0_RVT U31 ( .A(n167), .Y(n116) );
  INVX0_RVT U32 ( .A(n164), .Y(n115) );
  INVX0_RVT U33 ( .A(n476), .Y(n470) );
  INVX0_RVT U34 ( .A(n205), .Y(n102) );
  INVX0_RVT U35 ( .A(n202), .Y(n101) );
  INVX0_RVT U36 ( .A(n471), .Y(n473) );
  INVX0_RVT U37 ( .A(n464), .Y(n466) );
  INVX0_RVT U38 ( .A(n459), .Y(n461) );
  INVX0_RVT U39 ( .A(n451), .Y(n453) );
  INVX0_RVT U40 ( .A(n446), .Y(n448) );
  INVX0_RVT U41 ( .A(n217), .Y(n98) );
  INVX0_RVT U42 ( .A(n214), .Y(n97) );
  INVX0_RVT U43 ( .A(n442), .Y(n436) );
  INVX0_RVT U44 ( .A(n489), .Y(n31) );
  INVX0_RVT U45 ( .A(n437), .Y(n439) );
  INVX0_RVT U46 ( .A(n481), .Y(n483) );
  INVX0_RVT U47 ( .A(n155), .Y(n120) );
  INVX0_RVT U48 ( .A(n152), .Y(n119) );
  INVX0_RVT U49 ( .A(n131), .Y(n133) );
  INVX0_RVT U50 ( .A(n146), .Y(n122) );
  INVX0_RVT U51 ( .A(n143), .Y(n121) );
  INVX0_RVT U52 ( .A(n338), .Y(n55) );
  INVX0_RVT U53 ( .A(n341), .Y(n56) );
  INVX0_RVT U54 ( .A(n270), .Y(n82) );
  INVX0_RVT U55 ( .A(n267), .Y(n81) );
  INVX0_RVT U56 ( .A(n353), .Y(n52) );
  INVX0_RVT U57 ( .A(n261), .Y(n84) );
  INVX0_RVT U58 ( .A(n258), .Y(n83) );
  INVX0_RVT U59 ( .A(n294), .Y(n69) );
  INVX0_RVT U60 ( .A(n309), .Y(n66) );
  INVX0_RVT U61 ( .A(n306), .Y(n65) );
  INVX0_RVT U62 ( .A(n315), .Y(n63) );
  INVX0_RVT U63 ( .A(n318), .Y(n64) );
  INVX0_RVT U64 ( .A(n288), .Y(n72) );
  INVX0_RVT U65 ( .A(n329), .Y(n57) );
  INVX0_RVT U66 ( .A(n285), .Y(n71) );
  INVX0_RVT U67 ( .A(n332), .Y(n58) );
  INVX0_RVT U68 ( .A(n297), .Y(n70) );
  INVX0_RVT U69 ( .A(n377), .Y(n47) );
  INVX0_RVT U70 ( .A(n223), .Y(n95) );
  INVX0_RVT U71 ( .A(n410), .Y(n412) );
  INVX0_RVT U72 ( .A(n226), .Y(n96) );
  INVX0_RVT U73 ( .A(n384), .Y(n386) );
  INVX0_RVT U74 ( .A(n395), .Y(n397) );
  INVX0_RVT U75 ( .A(n240), .Y(n90) );
  INVX0_RVT U76 ( .A(n237), .Y(n89) );
  INVX0_RVT U77 ( .A(n391), .Y(n46) );
  INVX0_RVT U78 ( .A(n482), .Y(n32) );
  INVX0_RVT U79 ( .A(n350), .Y(n51) );
  INVX0_RVT U80 ( .A(n427), .Y(n420) );
  INVX0_RVT U81 ( .A(n422), .Y(n424) );
  INVX0_RVT U82 ( .A(n358), .Y(n50) );
  INVX0_RVT U83 ( .A(n415), .Y(n409) );
  INVX0_RVT U84 ( .A(n246), .Y(n87) );
  INVX0_RVT U85 ( .A(n249), .Y(n88) );
  INVX0_RVT U86 ( .A(addin_sum[1]), .Y(n488) );
  INVX0_RVT U87 ( .A(mul_step), .Y(n515) );
  INVX0_RVT U88 ( .A(mul_rst_l), .Y(n78) );
  INVX1_RVT U89 ( .A(n396), .Y(n389) );
  INVX1_RVT U90 ( .A(addin_sum[2]), .Y(n486) );
  AND2X1_RVT U91 ( .A1(n30), .A2(n489), .Y(n1) );
  OR2X1_RVT U92 ( .A1(addin_cout[32]), .A2(addin_sum[33]), .Y(n2) );
  AND2X1_RVT U93 ( .A1(n138), .A2(n126), .Y(n3) );
  AND2X1_RVT U94 ( .A1(n112), .A2(n183), .Y(n4) );
  INVX1_RVT U95 ( .A(addin_sum[16]), .Y(n394) );
  OR2X1_RVT U96 ( .A1(addin_sum[20]), .A2(addin_cout[19]), .Y(n5) );
  OR2X1_RVT U97 ( .A1(addin_sum[18]), .A2(addin_cout[17]), .Y(n6) );
  OR2X1_RVT U98 ( .A1(addin_cout[70]), .A2(addin_sum[71]), .Y(n7) );
  OR2X1_RVT U99 ( .A1(addin_cout[68]), .A2(addin_sum[69]), .Y(n8) );
  OR2X1_RVT U100 ( .A1(addin_cout[66]), .A2(addin_sum[67]), .Y(n9) );
  OR2X1_RVT U101 ( .A1(addin_cout[60]), .A2(addin_sum[61]), .Y(n10) );
  OR2X1_RVT U102 ( .A1(addin_cout[58]), .A2(addin_sum[59]), .Y(n11) );
  OR2X1_RVT U103 ( .A1(addin_cout[56]), .A2(addin_sum[57]), .Y(n12) );
  OR2X1_RVT U104 ( .A1(addin_cout[54]), .A2(addin_sum[55]), .Y(n13) );
  OR2X1_RVT U105 ( .A1(addin_cout[50]), .A2(addin_sum[51]), .Y(n14) );
  OR2X1_RVT U106 ( .A1(addin_cout[48]), .A2(addin_sum[49]), .Y(n15) );
  OR2X1_RVT U107 ( .A1(addin_cout[46]), .A2(addin_sum[47]), .Y(n16) );
  OR2X1_RVT U108 ( .A1(addin_cout[44]), .A2(addin_sum[45]), .Y(n17) );
  OR2X1_RVT U109 ( .A1(addin_cout[42]), .A2(addin_sum[43]), .Y(n18) );
  OR2X1_RVT U110 ( .A1(addin_cout[38]), .A2(addin_sum[39]), .Y(n19) );
  OR2X1_RVT U111 ( .A1(addin_cout[36]), .A2(addin_sum[37]), .Y(n20) );
  OR2X1_RVT U112 ( .A1(addin_cout[34]), .A2(addin_sum[35]), .Y(n21) );
  OR2X1_RVT U113 ( .A1(addin_cout[31]), .A2(addin_sum[32]), .Y(n22) );
  OR2X1_RVT U114 ( .A1(addin_sum[65]), .A2(addin_cout[64]), .Y(n23) );
  OR2X1_RVT U115 ( .A1(addin_sum[63]), .A2(addin_cout[62]), .Y(n24) );
  OR2X1_RVT U116 ( .A1(addin_sum[53]), .A2(addin_cout[52]), .Y(n25) );
  OR2X1_RVT U117 ( .A1(addin_sum[41]), .A2(addin_cout[40]), .Y(n26) );
  AO21X1_RVT U118 ( .A1(n112), .A2(n182), .A3(n111), .Y(n27) );
  AO21X1_RVT U119 ( .A1(n126), .A2(n137), .A3(n125), .Y(n28) );
  OR2X1_RVT U120 ( .A1(addin_sum[73]), .A2(addin_cout[72]), .Y(n29) );
  OR2X1_RVT U121 ( .A1(addin_sum[0]), .A2(addin_cin), .Y(n30) );
  NOR2X0_RVT U146 ( .A1(addin_cout[71]), .A2(addin_sum[72]), .Y(n131) );
  NOR2X0_RVT U147 ( .A1(addin_sum[64]), .A2(addin_cout[63]), .Y(n172) );
  INVX1_RVT U148 ( .A(n172), .Y(n177) );
  NAND2X0_RVT U149 ( .A1(n177), .A2(n23), .Y(n159) );
  NOR2X0_RVT U150 ( .A1(addin_cout[65]), .A2(addin_sum[66]), .Y(n163) );
  INVX1_RVT U151 ( .A(n163), .Y(n168) );
  NAND2X0_RVT U152 ( .A1(n9), .A2(n168), .Y(n118) );
  NOR2X0_RVT U153 ( .A1(n159), .A2(n118), .Y(n138) );
  NOR2X0_RVT U154 ( .A1(addin_cout[69]), .A2(addin_sum[70]), .Y(n142) );
  INVX1_RVT U155 ( .A(n142), .Y(n147) );
  NAND2X0_RVT U156 ( .A1(n7), .A2(n147), .Y(n124) );
  NOR2X0_RVT U157 ( .A1(addin_cout[67]), .A2(addin_sum[68]), .Y(n151) );
  INVX1_RVT U158 ( .A(n151), .Y(n156) );
  NAND2X0_RVT U159 ( .A1(n8), .A2(n156), .Y(n136) );
  NOR2X0_RVT U160 ( .A1(n124), .A2(n136), .Y(n126) );
  NOR2X0_RVT U161 ( .A1(addin_sum[52]), .A2(addin_cout[51]), .Y(n245) );
  INVX1_RVT U162 ( .A(n245), .Y(n250) );
  NAND2X0_RVT U163 ( .A1(n250), .A2(n25), .Y(n230) );
  NOR2X0_RVT U164 ( .A1(addin_cout[53]), .A2(addin_sum[54]), .Y(n236) );
  INVX1_RVT U165 ( .A(n236), .Y(n241) );
  NAND2X0_RVT U166 ( .A1(n13), .A2(n241), .Y(n92) );
  NOR2X0_RVT U167 ( .A1(n230), .A2(n92), .Y(n94) );
  NOR2X0_RVT U168 ( .A1(addin_cout[49]), .A2(addin_sum[50]), .Y(n257) );
  INVX1_RVT U169 ( .A(n257), .Y(n262) );
  NAND2X0_RVT U170 ( .A1(n14), .A2(n262), .Y(n86) );
  NOR2X0_RVT U171 ( .A1(addin_cout[47]), .A2(addin_sum[48]), .Y(n266) );
  INVX1_RVT U172 ( .A(n266), .Y(n271) );
  NAND2X0_RVT U173 ( .A1(n15), .A2(n271), .Y(n253) );
  NOR2X0_RVT U174 ( .A1(n86), .A2(n253), .Y(n232) );
  NAND2X0_RVT U175 ( .A1(n94), .A2(n232), .Y(n181) );
  NOR2X0_RVT U176 ( .A1(addin_cout[61]), .A2(addin_sum[62]), .Y(n192) );
  INVX1_RVT U177 ( .A(n192), .Y(n197) );
  NAND2X0_RVT U178 ( .A1(n197), .A2(n24), .Y(n106) );
  NOR2X0_RVT U179 ( .A1(addin_cout[59]), .A2(addin_sum[60]), .Y(n201) );
  INVX1_RVT U180 ( .A(n201), .Y(n206) );
  NAND2X0_RVT U181 ( .A1(n10), .A2(n206), .Y(n180) );
  NOR2X0_RVT U182 ( .A1(n106), .A2(n180), .Y(n108) );
  NOR2X0_RVT U183 ( .A1(addin_cout[57]), .A2(addin_sum[58]), .Y(n213) );
  INVX1_RVT U184 ( .A(n213), .Y(n218) );
  NAND2X0_RVT U185 ( .A1(n11), .A2(n218), .Y(n100) );
  NOR2X0_RVT U186 ( .A1(addin_cout[55]), .A2(addin_sum[56]), .Y(n222) );
  INVX1_RVT U187 ( .A(n222), .Y(n227) );
  NAND2X0_RVT U188 ( .A1(n12), .A2(n227), .Y(n209) );
  NOR2X0_RVT U189 ( .A1(n100), .A2(n209), .Y(n188) );
  NAND2X0_RVT U190 ( .A1(n108), .A2(n188), .Y(n110) );
  NOR2X0_RVT U191 ( .A1(n181), .A2(n110), .Y(n112) );
  NOR2X0_RVT U192 ( .A1(addin_sum[40]), .A2(addin_cout[39]), .Y(n314) );
  INVX1_RVT U193 ( .A(n314), .Y(n319) );
  NAND2X0_RVT U194 ( .A1(n319), .A2(n26), .Y(n301) );
  NOR2X0_RVT U195 ( .A1(addin_cout[41]), .A2(addin_sum[42]), .Y(n305) );
  INVX1_RVT U196 ( .A(n305), .Y(n310) );
  NAND2X0_RVT U197 ( .A1(n18), .A2(n310), .Y(n68) );
  NOR2X0_RVT U198 ( .A1(n301), .A2(n68), .Y(n280) );
  NOR2X0_RVT U199 ( .A1(addin_cout[45]), .A2(addin_sum[46]), .Y(n284) );
  INVX1_RVT U200 ( .A(n284), .Y(n289) );
  NAND2X0_RVT U201 ( .A1(n16), .A2(n289), .Y(n74) );
  NOR2X0_RVT U202 ( .A1(addin_cout[43]), .A2(addin_sum[44]), .Y(n293) );
  INVX1_RVT U203 ( .A(n293), .Y(n298) );
  NAND2X0_RVT U204 ( .A1(n17), .A2(n298), .Y(n274) );
  NOR2X0_RVT U205 ( .A1(n74), .A2(n274), .Y(n77) );
  NAND2X0_RVT U206 ( .A1(n280), .A2(n77), .Y(n80) );
  NOR2X0_RVT U207 ( .A1(addin_cout[37]), .A2(addin_sum[38]), .Y(n328) );
  INVX1_RVT U208 ( .A(n328), .Y(n333) );
  NAND2X0_RVT U209 ( .A1(n19), .A2(n333), .Y(n60) );
  NOR2X0_RVT U210 ( .A1(addin_cout[35]), .A2(addin_sum[36]), .Y(n337) );
  INVX1_RVT U211 ( .A(n337), .Y(n342) );
  NAND2X0_RVT U212 ( .A1(n20), .A2(n342), .Y(n322) );
  NOR2X0_RVT U213 ( .A1(n60), .A2(n322), .Y(n62) );
  NOR2X0_RVT U214 ( .A1(addin_cout[33]), .A2(addin_sum[34]), .Y(n349) );
  INVX1_RVT U215 ( .A(n349), .Y(n354) );
  NAND2X0_RVT U216 ( .A1(n21), .A2(n354), .Y(n54) );
  NAND2X0_RVT U217 ( .A1(n2), .A2(n22), .Y(n345) );
  NOR2X0_RVT U218 ( .A1(n54), .A2(n345), .Y(n324) );
  NAND2X0_RVT U219 ( .A1(n62), .A2(n324), .Y(n275) );
  NOR2X0_RVT U220 ( .A1(n80), .A2(n275), .Y(n183) );
  NOR2X0_RVT U221 ( .A1(addin_sum[19]), .A2(addin_cout[18]), .Y(n384) );
  NOR2X0_RVT U222 ( .A1(addin_sum[17]), .A2(addin_cout[16]), .Y(n395) );
  NOR2X0_RVT U223 ( .A1(n394), .A2(n395), .Y(n390) );
  NAND2X0_RVT U224 ( .A1(n6), .A2(n390), .Y(n380) );
  NOR2X0_RVT U225 ( .A1(n384), .A2(n380), .Y(n376) );
  NAND2X0_RVT U226 ( .A1(n5), .A2(n376), .Y(n49) );
  NOR2X0_RVT U227 ( .A1(addin_cout[12]), .A2(addin_sum[13]), .Y(n422) );
  NOR2X0_RVT U228 ( .A1(addin_cout[11]), .A2(addin_sum[12]), .Y(n419) );
  NOR2X0_RVT U229 ( .A1(n422), .A2(n419), .Y(n402) );
  NOR2X0_RVT U230 ( .A1(addin_sum[15]), .A2(addin_cout[14]), .Y(n410) );
  NOR2X0_RVT U231 ( .A1(addin_cout[13]), .A2(addin_sum[14]), .Y(n401) );
  NOR2X0_RVT U232 ( .A1(n410), .A2(n401), .Y(n41) );
  NAND2X0_RVT U233 ( .A1(n402), .A2(n41), .Y(n43) );
  NOR2X0_RVT U234 ( .A1(addin_sum[11]), .A2(addin_cout[10]), .Y(n437) );
  NOR2X0_RVT U235 ( .A1(addin_sum[10]), .A2(addin_cout[9]), .Y(n431) );
  NOR2X0_RVT U236 ( .A1(n437), .A2(n431), .Y(n39) );
  NOR2X0_RVT U237 ( .A1(addin_sum[9]), .A2(addin_cout[8]), .Y(n446) );
  NOR2X0_RVT U238 ( .A1(addin_sum[8]), .A2(addin_cout[7]), .Y(n451) );
  NOR2X0_RVT U239 ( .A1(n446), .A2(n451), .Y(n432) );
  NAND2X0_RVT U240 ( .A1(n39), .A2(n432), .Y(n405) );
  NOR2X0_RVT U241 ( .A1(n43), .A2(n405), .Y(n45) );
  NOR2X0_RVT U242 ( .A1(addin_cout[3]), .A2(addin_sum[4]), .Y(n469) );
  NOR2X0_RVT U243 ( .A1(addin_cout[4]), .A2(addin_sum[5]), .Y(n471) );
  NOR2X0_RVT U244 ( .A1(n469), .A2(n471), .Y(n458) );
  NOR2X0_RVT U245 ( .A1(addin_sum[7]), .A2(addin_cout[6]), .Y(n459) );
  NOR2X0_RVT U246 ( .A1(addin_sum[6]), .A2(addin_cout[5]), .Y(n464) );
  NOR2X0_RVT U247 ( .A1(n459), .A2(n464), .Y(n35) );
  NAND2X0_RVT U248 ( .A1(n458), .A2(n35), .Y(n37) );
  NOR2X0_RVT U249 ( .A1(addin_sum[3]), .A2(addin_cout[2]), .Y(n481) );
  NOR2X0_RVT U250 ( .A1(n486), .A2(n481), .Y(n33) );
  NAND2X0_RVT U251 ( .A1(addin_sum[0]), .A2(addin_cin), .Y(n489) );
  AND2X1_RVT U252 ( .A1(addin_sum[1]), .A2(n31), .Y(n480) );
  NAND2X0_RVT U253 ( .A1(addin_sum[3]), .A2(addin_cout[2]), .Y(n482) );
  AOI21X1_RVT U254 ( .A1(n33), .A2(n480), .A3(n32), .Y(n456) );
  NAND2X0_RVT U255 ( .A1(addin_cout[3]), .A2(addin_sum[4]), .Y(n476) );
  NAND2X0_RVT U256 ( .A1(addin_cout[4]), .A2(addin_sum[5]), .Y(n472) );
  OAI21X1_RVT U257 ( .A1(n476), .A2(n471), .A3(n472), .Y(n457) );
  NAND2X0_RVT U258 ( .A1(addin_sum[6]), .A2(addin_cout[5]), .Y(n465) );
  NAND2X0_RVT U259 ( .A1(addin_sum[7]), .A2(addin_cout[6]), .Y(n460) );
  OAI21X1_RVT U260 ( .A1(n465), .A2(n459), .A3(n460), .Y(n34) );
  AOI21X1_RVT U261 ( .A1(n35), .A2(n457), .A3(n34), .Y(n36) );
  OAI21X1_RVT U262 ( .A1(n37), .A2(n456), .A3(n36), .Y(n403) );
  NAND2X0_RVT U263 ( .A1(addin_sum[8]), .A2(addin_cout[7]), .Y(n452) );
  NAND2X0_RVT U264 ( .A1(addin_sum[9]), .A2(addin_cout[8]), .Y(n447) );
  OAI21X1_RVT U265 ( .A1(n452), .A2(n446), .A3(n447), .Y(n433) );
  NAND2X0_RVT U266 ( .A1(addin_sum[10]), .A2(addin_cout[9]), .Y(n442) );
  NAND2X0_RVT U267 ( .A1(addin_sum[11]), .A2(addin_cout[10]), .Y(n438) );
  OAI21X1_RVT U268 ( .A1(n442), .A2(n437), .A3(n438), .Y(n38) );
  AOI21X1_RVT U269 ( .A1(n39), .A2(n433), .A3(n38), .Y(n404) );
  NAND2X0_RVT U270 ( .A1(addin_cout[11]), .A2(addin_sum[12]), .Y(n427) );
  NAND2X0_RVT U271 ( .A1(addin_cout[12]), .A2(addin_sum[13]), .Y(n423) );
  OAI21X1_RVT U272 ( .A1(n427), .A2(n422), .A3(n423), .Y(n406) );
  NAND2X0_RVT U273 ( .A1(addin_cout[13]), .A2(addin_sum[14]), .Y(n415) );
  NAND2X0_RVT U274 ( .A1(addin_sum[15]), .A2(addin_cout[14]), .Y(n411) );
  OAI21X1_RVT U275 ( .A1(n415), .A2(n410), .A3(n411), .Y(n40) );
  AOI21X1_RVT U276 ( .A1(n41), .A2(n406), .A3(n40), .Y(n42) );
  OAI21X1_RVT U277 ( .A1(n43), .A2(n404), .A3(n42), .Y(n44) );
  AOI21X1_RVT U278 ( .A1(n45), .A2(n403), .A3(n44), .Y(n374) );
  NAND2X0_RVT U279 ( .A1(addin_sum[17]), .A2(addin_cout[16]), .Y(n396) );
  NAND2X0_RVT U280 ( .A1(addin_sum[18]), .A2(addin_cout[17]), .Y(n391) );
  AOI21X1_RVT U281 ( .A1(n6), .A2(n389), .A3(n46), .Y(n381) );
  NAND2X0_RVT U282 ( .A1(addin_sum[19]), .A2(addin_cout[18]), .Y(n385) );
  OAI21X1_RVT U283 ( .A1(n384), .A2(n381), .A3(n385), .Y(n375) );
  NAND2X0_RVT U284 ( .A1(addin_sum[20]), .A2(addin_cout[19]), .Y(n377) );
  AOI21X1_RVT U285 ( .A1(n5), .A2(n375), .A3(n47), .Y(n48) );
  OAI21X1_RVT U286 ( .A1(n49), .A2(n374), .A3(n48), .Y(n373) );
  NAND2X0_RVT U287 ( .A1(addin_cout[31]), .A2(addin_sum[32]), .Y(n361) );
  INVX1_RVT U288 ( .A(n361), .Y(n357) );
  NAND2X0_RVT U289 ( .A1(addin_cout[32]), .A2(addin_sum[33]), .Y(n358) );
  AOI21X1_RVT U290 ( .A1(n357), .A2(n2), .A3(n50), .Y(n346) );
  NAND2X0_RVT U291 ( .A1(addin_cout[33]), .A2(addin_sum[34]), .Y(n353) );
  NAND2X0_RVT U292 ( .A1(addin_cout[34]), .A2(addin_sum[35]), .Y(n350) );
  AOI21X1_RVT U293 ( .A1(n52), .A2(n21), .A3(n51), .Y(n53) );
  OAI21X1_RVT U294 ( .A1(n54), .A2(n346), .A3(n53), .Y(n323) );
  NAND2X0_RVT U295 ( .A1(addin_cout[35]), .A2(addin_sum[36]), .Y(n341) );
  NAND2X0_RVT U296 ( .A1(addin_cout[36]), .A2(addin_sum[37]), .Y(n338) );
  AOI21X1_RVT U297 ( .A1(n56), .A2(n20), .A3(n55), .Y(n325) );
  NAND2X0_RVT U298 ( .A1(addin_cout[37]), .A2(addin_sum[38]), .Y(n332) );
  NAND2X0_RVT U299 ( .A1(addin_cout[38]), .A2(addin_sum[39]), .Y(n329) );
  AOI21X1_RVT U300 ( .A1(n58), .A2(n19), .A3(n57), .Y(n59) );
  OAI21X1_RVT U301 ( .A1(n60), .A2(n325), .A3(n59), .Y(n61) );
  AOI21X1_RVT U302 ( .A1(n62), .A2(n323), .A3(n61), .Y(n276) );
  NAND2X0_RVT U303 ( .A1(addin_sum[40]), .A2(addin_cout[39]), .Y(n318) );
  NAND2X0_RVT U304 ( .A1(addin_sum[41]), .A2(addin_cout[40]), .Y(n315) );
  AOI21X1_RVT U305 ( .A1(n64), .A2(n26), .A3(n63), .Y(n302) );
  NAND2X0_RVT U306 ( .A1(addin_cout[41]), .A2(addin_sum[42]), .Y(n309) );
  NAND2X0_RVT U307 ( .A1(addin_cout[42]), .A2(addin_sum[43]), .Y(n306) );
  AOI21X1_RVT U308 ( .A1(n66), .A2(n18), .A3(n65), .Y(n67) );
  OAI21X1_RVT U309 ( .A1(n68), .A2(n302), .A3(n67), .Y(n279) );
  NAND2X0_RVT U310 ( .A1(addin_cout[43]), .A2(addin_sum[44]), .Y(n297) );
  NAND2X0_RVT U311 ( .A1(addin_cout[44]), .A2(addin_sum[45]), .Y(n294) );
  AOI21X1_RVT U312 ( .A1(n70), .A2(n17), .A3(n69), .Y(n281) );
  NAND2X0_RVT U313 ( .A1(addin_cout[45]), .A2(addin_sum[46]), .Y(n288) );
  NAND2X0_RVT U314 ( .A1(addin_cout[46]), .A2(addin_sum[47]), .Y(n285) );
  AOI21X1_RVT U315 ( .A1(n72), .A2(n16), .A3(n71), .Y(n73) );
  OAI21X1_RVT U316 ( .A1(n74), .A2(n281), .A3(n73), .Y(n75) );
  AOI21X1_RVT U317 ( .A1(n77), .A2(n279), .A3(n75), .Y(n79) );
  OAI21X1_RVT U318 ( .A1(n80), .A2(n276), .A3(n79), .Y(n182) );
  NAND2X0_RVT U319 ( .A1(addin_cout[47]), .A2(addin_sum[48]), .Y(n270) );
  NAND2X0_RVT U320 ( .A1(addin_cout[48]), .A2(addin_sum[49]), .Y(n267) );
  AOI21X1_RVT U321 ( .A1(n82), .A2(n15), .A3(n81), .Y(n254) );
  NAND2X0_RVT U322 ( .A1(addin_cout[49]), .A2(addin_sum[50]), .Y(n261) );
  NAND2X0_RVT U323 ( .A1(addin_cout[50]), .A2(addin_sum[51]), .Y(n258) );
  AOI21X1_RVT U324 ( .A1(n84), .A2(n14), .A3(n83), .Y(n85) );
  OAI21X1_RVT U325 ( .A1(n86), .A2(n254), .A3(n85), .Y(n231) );
  NAND2X0_RVT U326 ( .A1(addin_sum[52]), .A2(addin_cout[51]), .Y(n249) );
  NAND2X0_RVT U327 ( .A1(addin_sum[53]), .A2(addin_cout[52]), .Y(n246) );
  AOI21X1_RVT U328 ( .A1(n88), .A2(n25), .A3(n87), .Y(n233) );
  NAND2X0_RVT U329 ( .A1(addin_cout[53]), .A2(addin_sum[54]), .Y(n240) );
  NAND2X0_RVT U330 ( .A1(addin_cout[54]), .A2(addin_sum[55]), .Y(n237) );
  AOI21X1_RVT U331 ( .A1(n90), .A2(n13), .A3(n89), .Y(n91) );
  OAI21X1_RVT U332 ( .A1(n92), .A2(n233), .A3(n91), .Y(n93) );
  AOI21X1_RVT U333 ( .A1(n94), .A2(n231), .A3(n93), .Y(n184) );
  NAND2X0_RVT U334 ( .A1(addin_cout[55]), .A2(addin_sum[56]), .Y(n226) );
  NAND2X0_RVT U335 ( .A1(addin_cout[56]), .A2(addin_sum[57]), .Y(n223) );
  AOI21X1_RVT U336 ( .A1(n96), .A2(n12), .A3(n95), .Y(n210) );
  NAND2X0_RVT U337 ( .A1(addin_cout[57]), .A2(addin_sum[58]), .Y(n217) );
  NAND2X0_RVT U338 ( .A1(addin_cout[58]), .A2(addin_sum[59]), .Y(n214) );
  AOI21X1_RVT U339 ( .A1(n98), .A2(n11), .A3(n97), .Y(n99) );
  OAI21X1_RVT U340 ( .A1(n100), .A2(n210), .A3(n99), .Y(n187) );
  NAND2X0_RVT U341 ( .A1(addin_cout[59]), .A2(addin_sum[60]), .Y(n205) );
  NAND2X0_RVT U342 ( .A1(addin_cout[60]), .A2(addin_sum[61]), .Y(n202) );
  AOI21X1_RVT U343 ( .A1(n102), .A2(n10), .A3(n101), .Y(n189) );
  NAND2X0_RVT U344 ( .A1(addin_cout[61]), .A2(addin_sum[62]), .Y(n196) );
  NAND2X0_RVT U345 ( .A1(addin_sum[63]), .A2(addin_cout[62]), .Y(n193) );
  AOI21X1_RVT U346 ( .A1(n104), .A2(n24), .A3(n103), .Y(n105) );
  OAI21X1_RVT U347 ( .A1(n106), .A2(n189), .A3(n105), .Y(n107) );
  AOI21X1_RVT U348 ( .A1(n108), .A2(n187), .A3(n107), .Y(n109) );
  OAI21X1_RVT U349 ( .A1(n110), .A2(n184), .A3(n109), .Y(n111) );
  AOI21X1_RVT U350 ( .A1(n4), .A2(n490), .A3(n27), .Y(n171) );
  INVX1_RVT U351 ( .A(n171), .Y(n179) );
  NAND2X0_RVT U352 ( .A1(addin_sum[64]), .A2(addin_cout[63]), .Y(n176) );
  NAND2X0_RVT U353 ( .A1(addin_sum[65]), .A2(addin_cout[64]), .Y(n173) );
  AOI21X1_RVT U354 ( .A1(n114), .A2(n23), .A3(n113), .Y(n160) );
  NAND2X0_RVT U355 ( .A1(addin_cout[65]), .A2(addin_sum[66]), .Y(n167) );
  NAND2X0_RVT U356 ( .A1(addin_cout[66]), .A2(addin_sum[67]), .Y(n164) );
  AOI21X1_RVT U357 ( .A1(n116), .A2(n9), .A3(n115), .Y(n117) );
  OAI21X1_RVT U358 ( .A1(n118), .A2(n160), .A3(n117), .Y(n137) );
  NAND2X0_RVT U359 ( .A1(addin_cout[67]), .A2(addin_sum[68]), .Y(n155) );
  NAND2X0_RVT U360 ( .A1(addin_cout[68]), .A2(addin_sum[69]), .Y(n152) );
  AOI21X1_RVT U361 ( .A1(n120), .A2(n8), .A3(n119), .Y(n139) );
  NAND2X0_RVT U362 ( .A1(addin_cout[69]), .A2(addin_sum[70]), .Y(n146) );
  NAND2X0_RVT U363 ( .A1(addin_cout[70]), .A2(addin_sum[71]), .Y(n143) );
  AOI21X1_RVT U364 ( .A1(n122), .A2(n7), .A3(n121), .Y(n123) );
  OAI21X1_RVT U365 ( .A1(n124), .A2(n139), .A3(n123), .Y(n125) );
  AOI21X1_RVT U366 ( .A1(n3), .A2(n179), .A3(n28), .Y(n130) );
  NAND2X0_RVT U367 ( .A1(addin_cout[71]), .A2(addin_sum[72]), .Y(n132) );
  OAI21X1_RVT U368 ( .A1(n131), .A2(n130), .A3(n132), .Y(n129) );
  NAND2X0_RVT U369 ( .A1(addin_sum[73]), .A2(addin_cout[72]), .Y(n127) );
  NAND2X0_RVT U370 ( .A1(n29), .A2(n127), .Y(n128) );
  XNOR2X1_RVT U371 ( .A1(n129), .A2(n128), .Y(addout[73]) );
  INVX1_RVT U372 ( .A(n130), .Y(n135) );
  NAND2X0_RVT U373 ( .A1(n133), .A2(n132), .Y(n134) );
  XNOR2X1_RVT U374 ( .A1(n135), .A2(n134), .Y(addout[72]) );
  AOI21X1_RVT U375 ( .A1(n138), .A2(n179), .A3(n137), .Y(n150) );
  INVX1_RVT U376 ( .A(n150), .Y(n158) );
  INVX1_RVT U377 ( .A(n139), .Y(n140) );
  AOI21X1_RVT U378 ( .A1(n141), .A2(n158), .A3(n140), .Y(n149) );
  OAI21X1_RVT U379 ( .A1(n142), .A2(n149), .A3(n146), .Y(n145) );
  NAND2X0_RVT U380 ( .A1(n7), .A2(n143), .Y(n144) );
  XNOR2X1_RVT U381 ( .A1(n145), .A2(n144), .Y(addout[71]) );
  NAND2X0_RVT U382 ( .A1(n147), .A2(n146), .Y(n148) );
  XOR2X1_RVT U383 ( .A1(n149), .A2(n148), .Y(addout[70]) );
  OAI21X1_RVT U384 ( .A1(n151), .A2(n150), .A3(n155), .Y(n154) );
  NAND2X0_RVT U385 ( .A1(n8), .A2(n152), .Y(n153) );
  XNOR2X1_RVT U386 ( .A1(n154), .A2(n153), .Y(addout[69]) );
  NAND2X0_RVT U387 ( .A1(n156), .A2(n155), .Y(n157) );
  XNOR2X1_RVT U388 ( .A1(n158), .A2(n157), .Y(addout[68]) );
  AOI21X1_RVT U389 ( .A1(n162), .A2(n179), .A3(n161), .Y(n170) );
  OAI21X1_RVT U390 ( .A1(n163), .A2(n170), .A3(n167), .Y(n166) );
  NAND2X0_RVT U391 ( .A1(n9), .A2(n164), .Y(n165) );
  XNOR2X1_RVT U392 ( .A1(n166), .A2(n165), .Y(addout[67]) );
  NAND2X0_RVT U393 ( .A1(n168), .A2(n167), .Y(n169) );
  XOR2X1_RVT U394 ( .A1(n170), .A2(n169), .Y(addout[66]) );
  OAI21X1_RVT U395 ( .A1(n172), .A2(n171), .A3(n176), .Y(n175) );
  NAND2X0_RVT U396 ( .A1(n23), .A2(n173), .Y(n174) );
  XNOR2X1_RVT U397 ( .A1(n175), .A2(n174), .Y(addout[65]) );
  NAND2X0_RVT U398 ( .A1(n177), .A2(n176), .Y(n178) );
  XNOR2X1_RVT U399 ( .A1(n179), .A2(n178), .Y(addout[64]) );
  AOI21X1_RVT U400 ( .A1(n183), .A2(n490), .A3(n182), .Y(n265) );
  INVX1_RVT U401 ( .A(n265), .Y(n273) );
  INVX1_RVT U402 ( .A(n184), .Y(n185) );
  AOI21X1_RVT U403 ( .A1(n186), .A2(n273), .A3(n185), .Y(n221) );
  INVX1_RVT U404 ( .A(n221), .Y(n229) );
  AOI21X1_RVT U405 ( .A1(n188), .A2(n229), .A3(n187), .Y(n200) );
  INVX1_RVT U406 ( .A(n200), .Y(n208) );
  INVX1_RVT U407 ( .A(n189), .Y(n190) );
  AOI21X1_RVT U408 ( .A1(n191), .A2(n208), .A3(n190), .Y(n199) );
  OAI21X1_RVT U409 ( .A1(n192), .A2(n199), .A3(n196), .Y(n195) );
  NAND2X0_RVT U410 ( .A1(n24), .A2(n193), .Y(n194) );
  XNOR2X1_RVT U411 ( .A1(n195), .A2(n194), .Y(addout[63]) );
  NAND2X0_RVT U412 ( .A1(n197), .A2(n196), .Y(n198) );
  XOR2X1_RVT U413 ( .A1(n199), .A2(n198), .Y(addout[62]) );
  OAI21X1_RVT U414 ( .A1(n201), .A2(n200), .A3(n205), .Y(n204) );
  NAND2X0_RVT U415 ( .A1(n10), .A2(n202), .Y(n203) );
  XNOR2X1_RVT U416 ( .A1(n204), .A2(n203), .Y(addout[61]) );
  NAND2X0_RVT U417 ( .A1(n206), .A2(n205), .Y(n207) );
  XNOR2X1_RVT U418 ( .A1(n208), .A2(n207), .Y(addout[60]) );
  AOI21X1_RVT U419 ( .A1(n212), .A2(n229), .A3(n211), .Y(n220) );
  OAI21X1_RVT U420 ( .A1(n213), .A2(n220), .A3(n217), .Y(n216) );
  NAND2X0_RVT U421 ( .A1(n11), .A2(n214), .Y(n215) );
  XNOR2X1_RVT U422 ( .A1(n216), .A2(n215), .Y(addout[59]) );
  NAND2X0_RVT U423 ( .A1(n218), .A2(n217), .Y(n219) );
  XOR2X1_RVT U424 ( .A1(n220), .A2(n219), .Y(addout[58]) );
  OAI21X1_RVT U425 ( .A1(n222), .A2(n221), .A3(n226), .Y(n225) );
  NAND2X0_RVT U426 ( .A1(n12), .A2(n223), .Y(n224) );
  XNOR2X1_RVT U427 ( .A1(n225), .A2(n224), .Y(addout[57]) );
  NAND2X0_RVT U428 ( .A1(n227), .A2(n226), .Y(n228) );
  XNOR2X1_RVT U429 ( .A1(n229), .A2(n228), .Y(addout[56]) );
  AOI21X1_RVT U430 ( .A1(n232), .A2(n273), .A3(n231), .Y(n244) );
  INVX1_RVT U431 ( .A(n244), .Y(n252) );
  INVX1_RVT U432 ( .A(n233), .Y(n234) );
  AOI21X1_RVT U433 ( .A1(n235), .A2(n252), .A3(n234), .Y(n243) );
  OAI21X1_RVT U434 ( .A1(n236), .A2(n243), .A3(n240), .Y(n239) );
  NAND2X0_RVT U435 ( .A1(n13), .A2(n237), .Y(n238) );
  XNOR2X1_RVT U436 ( .A1(n239), .A2(n238), .Y(addout[55]) );
  NAND2X0_RVT U437 ( .A1(n241), .A2(n240), .Y(n242) );
  XOR2X1_RVT U438 ( .A1(n243), .A2(n242), .Y(addout[54]) );
  OAI21X1_RVT U439 ( .A1(n245), .A2(n244), .A3(n249), .Y(n248) );
  NAND2X0_RVT U440 ( .A1(n25), .A2(n246), .Y(n247) );
  XNOR2X1_RVT U441 ( .A1(n248), .A2(n247), .Y(addout[53]) );
  NAND2X0_RVT U442 ( .A1(n250), .A2(n249), .Y(n251) );
  XNOR2X1_RVT U443 ( .A1(n252), .A2(n251), .Y(addout[52]) );
  AOI21X1_RVT U444 ( .A1(n256), .A2(n273), .A3(n255), .Y(n264) );
  OAI21X1_RVT U445 ( .A1(n257), .A2(n264), .A3(n261), .Y(n260) );
  NAND2X0_RVT U446 ( .A1(n14), .A2(n258), .Y(n259) );
  XNOR2X1_RVT U447 ( .A1(n260), .A2(n259), .Y(addout[51]) );
  NAND2X0_RVT U448 ( .A1(n262), .A2(n261), .Y(n263) );
  XOR2X1_RVT U449 ( .A1(n264), .A2(n263), .Y(addout[50]) );
  OAI21X1_RVT U450 ( .A1(n266), .A2(n265), .A3(n270), .Y(n269) );
  NAND2X0_RVT U451 ( .A1(n15), .A2(n267), .Y(n268) );
  XNOR2X1_RVT U452 ( .A1(n269), .A2(n268), .Y(addout[49]) );
  NAND2X0_RVT U453 ( .A1(n271), .A2(n270), .Y(n272) );
  XNOR2X1_RVT U454 ( .A1(n273), .A2(n272), .Y(addout[48]) );
  AOI21X1_RVT U455 ( .A1(n278), .A2(n490), .A3(n277), .Y(n313) );
  INVX1_RVT U456 ( .A(n313), .Y(n321) );
  AOI21X1_RVT U457 ( .A1(n280), .A2(n321), .A3(n279), .Y(n292) );
  INVX1_RVT U458 ( .A(n292), .Y(n300) );
  INVX1_RVT U459 ( .A(n281), .Y(n282) );
  AOI21X1_RVT U460 ( .A1(n283), .A2(n300), .A3(n282), .Y(n291) );
  OAI21X1_RVT U461 ( .A1(n284), .A2(n291), .A3(n288), .Y(n287) );
  NAND2X0_RVT U462 ( .A1(n16), .A2(n285), .Y(n286) );
  XNOR2X1_RVT U463 ( .A1(n287), .A2(n286), .Y(addout[47]) );
  NAND2X0_RVT U464 ( .A1(n289), .A2(n288), .Y(n290) );
  XOR2X1_RVT U465 ( .A1(n291), .A2(n290), .Y(addout[46]) );
  OAI21X1_RVT U466 ( .A1(n293), .A2(n292), .A3(n297), .Y(n296) );
  NAND2X0_RVT U467 ( .A1(n17), .A2(n294), .Y(n295) );
  XNOR2X1_RVT U468 ( .A1(n296), .A2(n295), .Y(addout[45]) );
  NAND2X0_RVT U469 ( .A1(n298), .A2(n297), .Y(n299) );
  XNOR2X1_RVT U470 ( .A1(n300), .A2(n299), .Y(addout[44]) );
  AOI21X1_RVT U471 ( .A1(n304), .A2(n321), .A3(n303), .Y(n312) );
  OAI21X1_RVT U472 ( .A1(n305), .A2(n312), .A3(n309), .Y(n308) );
  NAND2X0_RVT U473 ( .A1(n18), .A2(n306), .Y(n307) );
  XNOR2X1_RVT U474 ( .A1(n308), .A2(n307), .Y(addout[43]) );
  NAND2X0_RVT U475 ( .A1(n310), .A2(n309), .Y(n311) );
  XOR2X1_RVT U476 ( .A1(n312), .A2(n311), .Y(addout[42]) );
  OAI21X1_RVT U477 ( .A1(n314), .A2(n313), .A3(n318), .Y(n317) );
  NAND2X0_RVT U478 ( .A1(n26), .A2(n315), .Y(n316) );
  XNOR2X1_RVT U479 ( .A1(n317), .A2(n316), .Y(addout[41]) );
  NAND2X0_RVT U480 ( .A1(n319), .A2(n318), .Y(n320) );
  XNOR2X1_RVT U481 ( .A1(n321), .A2(n320), .Y(addout[40]) );
  AOI21X1_RVT U482 ( .A1(n324), .A2(n490), .A3(n323), .Y(n336) );
  INVX1_RVT U483 ( .A(n336), .Y(n344) );
  AOI21X1_RVT U484 ( .A1(n327), .A2(n344), .A3(n326), .Y(n335) );
  OAI21X1_RVT U485 ( .A1(n328), .A2(n335), .A3(n332), .Y(n331) );
  NAND2X0_RVT U486 ( .A1(n19), .A2(n329), .Y(n330) );
  XNOR2X1_RVT U487 ( .A1(n331), .A2(n330), .Y(addout[39]) );
  NAND2X0_RVT U488 ( .A1(n333), .A2(n332), .Y(n334) );
  XOR2X1_RVT U489 ( .A1(n335), .A2(n334), .Y(addout[38]) );
  OAI21X1_RVT U490 ( .A1(n337), .A2(n336), .A3(n341), .Y(n340) );
  NAND2X0_RVT U491 ( .A1(n20), .A2(n338), .Y(n339) );
  XNOR2X1_RVT U492 ( .A1(n340), .A2(n339), .Y(addout[37]) );
  NAND2X0_RVT U493 ( .A1(n342), .A2(n341), .Y(n343) );
  XNOR2X1_RVT U494 ( .A1(n344), .A2(n343), .Y(addout[36]) );
  AOI21X1_RVT U495 ( .A1(n348), .A2(n490), .A3(n347), .Y(n356) );
  OAI21X1_RVT U496 ( .A1(n349), .A2(n356), .A3(n353), .Y(n352) );
  NAND2X0_RVT U497 ( .A1(n21), .A2(n350), .Y(n351) );
  XNOR2X1_RVT U498 ( .A1(n352), .A2(n351), .Y(addout[35]) );
  NAND2X0_RVT U499 ( .A1(n354), .A2(n353), .Y(n355) );
  XOR2X1_RVT U500 ( .A1(n356), .A2(n355), .Y(addout[34]) );
  AOI21X1_RVT U501 ( .A1(n22), .A2(n490), .A3(n357), .Y(n360) );
  NAND2X0_RVT U502 ( .A1(n2), .A2(n358), .Y(n359) );
  XOR2X1_RVT U503 ( .A1(n360), .A2(n359), .Y(addout[33]) );
  NAND2X0_RVT U504 ( .A1(n22), .A2(n361), .Y(n362) );
  XNOR2X1_RVT U505 ( .A1(n490), .A2(n362), .Y(addout[32]) );
  FADDX1_RVT U506 ( .A(addin_sum[31]), .B(addin_cout[30]), .CI(n363), .CO(n490), .S(addout[31]) );
  FADDX1_RVT U507 ( .A(addin_sum[30]), .B(addin_cout[29]), .CI(n364), .CO(n363), .S(addout[30]) );
  FADDX1_RVT U508 ( .A(addin_sum[29]), .B(addin_cout[28]), .CI(n365), .CO(n364), .S(addout[29]) );
  FADDX1_RVT U509 ( .A(addin_sum[28]), .B(addin_cout[27]), .CI(n366), .CO(n365), .S(addout[28]) );
  FADDX1_RVT U510 ( .A(addin_cout[26]), .B(addin_sum[27]), .CI(n367), .CO(n366), .S(addout[27]) );
  FADDX1_RVT U511 ( .A(addin_cout[25]), .B(addin_sum[26]), .CI(n368), .CO(n367), .S(addout[26]) );
  FADDX1_RVT U512 ( .A(addin_sum[25]), .B(addin_cout[24]), .CI(n369), .CO(n368), .S(addout[25]) );
  FADDX1_RVT U513 ( .A(addin_sum[24]), .B(addin_cout[23]), .CI(n370), .CO(n369), .S(addout[24]) );
  FADDX1_RVT U514 ( .A(addin_sum[23]), .B(addin_cout[22]), .CI(n371), .CO(n370), .S(addout[23]) );
  FADDX1_RVT U515 ( .A(addin_sum[22]), .B(addin_cout[21]), .CI(n372), .CO(n371), .S(addout[22]) );
  FADDX1_RVT U516 ( .A(addin_sum[21]), .B(addin_cout[20]), .CI(n373), .CO(n372), .S(addout[21]) );
  INVX1_RVT U517 ( .A(n374), .Y(n400) );
  AOI21X1_RVT U518 ( .A1(n376), .A2(n400), .A3(n375), .Y(n379) );
  NAND2X0_RVT U519 ( .A1(n5), .A2(n377), .Y(n378) );
  XOR2X1_RVT U520 ( .A1(n379), .A2(n378), .Y(addout[20]) );
  AOI21X1_RVT U521 ( .A1(n383), .A2(n400), .A3(n382), .Y(n388) );
  NAND2X0_RVT U522 ( .A1(n386), .A2(n385), .Y(n387) );
  XOR2X1_RVT U523 ( .A1(n388), .A2(n387), .Y(addout[19]) );
  AOI21X1_RVT U524 ( .A1(n390), .A2(n400), .A3(n389), .Y(n393) );
  NAND2X0_RVT U525 ( .A1(n6), .A2(n391), .Y(n392) );
  XOR2X1_RVT U526 ( .A1(n393), .A2(n392), .Y(addout[18]) );
  NAND2X0_RVT U527 ( .A1(addin_sum[16]), .A2(n400), .Y(n399) );
  NAND2X0_RVT U528 ( .A1(n397), .A2(n396), .Y(n398) );
  XOR2X1_RVT U529 ( .A1(n399), .A2(n398), .Y(addout[17]) );
  XNOR2X1_RVT U530 ( .A1(n400), .A2(n394), .Y(addout[16]) );
  INVX1_RVT U531 ( .A(n401), .Y(n416) );
  INVX1_RVT U532 ( .A(n403), .Y(n455) );
  OAI21X1_RVT U533 ( .A1(n405), .A2(n455), .A3(n404), .Y(n421) );
  INVX1_RVT U534 ( .A(n421), .Y(n430) );
  INVX1_RVT U535 ( .A(n406), .Y(n407) );
  OAI21X1_RVT U536 ( .A1(n408), .A2(n430), .A3(n407), .Y(n418) );
  AOI21X1_RVT U537 ( .A1(n416), .A2(n418), .A3(n409), .Y(n414) );
  NAND2X0_RVT U538 ( .A1(n412), .A2(n411), .Y(n413) );
  XOR2X1_RVT U539 ( .A1(n414), .A2(n413), .Y(addout[15]) );
  NAND2X0_RVT U540 ( .A1(n416), .A2(n415), .Y(n417) );
  XNOR2X1_RVT U541 ( .A1(n418), .A2(n417), .Y(addout[14]) );
  INVX1_RVT U542 ( .A(n419), .Y(n428) );
  AOI21X1_RVT U543 ( .A1(n428), .A2(n421), .A3(n420), .Y(n426) );
  NAND2X0_RVT U544 ( .A1(n424), .A2(n423), .Y(n425) );
  XOR2X1_RVT U545 ( .A1(n426), .A2(n425), .Y(addout[13]) );
  NAND2X0_RVT U546 ( .A1(n428), .A2(n427), .Y(n429) );
  XOR2X1_RVT U547 ( .A1(n430), .A2(n429), .Y(addout[12]) );
  INVX1_RVT U548 ( .A(n431), .Y(n443) );
  OAI21X1_RVT U549 ( .A1(n435), .A2(n455), .A3(n434), .Y(n445) );
  AOI21X1_RVT U550 ( .A1(n443), .A2(n445), .A3(n436), .Y(n441) );
  NAND2X0_RVT U551 ( .A1(n439), .A2(n438), .Y(n440) );
  XOR2X1_RVT U552 ( .A1(n441), .A2(n440), .Y(addout[11]) );
  NAND2X0_RVT U553 ( .A1(n443), .A2(n442), .Y(n444) );
  XNOR2X1_RVT U554 ( .A1(n445), .A2(n444), .Y(addout[10]) );
  OAI21X1_RVT U555 ( .A1(n451), .A2(n455), .A3(n452), .Y(n450) );
  NAND2X0_RVT U556 ( .A1(n448), .A2(n447), .Y(n449) );
  XNOR2X1_RVT U557 ( .A1(n450), .A2(n449), .Y(addout[9]) );
  NAND2X0_RVT U558 ( .A1(n453), .A2(n452), .Y(n454) );
  XOR2X1_RVT U559 ( .A1(n455), .A2(n454), .Y(addout[8]) );
  INVX1_RVT U560 ( .A(n456), .Y(n479) );
  AOI21X1_RVT U561 ( .A1(n458), .A2(n479), .A3(n457), .Y(n468) );
  OAI21X1_RVT U562 ( .A1(n464), .A2(n468), .A3(n465), .Y(n463) );
  NAND2X0_RVT U563 ( .A1(n461), .A2(n460), .Y(n462) );
  XNOR2X1_RVT U564 ( .A1(n463), .A2(n462), .Y(addout[7]) );
  NAND2X0_RVT U565 ( .A1(n466), .A2(n465), .Y(n467) );
  XOR2X1_RVT U566 ( .A1(n468), .A2(n467), .Y(addout[6]) );
  INVX1_RVT U567 ( .A(n469), .Y(n477) );
  AOI21X1_RVT U568 ( .A1(n477), .A2(n479), .A3(n470), .Y(n475) );
  NAND2X0_RVT U569 ( .A1(n473), .A2(n472), .Y(n474) );
  XOR2X1_RVT U570 ( .A1(n475), .A2(n474), .Y(addout[5]) );
  NAND2X0_RVT U571 ( .A1(n477), .A2(n476), .Y(n478) );
  XNOR2X1_RVT U572 ( .A1(n479), .A2(n478), .Y(addout[4]) );
  AND2X1_RVT U573 ( .A1(n480), .A2(addin_sum[2]), .Y(n485) );
  NAND2X0_RVT U574 ( .A1(n483), .A2(n482), .Y(n484) );
  XNOR2X1_RVT U575 ( .A1(n485), .A2(n484), .Y(addout[3]) );
  XOR2X1_RVT U576 ( .A1(n487), .A2(n486), .Y(addout[2]) );
  XOR2X1_RVT U577 ( .A1(n488), .A2(n489), .Y(addout[1]) );
  INVX1_RVT U578 ( .A(se), .Y(n516) );
  AND2X1_RVT U580 ( .A1(cyc3), .A2(cyc2), .Y(psum_in[98]) );
  AND2X1_RVT U581 ( .A1(cyc2), .A2(psum[97]), .Y(psum_in[97]) );
  AND2X1_RVT U582 ( .A1(cyc2), .A2(psum[96]), .Y(psum_in[96]) );
  AND2X1_RVT U583 ( .A1(cyc2), .A2(psum[95]), .Y(psum_in[95]) );
  AND2X1_RVT U584 ( .A1(cyc2), .A2(psum[94]), .Y(psum_in[94]) );
  AND2X1_RVT U585 ( .A1(cyc2), .A2(psum[93]), .Y(psum_in[93]) );
  AND2X1_RVT U586 ( .A1(cyc2), .A2(psum[92]), .Y(psum_in[92]) );
  AND2X1_RVT U587 ( .A1(cyc2), .A2(psum[91]), .Y(psum_in[91]) );
  AND2X1_RVT U588 ( .A1(cyc2), .A2(psum[90]), .Y(psum_in[90]) );
  AND2X1_RVT U589 ( .A1(cyc2), .A2(psum[89]), .Y(psum_in[89]) );
  AND2X1_RVT U590 ( .A1(cyc2), .A2(psum[88]), .Y(psum_in[88]) );
  AND2X1_RVT U591 ( .A1(cyc2), .A2(psum[87]), .Y(psum_in[87]) );
  AND2X1_RVT U592 ( .A1(cyc2), .A2(psum[86]), .Y(psum_in[86]) );
  AND2X1_RVT U593 ( .A1(cyc2), .A2(psum[85]), .Y(psum_in[85]) );
  AND2X1_RVT U594 ( .A1(cyc2), .A2(psum[84]), .Y(psum_in[84]) );
  AND2X1_RVT U595 ( .A1(cyc2), .A2(psum[83]), .Y(psum_in[83]) );
  AND2X1_RVT U596 ( .A1(cyc2), .A2(psum[82]), .Y(psum_in[82]) );
  AND2X1_RVT U597 ( .A1(cyc2), .A2(psum[81]), .Y(psum_in[81]) );
  AND2X1_RVT U598 ( .A1(cyc2), .A2(psum[80]), .Y(psum_in[80]) );
  AND2X1_RVT U599 ( .A1(cyc2), .A2(psum[79]), .Y(psum_in[79]) );
  AND2X1_RVT U600 ( .A1(cyc2), .A2(psum[78]), .Y(psum_in[78]) );
  AND2X1_RVT U601 ( .A1(cyc2), .A2(psum[77]), .Y(psum_in[77]) );
  AND2X1_RVT U602 ( .A1(cyc2), .A2(psum[76]), .Y(psum_in[76]) );
  AND2X1_RVT U603 ( .A1(cyc2), .A2(psum[75]), .Y(psum_in[75]) );
  AND2X1_RVT U604 ( .A1(cyc2), .A2(psum[74]), .Y(psum_in[74]) );
  AND2X1_RVT U605 ( .A1(cyc2), .A2(psum[73]), .Y(psum_in[73]) );
  AND2X1_RVT U606 ( .A1(cyc2), .A2(psum[72]), .Y(psum_in[72]) );
  AND2X1_RVT U607 ( .A1(cyc2), .A2(psum[71]), .Y(psum_in[71]) );
  AND2X1_RVT U608 ( .A1(cyc2), .A2(psum[70]), .Y(psum_in[70]) );
  AND2X1_RVT U609 ( .A1(cyc2), .A2(psum[69]), .Y(psum_in[69]) );
  AND2X1_RVT U610 ( .A1(cyc2), .A2(psum[68]), .Y(psum_in[68]) );
  AND2X1_RVT U611 ( .A1(cyc2), .A2(psum[67]), .Y(psum_in[67]) );
  AND2X1_RVT U612 ( .A1(cyc2), .A2(psum[66]), .Y(psum_in[66]) );
  AND2X1_RVT U613 ( .A1(cyc2), .A2(psum[65]), .Y(psum_in[65]) );
  AND2X1_RVT U614 ( .A1(cyc2), .A2(psum[64]), .Y(psum_in[64]) );
  AND2X1_RVT U615 ( .A1(cyc2), .A2(psum[63]), .Y(psum_in[63]) );
  AND2X1_RVT U616 ( .A1(cyc2), .A2(psum[62]), .Y(psum_in[62]) );
  AND2X1_RVT U617 ( .A1(cyc2), .A2(psum[61]), .Y(psum_in[61]) );
  AND2X1_RVT U618 ( .A1(cyc2), .A2(psum[60]), .Y(psum_in[60]) );
  AND2X1_RVT U619 ( .A1(cyc2), .A2(psum[59]), .Y(psum_in[59]) );
  AND2X1_RVT U620 ( .A1(cyc2), .A2(psum[58]), .Y(psum_in[58]) );
  AND2X1_RVT U621 ( .A1(cyc2), .A2(psum[57]), .Y(psum_in[57]) );
  AND2X1_RVT U622 ( .A1(cyc2), .A2(psum[56]), .Y(psum_in[56]) );
  AND2X1_RVT U623 ( .A1(cyc2), .A2(psum[55]), .Y(psum_in[55]) );
  AND2X1_RVT U624 ( .A1(cyc2), .A2(psum[54]), .Y(psum_in[54]) );
  AND2X1_RVT U625 ( .A1(cyc2), .A2(psum[53]), .Y(psum_in[53]) );
  AND2X1_RVT U626 ( .A1(cyc2), .A2(psum[52]), .Y(psum_in[52]) );
  AND2X1_RVT U627 ( .A1(cyc2), .A2(psum[51]), .Y(psum_in[51]) );
  AND2X1_RVT U628 ( .A1(cyc2), .A2(psum[50]), .Y(psum_in[50]) );
  AND2X1_RVT U629 ( .A1(cyc2), .A2(psum[49]), .Y(psum_in[49]) );
  AND2X1_RVT U630 ( .A1(cyc2), .A2(psum[48]), .Y(psum_in[48]) );
  AND2X1_RVT U631 ( .A1(cyc2), .A2(psum[47]), .Y(psum_in[47]) );
  AND2X1_RVT U632 ( .A1(cyc2), .A2(psum[46]), .Y(psum_in[46]) );
  AND2X1_RVT U633 ( .A1(cyc2), .A2(psum[45]), .Y(psum_in[45]) );
  AND2X1_RVT U634 ( .A1(cyc2), .A2(psum[44]), .Y(psum_in[44]) );
  AND2X1_RVT U635 ( .A1(cyc2), .A2(psum[43]), .Y(psum_in[43]) );
  AND2X1_RVT U636 ( .A1(cyc2), .A2(psum[42]), .Y(psum_in[42]) );
  AND2X1_RVT U637 ( .A1(cyc2), .A2(psum[41]), .Y(psum_in[41]) );
  AND2X1_RVT U638 ( .A1(cyc2), .A2(psum[40]), .Y(psum_in[40]) );
  AND2X1_RVT U639 ( .A1(cyc2), .A2(psum[39]), .Y(psum_in[39]) );
  AND2X1_RVT U640 ( .A1(cyc2), .A2(psum[38]), .Y(psum_in[38]) );
  AND2X1_RVT U641 ( .A1(cyc2), .A2(psum[37]), .Y(psum_in[37]) );
  AND2X1_RVT U642 ( .A1(cyc2), .A2(psum[36]), .Y(psum_in[36]) );
  AND2X1_RVT U643 ( .A1(cyc2), .A2(psum[35]), .Y(psum_in[35]) );
  AND2X1_RVT U644 ( .A1(cyc2), .A2(psum[34]), .Y(psum_in[34]) );
  AND2X1_RVT U645 ( .A1(cyc2), .A2(psum[33]), .Y(psum_in[33]) );
  AND2X1_RVT U646 ( .A1(cyc2), .A2(psum[32]), .Y(psum_in[32]) );
  AND2X1_RVT U647 ( .A1(cyc2), .A2(pcout[97]), .Y(pcout_in[97]) );
  AND2X1_RVT U648 ( .A1(cyc2), .A2(pcout[96]), .Y(pcout_in[96]) );
  AND2X1_RVT U649 ( .A1(cyc2), .A2(pcout[95]), .Y(pcout_in[95]) );
  AND2X1_RVT U650 ( .A1(cyc2), .A2(pcout[94]), .Y(pcout_in[94]) );
  AND2X1_RVT U651 ( .A1(cyc2), .A2(pcout[93]), .Y(pcout_in[93]) );
  AND2X1_RVT U652 ( .A1(cyc2), .A2(pcout[92]), .Y(pcout_in[92]) );
  AND2X1_RVT U653 ( .A1(cyc2), .A2(pcout[91]), .Y(pcout_in[91]) );
  AND2X1_RVT U654 ( .A1(cyc2), .A2(pcout[90]), .Y(pcout_in[90]) );
  AND2X1_RVT U655 ( .A1(cyc2), .A2(pcout[89]), .Y(pcout_in[89]) );
  AND2X1_RVT U656 ( .A1(cyc2), .A2(pcout[88]), .Y(pcout_in[88]) );
  AND2X1_RVT U657 ( .A1(cyc2), .A2(pcout[87]), .Y(pcout_in[87]) );
  AND2X1_RVT U658 ( .A1(cyc2), .A2(pcout[86]), .Y(pcout_in[86]) );
  AND2X1_RVT U659 ( .A1(cyc2), .A2(pcout[85]), .Y(pcout_in[85]) );
  AND2X1_RVT U660 ( .A1(cyc2), .A2(pcout[84]), .Y(pcout_in[84]) );
  AND2X1_RVT U661 ( .A1(cyc2), .A2(pcout[83]), .Y(pcout_in[83]) );
  AND2X1_RVT U662 ( .A1(cyc2), .A2(pcout[82]), .Y(pcout_in[82]) );
  AND2X1_RVT U663 ( .A1(cyc2), .A2(pcout[81]), .Y(pcout_in[81]) );
  AND2X1_RVT U664 ( .A1(cyc2), .A2(pcout[80]), .Y(pcout_in[80]) );
  AND2X1_RVT U665 ( .A1(cyc2), .A2(pcout[79]), .Y(pcout_in[79]) );
  AND2X1_RVT U666 ( .A1(cyc2), .A2(pcout[78]), .Y(pcout_in[78]) );
  AND2X1_RVT U667 ( .A1(cyc2), .A2(pcout[77]), .Y(pcout_in[77]) );
  AND2X1_RVT U668 ( .A1(cyc2), .A2(pcout[76]), .Y(pcout_in[76]) );
  AND2X1_RVT U669 ( .A1(cyc2), .A2(pcout[75]), .Y(pcout_in[75]) );
  AND2X1_RVT U670 ( .A1(cyc2), .A2(pcout[74]), .Y(pcout_in[74]) );
  AND2X1_RVT U671 ( .A1(cyc2), .A2(pcout[73]), .Y(pcout_in[73]) );
  AND2X1_RVT U672 ( .A1(cyc2), .A2(pcout[72]), .Y(pcout_in[72]) );
  AND2X1_RVT U673 ( .A1(cyc2), .A2(pcout[71]), .Y(pcout_in[71]) );
  AND2X1_RVT U674 ( .A1(cyc2), .A2(pcout[70]), .Y(pcout_in[70]) );
  AND2X1_RVT U675 ( .A1(cyc2), .A2(pcout[69]), .Y(pcout_in[69]) );
  AND2X1_RVT U676 ( .A1(cyc2), .A2(pcout[68]), .Y(pcout_in[68]) );
  AND2X1_RVT U677 ( .A1(cyc2), .A2(pcout[67]), .Y(pcout_in[67]) );
  AND2X1_RVT U678 ( .A1(cyc2), .A2(pcout[66]), .Y(pcout_in[66]) );
  AND2X1_RVT U679 ( .A1(cyc2), .A2(pcout[65]), .Y(pcout_in[65]) );
  AND2X1_RVT U680 ( .A1(cyc2), .A2(pcout[64]), .Y(pcout_in[64]) );
  AND2X1_RVT U681 ( .A1(cyc2), .A2(pcout[63]), .Y(pcout_in[63]) );
  AND2X1_RVT U682 ( .A1(cyc2), .A2(pcout[62]), .Y(pcout_in[62]) );
  AND2X1_RVT U683 ( .A1(cyc2), .A2(pcout[61]), .Y(pcout_in[61]) );
  AND2X1_RVT U684 ( .A1(cyc2), .A2(pcout[60]), .Y(pcout_in[60]) );
  AND2X1_RVT U685 ( .A1(cyc2), .A2(pcout[59]), .Y(pcout_in[59]) );
  AND2X1_RVT U686 ( .A1(cyc2), .A2(pcout[58]), .Y(pcout_in[58]) );
  AND2X1_RVT U687 ( .A1(cyc2), .A2(pcout[57]), .Y(pcout_in[57]) );
  AND2X1_RVT U688 ( .A1(cyc2), .A2(pcout[56]), .Y(pcout_in[56]) );
  AND2X1_RVT U689 ( .A1(cyc2), .A2(pcout[55]), .Y(pcout_in[55]) );
  AND2X1_RVT U690 ( .A1(cyc2), .A2(pcout[54]), .Y(pcout_in[54]) );
  AND2X1_RVT U691 ( .A1(cyc2), .A2(pcout[53]), .Y(pcout_in[53]) );
  AND2X1_RVT U692 ( .A1(cyc2), .A2(pcout[52]), .Y(pcout_in[52]) );
  AND2X1_RVT U693 ( .A1(cyc2), .A2(pcout[51]), .Y(pcout_in[51]) );
  AND2X1_RVT U694 ( .A1(cyc2), .A2(pcout[50]), .Y(pcout_in[50]) );
  AND2X1_RVT U695 ( .A1(cyc2), .A2(pcout[49]), .Y(pcout_in[49]) );
  AND2X1_RVT U696 ( .A1(cyc2), .A2(pcout[48]), .Y(pcout_in[48]) );
  AND2X1_RVT U697 ( .A1(cyc2), .A2(pcout[47]), .Y(pcout_in[47]) );
  AND2X1_RVT U698 ( .A1(cyc2), .A2(pcout[46]), .Y(pcout_in[46]) );
  AND2X1_RVT U699 ( .A1(cyc2), .A2(pcout[45]), .Y(pcout_in[45]) );
  AND2X1_RVT U700 ( .A1(cyc2), .A2(pcout[44]), .Y(pcout_in[44]) );
  AND2X1_RVT U701 ( .A1(cyc2), .A2(pcout[43]), .Y(pcout_in[43]) );
  AND2X1_RVT U702 ( .A1(cyc2), .A2(pcout[42]), .Y(pcout_in[42]) );
  AND2X1_RVT U703 ( .A1(cyc2), .A2(pcout[41]), .Y(pcout_in[41]) );
  AND2X1_RVT U704 ( .A1(cyc2), .A2(pcout[40]), .Y(pcout_in[40]) );
  AND2X1_RVT U705 ( .A1(cyc2), .A2(pcout[39]), .Y(pcout_in[39]) );
  AND2X1_RVT U706 ( .A1(cyc2), .A2(pcout[38]), .Y(pcout_in[38]) );
  AND2X1_RVT U707 ( .A1(cyc2), .A2(pcout[37]), .Y(pcout_in[37]) );
  AND2X1_RVT U708 ( .A1(cyc2), .A2(pcout[36]), .Y(pcout_in[36]) );
  AND2X1_RVT U709 ( .A1(cyc2), .A2(pcout[35]), .Y(pcout_in[35]) );
  AND2X1_RVT U710 ( .A1(cyc2), .A2(pcout[34]), .Y(pcout_in[34]) );
  AND2X1_RVT U711 ( .A1(cyc2), .A2(pcout[33]), .Y(pcout_in[33]) );
  AND2X1_RVT U712 ( .A1(cyc2), .A2(pcout[32]), .Y(pcout_in[32]) );
  AND2X1_RVT U713 ( .A1(cyc2), .A2(pcout[31]), .Y(pcout_in[31]) );
  AND2X1_RVT U714 ( .A1(cyc3), .A2(n490), .Y(add_cin) );
  NAND2X0_RVT U715 ( .A1(mul_step), .A2(valid), .Y(n76) );
endmodule


module fpu_mul ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_mul, 
        fmul_clken_l, fmul_clken_l_buf1, arst_l, grst_l, rclk, mul_pipe_active, 
        m1stg_step, m6stg_fmul_in, m6stg_id_in, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, se_mul, se_mul64, si, so, mul_dest_rdy_BAR, 
        mul_dest_rdya_BAR );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] m6stg_id_in;
  output [4:0] mul_exc_out;
  output [10:0] mul_exp_out;
  output [51:0] mul_frac_out;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_mul, fmul_clken_l, fmul_clken_l_buf1, arst_l,
         grst_l, rclk, se_mul, se_mul64, si, mul_dest_rdy_BAR,
         mul_dest_rdya_BAR;
  output mul_pipe_active, m1stg_step, m6stg_fmul_in, m6stg_fmul_dbl_dst,
         m6stg_fmuls, mul_sign_out, so;
  wire   mul_dest_rdya, m5stg_fracadd_cout, m5stg_frac_neq_0,
         m5stg_frac_dbl_nx, m5stg_frac_sng_nx, m3stg_expadd_eq_0,
         m3stg_expadd_lte_0_inv, m4stg_frac_105, mul_rst_l, m1stg_snan_sng_in1,
         m1stg_snan_dbl_in1, m1stg_snan_sng_in2, m1stg_snan_dbl_in2,
         m1stg_sngop, m1stg_dblop, m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld,
         m2stg_fmuls, m2stg_fmuld, m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld,
         m5stg_fmulda, m6stg_step, m5stg_in_of, m2stg_frac1_dbl_norm,
         m2stg_frac1_dbl_dnrm, m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm,
         m2stg_frac1_inf, m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm,
         m2stg_frac2_sng_norm, m2stg_frac2_sng_dnrm, m2stg_frac2_inf,
         m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, m2stg_exp_expadd,
         m2stg_exp_0bff, m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero,
         m4stg_inc_exp_54, m4stg_inc_exp_55, m4stg_inc_exp_105,
         m4stg_left_shift_step, m4stg_right_shift_step, m5stg_to_0,
         m5stg_to_0_inv, mul_frac_out_fracadd, mul_frac_out_frac,
         mul_exp_out_exp_plus1, mul_exp_out_exp, m4stg_shl_54, m4stg_shl_55,
         net211155, net211156, net211157, net211158, net211159, net211160;
  wire   [12:0] m5stg_exp;
  wire   [5:0] m1stg_ld0_1;
  wire   [5:0] m1stg_ld0_2;
  wire   [12:0] m3stg_exp;
  wire   [6:0] m3stg_ld0_inv;
  wire   [12:0] m4stg_exp;
  wire   [32:0] m5stg_frac_32_0;
  wire   [6:0] m3bstg_ld0_inv;
  wire   [5:0] m4stg_sh_cnt_in;
  wire   [105:0] m4stg_frac;
  wire   [52:0] m2stg_frac1_array_in;
  wire   [52:0] m2stg_frac2_array_in;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;
  assign mul_dest_rdya = mul_dest_rdya_BAR;

  fpu_mul_ctl fpu_mul_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_51(inq_in2[51]), .inq_in2_54(
        inq_in2[54]), .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(inq_op), .inq_mul(
        inq_mul), .inq_rnd_mode(inq_rnd_mode), .inq_id(inq_id), .inq_in1_63(
        inq_in1[63]), .inq_in2_63(inq_in2[63]), .mul_dest_rdy(net211158), 
        .m5stg_exp(m5stg_exp), .m5stg_fracadd_cout(m5stg_fracadd_cout), 
        .m5stg_frac_neq_0(m5stg_frac_neq_0), .m5stg_frac_dbl_nx(
        m5stg_frac_dbl_nx), .m5stg_frac_sng_nx(m5stg_frac_sng_nx), 
        .m1stg_ld0_1(m1stg_ld0_1), .m1stg_ld0_2(m1stg_ld0_2), .m3stg_exp(
        m3stg_exp), .m3stg_expadd_eq_0(m3stg_expadd_eq_0), 
        .m3stg_expadd_lte_0_inv(m3stg_expadd_lte_0_inv), .m3stg_ld0_inv(
        m3stg_ld0_inv[5:0]), .m4stg_exp({net211159, m4stg_exp[11:0]}), 
        .m4stg_frac_105(m4stg_frac_105), .m5stg_frac(m5stg_frac_32_0), 
        .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), .mul_pipe_active(
        mul_pipe_active), .m1stg_snan_sng_in1(m1stg_snan_sng_in1), 
        .m1stg_snan_dbl_in1(m1stg_snan_dbl_in1), .m1stg_snan_sng_in2(
        m1stg_snan_sng_in2), .m1stg_snan_dbl_in2(m1stg_snan_dbl_in2), 
        .m1stg_step(m1stg_step), .m1stg_sngop(m1stg_sngop), .m1stg_dblop(
        m1stg_dblop), .m1stg_dblop_inv(m1stg_dblop_inv), .m1stg_fmul(
        m1stg_fmul), .m1stg_fsmuld(m1stg_fsmuld), .m2stg_fmuls(m2stg_fmuls), 
        .m2stg_fmuld(m2stg_fmuld), .m2stg_fsmuld(m2stg_fsmuld), .m5stg_fmuls(
        m5stg_fmuls), .m5stg_fmuld(m5stg_fmuld), .m5stg_fmulda(m5stg_fmulda), 
        .m6stg_fmul_in(m6stg_fmul_in), .m6stg_id_in(m6stg_id_in), 
        .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), .m6stg_fmuls(m6stg_fmuls), 
        .m6stg_step(m6stg_step), .mul_sign_out(mul_sign_out), .m5stg_in_of(
        m5stg_in_of), .mul_exc_out({mul_exc_out[4:2], SYNOPSYS_UNCONNECTED__0, 
        mul_exc_out[0]}), .m2stg_frac1_dbl_norm(m2stg_frac1_dbl_norm), 
        .m2stg_frac1_dbl_dnrm(m2stg_frac1_dbl_dnrm), .m2stg_frac1_sng_norm(
        m2stg_frac1_sng_norm), .m2stg_frac1_sng_dnrm(m2stg_frac1_sng_dnrm), 
        .m2stg_frac1_inf(m2stg_frac1_inf), .m2stg_frac2_dbl_norm(
        m2stg_frac2_dbl_norm), .m2stg_frac2_dbl_dnrm(m2stg_frac2_dbl_dnrm), 
        .m2stg_frac2_sng_norm(m2stg_frac2_sng_norm), .m2stg_frac2_sng_dnrm(
        m2stg_frac2_sng_dnrm), .m2stg_frac2_inf(m2stg_frac2_inf), 
        .m1stg_inf_zero_in(m1stg_inf_zero_in), .m1stg_inf_zero_in_dbl(
        m1stg_inf_zero_in_dbl), .m2stg_exp_expadd(m2stg_exp_expadd), 
        .m2stg_exp_0bff(m2stg_exp_0bff), .m2stg_exp_017f(m2stg_exp_017f), 
        .m2stg_exp_04ff(m2stg_exp_04ff), .m2stg_exp_zero(m2stg_exp_zero), 
        .m3bstg_ld0_inv(m3bstg_ld0_inv), .m4stg_sh_cnt_in(m4stg_sh_cnt_in), 
        .m4stg_inc_exp_54(m4stg_inc_exp_54), .m4stg_inc_exp_55(
        m4stg_inc_exp_55), .m4stg_inc_exp_105(m4stg_inc_exp_105), 
        .m4stg_left_shift_step(m4stg_left_shift_step), 
        .m4stg_right_shift_step(m4stg_right_shift_step), .m5stg_to_0(
        m5stg_to_0), .m5stg_to_0_inv(m5stg_to_0_inv), .mul_frac_out_fracadd(
        mul_frac_out_fracadd), .mul_frac_out_frac(mul_frac_out_frac), 
        .mul_exp_out_exp_plus1(mul_exp_out_exp_plus1), .mul_exp_out_exp(
        mul_exp_out_exp), .mula_rst_l(mul_rst_l), .se(se_mul), .si(net211160), 
        .mul_dest_rdya_BAR(mul_dest_rdya) );
  fpu_mul_exp_dp fpu_mul_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .m6stg_step(m6stg_step), .m1stg_dblop(m1stg_dblop), 
        .m1stg_sngop(m1stg_sngop), .m2stg_exp_expadd(m2stg_exp_expadd), 
        .m2stg_exp_0bff(m2stg_exp_0bff), .m2stg_exp_017f(m2stg_exp_017f), 
        .m2stg_exp_04ff(m2stg_exp_04ff), .m2stg_exp_zero(m2stg_exp_zero), 
        .m1stg_fsmuld(m1stg_fsmuld), .m2stg_fmuld(m2stg_fmuld), .m2stg_fmuls(
        m2stg_fmuls), .m2stg_fsmuld(m2stg_fsmuld), .m3stg_ld0_inv(
        m3stg_ld0_inv), .m5stg_fracadd_cout(m5stg_fracadd_cout), 
        .mul_exp_out_exp_plus1(mul_exp_out_exp_plus1), .mul_exp_out_exp(
        mul_exp_out_exp), .m5stg_in_of(m5stg_in_of), .m5stg_fmuld(m5stg_fmuld), 
        .m5stg_to_0_inv(m5stg_to_0_inv), .m4stg_shl_54(m4stg_shl_54), 
        .m4stg_shl_55(m4stg_shl_55), .m4stg_inc_exp_54(m4stg_inc_exp_54), 
        .m4stg_inc_exp_55(m4stg_inc_exp_55), .m4stg_inc_exp_105(
        m4stg_inc_exp_105), .fmul_clken_l(fmul_clken_l_buf1), .rclk(rclk), 
        .m3stg_exp(m3stg_exp), .m3stg_expadd_eq_0(m3stg_expadd_eq_0), 
        .m3stg_expadd_lte_0_inv(m3stg_expadd_lte_0_inv), .m4stg_exp({
        SYNOPSYS_UNCONNECTED__1, m4stg_exp[11:0]}), .m5stg_exp(m5stg_exp), 
        .mul_exp_out(mul_exp_out), .se(se_mul), .si(net211157) );
  fpu_mul_frac_dp fpu_mul_frac_dp ( .inq_in1(inq_in1[54:0]), .inq_in2(
        inq_in2[54:0]), .m6stg_step(m6stg_step), .m2stg_frac1_dbl_norm(
        m2stg_frac1_dbl_norm), .m2stg_frac1_dbl_dnrm(m2stg_frac1_dbl_dnrm), 
        .m2stg_frac1_sng_norm(m2stg_frac1_sng_norm), .m2stg_frac1_sng_dnrm(
        m2stg_frac1_sng_dnrm), .m2stg_frac1_inf(m2stg_frac1_inf), 
        .m1stg_snan_dbl_in1(m1stg_snan_dbl_in1), .m1stg_snan_sng_in1(
        m1stg_snan_sng_in1), .m2stg_frac2_dbl_norm(m2stg_frac2_dbl_norm), 
        .m2stg_frac2_dbl_dnrm(m2stg_frac2_dbl_dnrm), .m2stg_frac2_sng_norm(
        m2stg_frac2_sng_norm), .m2stg_frac2_sng_dnrm(m2stg_frac2_sng_dnrm), 
        .m2stg_frac2_inf(m2stg_frac2_inf), .m1stg_snan_dbl_in2(
        m1stg_snan_dbl_in2), .m1stg_snan_sng_in2(m1stg_snan_sng_in2), 
        .m1stg_inf_zero_in(m1stg_inf_zero_in), .m1stg_inf_zero_in_dbl(
        m1stg_inf_zero_in_dbl), .m1stg_dblop(m1stg_dblop), .m1stg_dblop_inv(
        m1stg_dblop_inv), .m4stg_frac(m4stg_frac), .m4stg_sh_cnt_in(
        m4stg_sh_cnt_in), .m3bstg_ld0_inv(m3bstg_ld0_inv), 
        .m4stg_left_shift_step(m4stg_left_shift_step), 
        .m4stg_right_shift_step(m4stg_right_shift_step), .m5stg_fmuls(
        m5stg_fmuls), .m5stg_fmulda(m5stg_fmulda), .mul_frac_out_fracadd(
        mul_frac_out_fracadd), .mul_frac_out_frac(mul_frac_out_frac), 
        .m5stg_in_of(m5stg_in_of), .m5stg_to_0(m5stg_to_0), .fmul_clken_l(
        fmul_clken_l), .rclk(rclk), .m2stg_frac1_array_in(m2stg_frac1_array_in), .m2stg_frac2_array_in(m2stg_frac2_array_in), .m1stg_ld0_1(m1stg_ld0_1), 
        .m1stg_ld0_2(m1stg_ld0_2), .m4stg_frac_105(m4stg_frac_105), 
        .m3stg_ld0_inv(m3stg_ld0_inv), .m4stg_shl_54(m4stg_shl_54), 
        .m4stg_shl_55(m4stg_shl_55), .m5stg_frac_32_0(m5stg_frac_32_0), 
        .m5stg_frac_dbl_nx(m5stg_frac_dbl_nx), .m5stg_frac_sng_nx(
        m5stg_frac_sng_nx), .m5stg_frac_neq_0(m5stg_frac_neq_0), 
        .m5stg_fracadd_cout(m5stg_fracadd_cout), .mul_frac_out(mul_frac_out), 
        .se(se_mul), .si(net211156) );
  mul64 i_m4stg_frac ( .rs1_l({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, m2stg_frac1_array_in}), .rs2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m2stg_frac2_array_in}), 
        .valid(m1stg_fmul), .areg({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .accreg({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .x2(1'b0), .out({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, m4stg_frac}), .rclk(rclk), .si(net211155), 
        .se(se_mul64), .mul_rst_l(mul_rst_l), .mul_step(m6stg_step) );
endmodule


module dffrl_async_SIZE1_2 ( din, clk, rst_l, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  wire   N4, n1;

  DFFARX1_RVT \q_reg[0]  ( .D(N4), .CLK(clk), .RSTB(rst_l), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
endmodule


module dffe_SIZE1_30 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_29 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_28 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_27 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_26 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_25 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_24 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_23 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_22 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_21 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_20 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_19 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_18 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_17 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dff_SIZE1_28 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_27 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_26 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_25 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_24 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_23 ( din, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0]_BAR ;


  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\q[0]_BAR ) );
endmodule


module dff_SIZE1_22 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_21 ( din, clk, se, si, so, \q[0]  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0] ;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(\q[0] ) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_20 ( din, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0]_BAR ;


  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\q[0]_BAR ) );
endmodule


module dff_SIZE1_19 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_18 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_16 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_13 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_11 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_10 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_9 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dffr_SIZE8 ( din, clk, rst, se, si, so, \q[7] , \q[6] , \q[5]_BAR , 
        \q[4] , \q[3] , \q[2] , \q[1] , \q[0]  );
  input [7:0] din;
  input [7:0] si;
  output [7:0] so;
  input clk, rst, se;
  output \q[7] , \q[6] , \q[5]_BAR , \q[4] , \q[3] , \q[2] , \q[1] , \q[0] ;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, n1;
  wire   [7:0] q;

  DFFX1_RVT \q_reg[7]  ( .D(N21), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N20), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N19), .CLK(clk), .QN(\q[5]_BAR ) );
  DFFX1_RVT \q_reg[4]  ( .D(N18), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N17), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N16), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N15), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N14), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N14) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N15) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N16) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[3]), .Y(N17) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[4]), .Y(N18) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[5]), .Y(N19) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[6]), .Y(N20) );
  AND2X1_RVT U11 ( .A1(n1), .A2(din[7]), .Y(N21) );
endmodule


module dffr_SIZE1_3 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_3 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_3 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE1_16 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_2 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_2 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N4), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N4), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N4), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  OR2X1_RVT U5 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffr_SIZE3_0 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N9, N10, N11, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N11) );
endmodule


module dffr_SIZE1_2 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dffr_SIZE3_4 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N9, N10, N11, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N11) );
endmodule


module dffr_SIZE3_3 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N9, N10, N11, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_2 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_2 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffre_SIZE1_7 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dff_SIZE1_8 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dffr_SIZE3_2 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N9, N10, N11, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N11) );
endmodule


module dffr_SIZE3_1 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N9, N10, N11, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n1) );
  AND2X1_RVT U4 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[2]), .Y(N11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE3_1 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N9, N10, N11, net24318, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE3_1 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24318), .TE(1'b0) );
  DFFX1_RVT \q_reg[2]  ( .D(N11), .CLK(net24318), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N10), .CLK(net24318), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N9), .CLK(net24318), .Q(q[0]) );
  INVX1_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N9) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N10) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N11) );
  NAND2X0_RVT U9 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffre_SIZE1_6 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2;

  DFFX1_RVT \q_reg[0]  ( .D(n2), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U2 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U3 ( .A1(rst), .A2(se), .A3(n1), .Y(n2) );
endmodule


module dffe_SIZE2_2 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE5_1 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, net24300, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE5_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24300), .TE(1'b0) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24300), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24300), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24300), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24300), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24300), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  OR2X1_RVT U9 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module dffe_SIZE1_15 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_14 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE2_1 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[1]  ( .D(n4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(q[0]) );
  NOR2X0_RVT U2 ( .A1(se), .A2(en), .Y(n3) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(en), .A2(n1), .Y(n2) );
  AO22X1_RVT U5 ( .A1(n3), .A2(q[1]), .A3(din[1]), .A4(n2), .Y(n4) );
  AO22X1_RVT U6 ( .A1(n3), .A2(q[0]), .A3(n2), .A4(din[0]), .Y(n5) );
endmodule


module dff_SIZE10_1 ( din, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, n1;

  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
endmodule


module dffe_SIZE1_13 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffre_SIZE6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffre_SIZE6_1 ( din, rst, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input rst, en, clk, se;
  wire   N12, N13, N14, N15, N16, N17, net24282, n1, n2, n3, n5;

  SNPS_CLOCK_GATE_HIGH_dffre_SIZE6_1 clk_gate_q_reg ( .CLK(clk), .EN(n5), 
        .ENCLK(net24282), .TE(1'b0) );
  DFFX1_RVT \q_reg[5]  ( .D(N17), .CLK(net24282), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N16), .CLK(net24282), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N15), .CLK(net24282), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N14), .CLK(net24282), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N13), .CLK(net24282), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N12), .CLK(net24282), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(se), .A2(rst), .Y(n3) );
  AND2X1_RVT U4 ( .A1(en), .A2(n3), .Y(n1) );
  AND2X1_RVT U5 ( .A1(n1), .A2(din[0]), .Y(N12) );
  AND2X1_RVT U6 ( .A1(n1), .A2(din[1]), .Y(N13) );
  AND2X1_RVT U7 ( .A1(n1), .A2(din[2]), .Y(N14) );
  AND2X1_RVT U8 ( .A1(n1), .A2(din[3]), .Y(N15) );
  AND2X1_RVT U9 ( .A1(n1), .A2(din[4]), .Y(N16) );
  AND2X1_RVT U10 ( .A1(n1), .A2(din[5]), .Y(N17) );
  NAND2X0_RVT U12 ( .A1(n3), .A2(n2), .Y(n5) );
endmodule


module dffre_SIZE1_5 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffre_SIZE1_4 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffre_SIZE1_3 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffre_SIZE1_2 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  NOR2X0_RVT U3 ( .A1(rst), .A2(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_12 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_11 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_10 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_9 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_8 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_7 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_6 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_5 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_4 ( din, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(\q[0] ), .A3(n2), .A4(din[0]), .A5(n1), .Y(n5)
         );
endmodule


module dffe_SIZE1_3 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dffe_SIZE1_2 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX0_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module dff_SIZE1_7 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dff_SIZE1_6 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N3, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
endmodule


module dffr_SIZE1_1 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N7, n1;

  DFFX1_RVT \q_reg[0]  ( .D(N7), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(din[0]), .Y(n1) );
  NOR3X0_RVT U4 ( .A1(se), .A2(rst), .A3(n1), .Y(N7) );
endmodule


module dffe_SIZE1_1 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   n1, n2, n3;

  DFFX1_RVT \q_reg[0]  ( .D(n3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U2 ( .A(en), .Y(n2) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(en), .A2(q[0]), .A3(n2), .A4(din[0]), .A5(n1), .Y(n3)
         );
endmodule


module fpu_div_ctl ( inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, inq_op, div_exp1, inq_rnd_mode, inq_id, 
        inq_in1_63, inq_in2_63, inq_div, div_exp_out, div_frac_add_52_inva, 
        div_frac_add_in1_neq_0, div_frac_out_54, d6stg_frac_0, d6stg_frac_1, 
        d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, d6stg_frac_31, 
        div_frac_out_53, div_expadd2_12, arst_l, grst_l, rclk, div_pipe_active, 
        d1stg_snan_sng_in1, d1stg_snan_dbl_in1, d1stg_snan_sng_in2, 
        d1stg_snan_dbl_in2, d1stg_step, d1stg_dblop, d234stg_fdiv, d3stg_fdiv, 
        d4stg_fdiv, d5stg_fdiva, d5stg_fdivb, d5stg_fdivs, d5stg_fdivd, 
        d6stg_fdiv, d6stg_fdivs, d6stg_fdivd, d7stg_fdiv, d7stg_fdivd, 
        d8stg_fdiv_in, d8stg_fdivs, d8stg_fdivd, div_id_out_in, div_sign_out, 
        div_exc_out, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm, 
        div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm, 
        div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm, 
        div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf, 
        div_norm_qnan, div_norm_zero, div_frac_add_in2_load, 
        d6stg_frac_out_shl1, d6stg_frac_out_nosh, div_frac_add_in1_add, 
        div_frac_add_in1_load, d7stg_rndup_inv, d7stg_to_0, d7stg_to_0_inv, 
        div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl, 
        div_frac_out_shl1_sng, div_frac_out_of, div_frac_out_load, 
        div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl, 
        div_expadd1_in2_exp_in2_sng, div_exp1_expadd1, div_exp1_0835, 
        div_exp1_0118, div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out, 
        div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd22_inv, 
        div_exp_out_expadd2, div_exp_out_of, div_exp_out_exp_out, 
        div_exp_out_load, se, si, so, div_dest_rdy_BAR );
  input [7:0] inq_op;
  input [12:0] div_exp1;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [12:0] div_exp_out;
  output [9:0] div_id_out_in;
  output [4:0] div_exc_out;
  input inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs,
         inq_in1_63, inq_in2_63, inq_div, div_frac_add_52_inva,
         div_frac_add_in1_neq_0, div_frac_out_54, d6stg_frac_0, d6stg_frac_1,
         d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, d6stg_frac_31,
         div_frac_out_53, div_expadd2_12, arst_l, grst_l, rclk, se, si,
         div_dest_rdy_BAR;
  output div_pipe_active, d1stg_snan_sng_in1, d1stg_snan_dbl_in1,
         d1stg_snan_sng_in2, d1stg_snan_dbl_in2, d1stg_step, d1stg_dblop,
         d234stg_fdiv, d3stg_fdiv, d4stg_fdiv, d5stg_fdiva, d5stg_fdivb,
         d5stg_fdivs, d5stg_fdivd, d6stg_fdiv, d6stg_fdivs, d6stg_fdivd,
         d7stg_fdiv, d7stg_fdivd, d8stg_fdiv_in, d8stg_fdivs, d8stg_fdivd,
         div_sign_out, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm,
         div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm,
         div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm,
         div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf,
         div_norm_qnan, div_norm_zero, div_frac_add_in2_load,
         d6stg_frac_out_shl1, d6stg_frac_out_nosh, div_frac_add_in1_add,
         div_frac_add_in1_load, d7stg_rndup_inv, d7stg_to_0, d7stg_to_0_inv,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, div_frac_out_load,
         div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl,
         div_expadd1_in2_exp_in2_sng, div_exp1_expadd1, div_exp1_0835,
         div_exp1_0118, div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd22_inv,
         div_exp_out_expadd2, div_exp_out_of, div_exp_out_exp_out,
         div_exp_out_load, so;
  wire   div_dest_rdy, div_frac_out_of, div_ctl_rst_l, div_frac_in1_51,
         div_frac_in1_54, div_frac_in1_53_0_neq_0, div_frac_in1_50_0_neq_0,
         div_frac_in1_53_32_neq_0, div_exp_in1_exp_eq_0,
         div_exp_in1_exp_neq_ffs, div_frac_in2_51, div_frac_in2_54,
         div_frac_in2_53_0_neq_0, div_frac_in2_50_0_neq_0,
         div_frac_in2_53_32_neq_0, div_exp_in2_exp_eq_0,
         div_exp_in2_exp_neq_ffs, d1stg_denorm_sng_in2, d1stg_denorm_dbl_in2,
         d2stg_denorm_sng_in2, d2stg_denorm_dbl_in2, d1stg_norm_sng_in2,
         d1stg_norm_dbl_in2, d2stg_norm_sng_in2, d2stg_norm_dbl_in2,
         d1stg_snan_in1, d1stg_snan_in2, d1stg_qnan_in1, d1stg_qnan_in2,
         d1stg_nan_in2, d1stg_nan_in, d2stg_snan_in1, d2stg_snan_in2,
         d2stg_qnan_in1, d2stg_qnan_in2, d2stg_nan_in2, d2stg_nan_in,
         d1stg_inf_in1, d1stg_2inf_in, d2stg_inf_in1, d2stg_2inf_in,
         d1stg_infnan_in, d2stg_infnan_in, d1stg_zero_in2, d1stg_zero_in,
         d1stg_2zero_in, d2stg_zero_in2, d2stg_zero_in, d2stg_2zero_in,
         d1stg_div, divs_cnt_lt_23, divd_cnt_lt_52, divs_cnt_lt_23a,
         divd_cnt_lt_52a, d1stg_div_in, \d1stg_opdec[2] , d234stg_fdiv_in,
         \d2stg_opdec[2] , d5stg_step, \d5stg_opdec[2] , d5stg_fdivb_in,
         \d7stg_opdec[1] , \d8stg_opdec[2] , div_pipe_active_in, d1stg_sign1,
         d1stg_sign2, d1stg_sign, div_bkend_step, div_cnt_step,
         div_cnt_lt_step, divs_cnt_lt_23_in, divd_cnt_lt_52_in, div_of_mask,
         div_nv_out_in, div_dz_out_in, d7stg_in_of, div_of_out_tmp1_in,
         div_of_out_tmp1, div_of_out_tmp2, div_out_52_inv, d7stg_grd,
         d7stg_stk, div_uf_out_in, div_nx_out_in, div_nx_out, d7stg_lsb_in,
         d7stg_grd_in, d7stg_stk_in, d7stg_lsb, div_expadd1_in1_dbl_in,
         div_expadd1_in1_sng_in, div_expadd2_in1_exp_out_in,
         div_expadd2_no_decr_load, n148, n149, n150, n151, n154, n156, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n152, n153, n155, n157, n158, n159, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n183;
  wire   [4:0] d1stg_sngopa;
  wire   [4:0] d1stg_dblopa;
  wire   [7:0] d1stg_op_in;
  wire   [7:0] d1stg_op;
  wire   [1:0] d3stg_opdec;
  wire   [1:0] d4stg_opdec;
  wire   [5:0] div_cnt;
  wire   [2:0] d6stg_opdec_in;
  wire   [1:0] d1stg_rnd_mode;
  wire   [4:0] d1stg_id;
  wire   [1:0] div_rnd_mode;
  wire   [9:0] div_id_out;
  wire   [5:0] div_cnt_in;
  assign div_dest_rdy = div_dest_rdy_BAR;
  assign div_exp_out_of = div_frac_out_of;
  assign so = 1'b0;

  dffrl_async_SIZE1_2 dffrl_div_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(div_ctl_rst_l), .se(se), .si(1'b0) );
  dffe_SIZE1_30 i_div_frac_in1_51 ( .din(inq_in1_51), .en(d1stg_step), .clk(
        rclk), .q(div_frac_in1_51), .se(se), .si(1'b0) );
  dffe_SIZE1_29 i_div_frac_in1_54 ( .din(inq_in1_54), .en(d1stg_step), .clk(
        rclk), .q(div_frac_in1_54), .se(se), .si(1'b0) );
  dffe_SIZE1_28 i_div_frac_in1_53_0_neq_0 ( .din(inq_in1_53_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_53_0_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_27 i_div_frac_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_50_0_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_26 i_div_frac_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_53_32_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_25 i_div_exp_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(
        d1stg_step), .clk(rclk), .q(div_exp_in1_exp_eq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_24 i_div_exp_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        d1stg_step), .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (
        div_exp_in1_exp_neq_ffs) );
  dffe_SIZE1_23 i_div_frac_in2_51 ( .din(inq_in2_51), .en(d1stg_step), .clk(
        rclk), .q(div_frac_in2_51), .se(se), .si(1'b0) );
  dffe_SIZE1_22 i_div_frac_in2_54 ( .din(inq_in2_54), .en(d1stg_step), .clk(
        rclk), .q(div_frac_in2_54), .se(se), .si(1'b0) );
  dffe_SIZE1_21 i_div_frac_in2_53_0_neq_0 ( .din(inq_in2_53_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_53_0_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_20 i_div_frac_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_50_0_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_19 i_div_frac_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_53_32_neq_0), .se(se), .si(
        1'b0) );
  dffe_SIZE1_18 i_div_exp_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(
        d1stg_step), .clk(rclk), .q(div_exp_in2_exp_eq_0), .se(se), .si(1'b0)
         );
  dffe_SIZE1_17 i_div_exp_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        d1stg_step), .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (
        div_exp_in2_exp_neq_ffs) );
  dff_SIZE1_28 i_d2stg_denorm_sng_in2 ( .din(d1stg_denorm_sng_in2), .clk(rclk), 
        .q(d2stg_denorm_sng_in2), .se(se), .si(1'b0) );
  dff_SIZE1_27 i_d2stg_denorm_dbl_in2 ( .din(d1stg_denorm_dbl_in2), .clk(rclk), 
        .q(d2stg_denorm_dbl_in2), .se(se), .si(1'b0) );
  dff_SIZE1_26 i_d2stg_norm_sng_in2 ( .din(d1stg_norm_sng_in2), .clk(rclk), 
        .q(d2stg_norm_sng_in2), .se(se), .si(1'b0) );
  dff_SIZE1_25 i_d2stg_norm_dbl_in2 ( .din(d1stg_norm_dbl_in2), .clk(rclk), 
        .q(d2stg_norm_dbl_in2), .se(se), .si(1'b0) );
  dff_SIZE1_24 i_d2stg_snan_in1 ( .din(d1stg_snan_in1), .clk(rclk), .q(
        d2stg_snan_in1), .se(se), .si(1'b0) );
  dff_SIZE1_23 i_d2stg_snan_in2 ( .din(d1stg_snan_in2), .clk(rclk), .se(se), 
        .si(1'b0), .\q[0]_BAR (d2stg_snan_in2) );
  dff_SIZE1_22 i_d2stg_qnan_in1 ( .din(d1stg_qnan_in1), .clk(rclk), .q(
        d2stg_qnan_in1), .se(se), .si(1'b0) );
  dff_SIZE1_21 i_d2stg_qnan_in2 ( .din(d1stg_qnan_in2), .clk(rclk), .se(se), 
        .si(1'b0), .\q[0] (d2stg_qnan_in2) );
  dff_SIZE1_20 i_d2stg_nan_in2 ( .din(d1stg_nan_in2), .clk(rclk), .se(se), 
        .si(1'b0), .\q[0]_BAR (d2stg_nan_in2) );
  dff_SIZE1_19 i_d2stg_nan_in ( .din(d1stg_nan_in), .clk(rclk), .q(
        d2stg_nan_in), .se(se), .si(1'b0) );
  dff_SIZE1_18 i_d2stg_inf_in1 ( .din(d1stg_inf_in1), .clk(rclk), .q(
        d2stg_inf_in1), .se(se), .si(1'b0) );
  dff_SIZE1_16 i_d2stg_2inf_in ( .din(d1stg_2inf_in), .clk(rclk), .q(
        d2stg_2inf_in), .se(se), .si(1'b0) );
  dff_SIZE1_13 i_d2stg_infnan_in ( .din(d1stg_infnan_in), .clk(rclk), .q(
        d2stg_infnan_in), .se(se), .si(1'b0) );
  dff_SIZE1_11 i_d2stg_zero_in2 ( .din(d1stg_zero_in2), .clk(rclk), .q(
        d2stg_zero_in2), .se(se), .si(1'b0) );
  dff_SIZE1_10 i_d2stg_zero_in ( .din(d1stg_zero_in), .clk(rclk), .q(
        d2stg_zero_in), .se(se), .si(1'b0) );
  dff_SIZE1_9 i_d2stg_2zero_in ( .din(d1stg_2zero_in), .clk(rclk), .q(
        d2stg_2zero_in), .se(se), .si(1'b0) );
  dffr_SIZE8 i_d1stg_op ( .din(d1stg_op_in), .clk(rclk), .rst(n148), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\q[7] (
        d1stg_op[7]), .\q[6] (d1stg_op[6]), .\q[5]_BAR (d1stg_op[5]), .\q[4] (
        d1stg_op[4]), .\q[3] (d1stg_op[3]), .\q[2] (d1stg_op[2]), .\q[1] (
        d1stg_op[1]), .\q[0] (d1stg_op[0]) );
  dffr_SIZE1_3 i_d1stg_div ( .din(d1stg_div_in), .clk(rclk), .rst(n148), .q(
        d1stg_div), .se(se), .si(1'b0) );
  dffe_SIZE5_3 i_d1stg_sngopa ( .din({1'b0, 1'b0, 1'b0, 1'b0, inq_op[0]}), 
        .en(n183), .clk(rclk), .q(d1stg_sngopa), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffe_SIZE1_16 i_d1stg_dblop ( .din(inq_op[1]), .en(n183), .clk(rclk), .q(
        d1stg_dblop), .se(se), .si(1'b0) );
  dffe_SIZE5_2 i_d1stg_dblopa ( .din({1'b0, 1'b0, 1'b0, 1'b0, inq_op[1]}), 
        .en(n183), .clk(rclk), .q(d1stg_dblopa), .se(se), .si({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}) );
  dffr_SIZE3_0 i_d2stg_opdec ( .din({\d1stg_opdec[2] , n150, n151}), .clk(rclk), .rst(n148), .q({\d2stg_opdec[2] , div_expadd1_in2_exp_in2_sng, 
        div_expadd1_in2_exp_in2_dbl}), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dffr_SIZE1_2 i_d234stg_fdiv ( .din(d234stg_fdiv_in), .clk(rclk), .rst(n148), 
        .q(d234stg_fdiv), .se(se), .si(1'b0) );
  dffr_SIZE3_4 i_d3stg_opdec ( .din({\d2stg_opdec[2] , 
        div_expadd1_in2_exp_in2_sng, div_expadd1_in2_exp_in2_dbl}), .clk(rclk), 
        .rst(n148), .q({d3stg_fdiv, d3stg_opdec}), .se(se), .si({1'b0, 1'b0, 
        1'b0}) );
  dffr_SIZE3_3 i_d4stg_opdec ( .din({d3stg_fdiv, d3stg_opdec}), .clk(rclk), 
        .rst(n148), .q({d4stg_fdiv, d4stg_opdec}), .se(se), .si({1'b0, 1'b0, 
        1'b0}) );
  dffre_SIZE3_2 i_d5stg_opdec ( .din({d4stg_fdiv, d4stg_opdec}), .rst(n148), 
        .en(d5stg_step), .clk(rclk), .q({\d5stg_opdec[2] , d5stg_fdivs, 
        d5stg_fdivd}), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_7 i_d5stg_fdiva ( .din(d4stg_fdiv), .rst(n148), .en(d5stg_step), 
        .clk(rclk), .q(d5stg_fdiva), .se(se), .si(1'b0) );
  dff_SIZE1_8 i_d5stg_fdivb ( .din(d5stg_fdivb_in), .clk(rclk), .q(d5stg_fdivb), .se(se), .si(1'b0) );
  dffr_SIZE3_2 i_d6stg_opdec ( .din(d6stg_opdec_in), .clk(rclk), .rst(n148), 
        .q({d6stg_fdiv, d6stg_fdivs, d6stg_fdivd}), .se(se), .si({1'b0, 1'b0, 
        1'b0}) );
  dffr_SIZE3_1 i_d7stg_opdec ( .din({d6stg_fdiv, d6stg_fdivs, d6stg_fdivd}), 
        .clk(rclk), .rst(n148), .q({d7stg_fdiv, \d7stg_opdec[1] , d7stg_fdivd}), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE3_1 i_d8stg_opdec ( .din({d7stg_fdiv, \d7stg_opdec[1] , 
        d7stg_fdivd}), .rst(n148), .en(n156), .clk(rclk), .q({\d8stg_opdec[2] , 
        d8stg_fdivs, d8stg_fdivd}), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dffre_SIZE1_6 i_div_pipe_active ( .din(div_pipe_active_in), .rst(n148), .en(
        1'b1), .clk(rclk), .q(div_pipe_active), .se(se), .si(1'b0) );
  dffe_SIZE2_2 i_d1stg_rnd_mode ( .din(inq_rnd_mode), .en(n183), .clk(rclk), 
        .q(d1stg_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dffe_SIZE5_1 i_d1stg_id ( .din(inq_id), .en(n183), .clk(rclk), .q(d1stg_id), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE1_15 i_d1stg_sign1 ( .din(inq_in1_63), .en(n183), .clk(rclk), .q(
        d1stg_sign1), .se(se), .si(1'b0) );
  dffe_SIZE1_14 i_d1stg_sign2 ( .din(inq_in2_63), .en(n183), .clk(rclk), .q(
        d1stg_sign2), .se(se), .si(1'b0) );
  dffe_SIZE2_1 i_div_rnd_mode ( .din(d1stg_rnd_mode), .en(div_bkend_step), 
        .clk(rclk), .q(div_rnd_mode), .se(se), .si({1'b0, 1'b0}) );
  dff_SIZE10_1 i_div_id_out ( .din(div_id_out_in), .clk(rclk), .q(div_id_out), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE1_13 i_div_sign_out ( .din(d1stg_sign), .en(div_bkend_step), .clk(
        rclk), .q(div_sign_out), .se(se), .si(1'b0) );
  dffre_SIZE6_1 i_div_cnt ( .din(div_cnt_in), .rst(n148), .en(div_cnt_step), 
        .clk(rclk), .q(div_cnt), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffre_SIZE1_5 i_divs_cnt_lt_23 ( .din(divs_cnt_lt_23_in), .rst(n148), .en(
        div_cnt_lt_step), .clk(rclk), .q(divs_cnt_lt_23), .se(se), .si(1'b0)
         );
  dffre_SIZE1_4 i_divs_cnt_lt_23a ( .din(divs_cnt_lt_23_in), .rst(n148), .en(
        div_cnt_lt_step), .clk(rclk), .q(divs_cnt_lt_23a), .se(se), .si(1'b0)
         );
  dffre_SIZE1_3 i_divd_cnt_lt_52 ( .din(divd_cnt_lt_52_in), .rst(n148), .en(
        div_cnt_lt_step), .clk(rclk), .q(divd_cnt_lt_52), .se(se), .si(1'b0)
         );
  dffre_SIZE1_2 i_divd_cnt_lt_52a ( .din(divd_cnt_lt_52_in), .rst(n148), .en(
        div_cnt_lt_step), .clk(rclk), .q(divd_cnt_lt_52a), .se(se), .si(1'b0)
         );
  dffe_SIZE1_12 i_div_of_mask ( .din(n149), .en(div_bkend_step), .clk(rclk), 
        .q(div_of_mask), .se(se), .si(1'b0) );
  dffe_SIZE1_11 i_div_nv_out ( .din(div_nv_out_in), .en(div_bkend_step), .clk(
        rclk), .q(div_exc_out[4]), .se(se), .si(1'b0) );
  dffe_SIZE1_10 i_div_dz_out ( .din(div_dz_out_in), .en(div_bkend_step), .clk(
        rclk), .q(div_exc_out[1]), .se(se), .si(1'b0) );
  dffe_SIZE1_9 i_div_of_out_tmp1 ( .din(div_of_out_tmp1_in), .en(d7stg_fdiv), 
        .clk(rclk), .q(div_of_out_tmp1), .se(se), .si(1'b0) );
  dffe_SIZE1_8 i_div_of_out_tmp2 ( .din(d7stg_in_of), .en(d7stg_fdiv), .clk(
        rclk), .q(div_of_out_tmp2), .se(se), .si(1'b0) );
  dffe_SIZE1_7 i_div_out_52_inv ( .din(div_frac_add_52_inva), .en(d7stg_fdiv), 
        .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (div_out_52_inv) );
  dffe_SIZE1_6 i_div_uf_out ( .din(div_uf_out_in), .en(d7stg_fdiv), .clk(rclk), 
        .q(div_exc_out[2]), .se(se), .si(1'b0) );
  dffe_SIZE1_5 i_div_nx_out ( .din(div_nx_out_in), .en(d7stg_fdiv), .clk(rclk), 
        .q(div_nx_out), .se(se), .si(1'b0) );
  dffe_SIZE1_4 i_d7stg_lsb ( .din(d7stg_lsb_in), .en(d6stg_fdiv), .clk(rclk), 
        .se(se), .si(1'b0), .\q[0]_BAR (d7stg_lsb) );
  dffe_SIZE1_3 i_d7stg_grd ( .din(d7stg_grd_in), .en(d6stg_fdiv), .clk(rclk), 
        .q(d7stg_grd), .se(se), .si(1'b0) );
  dffe_SIZE1_2 i_d7stg_stk ( .din(d7stg_stk_in), .en(d6stg_fdiv), .clk(rclk), 
        .q(d7stg_stk), .se(se), .si(1'b0) );
  dff_SIZE1_7 i_div_expadd1_in1_dbl ( .din(div_expadd1_in1_dbl_in), .clk(rclk), 
        .q(div_expadd1_in1_dbl), .se(se), .si(1'b0) );
  dff_SIZE1_6 i_div_expadd1_in1_sng ( .din(div_expadd1_in1_sng_in), .clk(rclk), 
        .q(div_expadd1_in1_sng), .se(se), .si(1'b0) );
  dffr_SIZE1_1 i_div_expadd2_in1_exp_out ( .din(div_expadd2_in1_exp_out_in), 
        .clk(rclk), .rst(n148), .q(div_expadd2_in1_exp_out), .se(se), .si(1'b0) );
  dffe_SIZE1_1 i_div_expadd2_no_decr_inv ( .din(n154), .en(
        div_expadd2_no_decr_load), .clk(rclk), .q(div_expadd2_no_decr_inv), 
        .se(se), .si(1'b0) );
  INVX0_RVT U3 ( .A(d5stg_step), .Y(n87) );
  INVX0_RVT U4 ( .A(n157), .Y(d7stg_in_of) );
  INVX0_RVT U5 ( .A(div_frac_add_in1_neq_0), .Y(n131) );
  OR3X1_RVT U6 ( .A1(d3stg_fdiv), .A2(\d2stg_opdec[2] ), .A3(\d1stg_opdec[2] ), 
        .Y(d234stg_fdiv_in) );
  INVX0_RVT U7 ( .A(div_exp_out[0]), .Y(n129) );
  INVX0_RVT U8 ( .A(div_exp1[2]), .Y(n165) );
  INVX0_RVT U9 ( .A(div_exp1[3]), .Y(n168) );
  INVX0_RVT U10 ( .A(div_exp1[5]), .Y(n164) );
  OR3X1_RVT U11 ( .A1(div_exp1[8]), .A2(div_exp1[11]), .A3(div_exp1[7]), .Y(
        n49) );
  INVX0_RVT U12 ( .A(div_exp1[12]), .Y(n141) );
  INVX0_RVT U13 ( .A(n66), .Y(d1stg_inf_in1) );
  INVX0_RVT U14 ( .A(n117), .Y(n118) );
  INVX0_RVT U15 ( .A(n116), .Y(n119) );
  INVX0_RVT U16 ( .A(n107), .Y(div_expadd2_no_decr_load) );
  INVX0_RVT U17 ( .A(n125), .Y(d1stg_snan_sng_in1) );
  INVX0_RVT U18 ( .A(n126), .Y(d1stg_snan_dbl_in1) );
  INVX0_RVT U19 ( .A(n123), .Y(d1stg_snan_sng_in2) );
  INVX0_RVT U20 ( .A(n124), .Y(d1stg_snan_dbl_in2) );
  INVX1_RVT U21 ( .A(d7stg_to_0_inv), .Y(d7stg_to_0) );
  INVX1_RVT U22 ( .A(n156), .Y(n65) );
  INVX0_RVT U23 ( .A(n136), .Y(d1stg_zero_in2) );
  INVX0_RVT U24 ( .A(n78), .Y(n79) );
  OR3X2_RVT U25 ( .A1(div_cnt[2]), .A2(div_cnt[3]), .A3(n108), .Y(n109) );
  OR3X1_RVT U26 ( .A1(n14), .A2(div_frac_in2_51), .A3(div_frac_in2_50_0_neq_0), 
        .Y(n13) );
  INVX0_RVT U27 ( .A(n183), .Y(n152) );
  INVX1_RVT U28 ( .A(div_cnt[2]), .Y(n75) );
  INVX0_RVT U29 ( .A(div_cnt[4]), .Y(n80) );
  INVX0_RVT U30 ( .A(d5stg_fdivs), .Y(n169) );
  INVX1_RVT U31 ( .A(div_cnt[5]), .Y(n51) );
  INVX0_RVT U32 ( .A(div_nx_out_in), .Y(n130) );
  OR3X1_RVT U33 ( .A1(div_frac_in1_54), .A2(div_frac_in1_53_0_neq_0), .A3(n38), 
        .Y(n135) );
  OR3X1_RVT U34 ( .A1(div_frac_in2_54), .A2(div_frac_in2_53_0_neq_0), .A3(n83), 
        .Y(n136) );
  INVX0_RVT U35 ( .A(d4stg_fdiv), .Y(n146) );
  INVX1_RVT U36 ( .A(d6stg_fdivd), .Y(n143) );
  INVX0_RVT U37 ( .A(d1stg_op[0]), .Y(n24) );
  INVX0_RVT U38 ( .A(div_rnd_mode[1]), .Y(n1) );
  OR3X1_RVT U39 ( .A1(d2stg_zero_in2), .A2(d2stg_nan_in), .A3(d2stg_inf_in1), 
        .Y(n153) );
  INVX1_RVT U40 ( .A(div_rnd_mode[0]), .Y(n3) );
  INVX1_RVT U41 ( .A(div_sign_out), .Y(n2) );
  INVX0_RVT U42 ( .A(\d7stg_opdec[1] ), .Y(n11) );
  INVX0_RVT U43 ( .A(d7stg_fdiv), .Y(n163) );
  INVX0_RVT U44 ( .A(d6stg_fdiv), .Y(n142) );
  INVX0_RVT U45 ( .A(d1stg_op[1]), .Y(n25) );
  INVX0_RVT U46 ( .A(div_frac_in1_54), .Y(n37) );
  INVX0_RVT U47 ( .A(div_frac_in1_51), .Y(n30) );
  INVX0_RVT U48 ( .A(div_frac_in2_54), .Y(n35) );
  INVX0_RVT U49 ( .A(div_frac_in2_51), .Y(n28) );
  INVX0_RVT U50 ( .A(div_exp_in2_exp_neq_ffs), .Y(n137) );
  NAND3X0_RVT U51 ( .A1(d7stg_grd), .A2(n1), .A3(n3), .Y(n7) );
  INVX1_RVT U52 ( .A(d7stg_stk), .Y(n6) );
  AO22X1_RVT U53 ( .A1(div_rnd_mode[0]), .A2(div_sign_out), .A3(n3), .A4(n2), 
        .Y(n4) );
  OR2X1_RVT U54 ( .A1(d7stg_stk), .A2(d7stg_grd), .Y(div_nx_out_in) );
  NAND3X0_RVT U55 ( .A1(div_rnd_mode[1]), .A2(n4), .A3(div_nx_out_in), .Y(n5)
         );
  OA221X1_RVT U56 ( .A1(n7), .A2(d7stg_lsb), .A3(n7), .A4(n6), .A5(n5), .Y(
        d7stg_rndup_inv) );
  INVX1_RVT U57 ( .A(div_exp_out[12]), .Y(n158) );
  OR4X1_RVT U58 ( .A1(div_exp_out[10]), .A2(div_exp_out[9]), .A3(
        div_exp_out[8]), .A4(div_exp_out[11]), .Y(n68) );
  NAND4X0_RVT U59 ( .A1(d7stg_fdivd), .A2(div_exp_out[10]), .A3(div_exp_out[9]), .A4(div_exp_out[8]), .Y(n10) );
  AND4X1_RVT U60 ( .A1(div_exp_out[2]), .A2(div_exp_out[1]), .A3(
        div_exp_out[7]), .A4(div_exp_out[4]), .Y(n8) );
  NAND4X0_RVT U61 ( .A1(div_exp_out[6]), .A2(div_exp_out[5]), .A3(
        div_exp_out[3]), .A4(n8), .Y(n9) );
  AOI21X1_RVT U62 ( .A1(n11), .A2(n10), .A3(n9), .Y(n127) );
  AO222X1_RVT U63 ( .A1(n68), .A2(\d7stg_opdec[1] ), .A3(n127), .A4(
        div_exp_out[0]), .A5(d7stg_fdivd), .A6(div_exp_out[11]), .Y(n12) );
  NAND3X0_RVT U64 ( .A1(div_of_mask), .A2(n158), .A3(n12), .Y(n157) );
  AND3X1_RVT U65 ( .A1(d7stg_fdiv), .A2(d7stg_rndup_inv), .A3(n157), .Y(
        div_frac_out_add_in1) );
  INVX1_RVT U66 ( .A(d7stg_rndup_inv), .Y(n162) );
  AND3X1_RVT U67 ( .A1(d7stg_fdiv), .A2(n157), .A3(n162), .Y(div_frac_out_add)
         );
  NAND2X0_RVT U68 ( .A1(\d8stg_opdec[2] ), .A2(div_dest_rdy), .Y(n156) );
  OA21X1_RVT U69 ( .A1(n65), .A2(d7stg_fdiv), .A3(div_ctl_rst_l), .Y(
        d8stg_fdiv_in) );
  INVX1_RVT U70 ( .A(div_exp_in2_exp_eq_0), .Y(n83) );
  INVX1_RVT U71 ( .A(div_exp_in1_exp_eq_0), .Y(n38) );
  INVX1_RVT U72 ( .A(d1stg_dblopa[2]), .Y(n14) );
  INVX1_RVT U73 ( .A(d1stg_sngopa[2]), .Y(n15) );
  OR2X1_RVT U74 ( .A1(div_frac_in2_53_32_neq_0), .A2(div_frac_in2_54), .Y(n19)
         );
  AO221X1_RVT U75 ( .A1(n13), .A2(n15), .A3(n13), .A4(n19), .A5(n137), .Y(n29)
         );
  OR2X1_RVT U76 ( .A1(div_frac_in1_54), .A2(div_frac_in1_53_32_neq_0), .Y(n18)
         );
  OR2X1_RVT U77 ( .A1(div_frac_in1_50_0_neq_0), .A2(div_frac_in1_51), .Y(n17)
         );
  OAI22X1_RVT U78 ( .A1(n15), .A2(n18), .A3(n14), .A4(n17), .Y(n16) );
  NAND2X0_RVT U79 ( .A1(div_exp_in1_exp_neq_ffs), .A2(n16), .Y(n66) );
  AND4X1_RVT U80 ( .A1(n136), .A2(n135), .A3(n29), .A4(n66), .Y(n27) );
  AO22X1_RVT U81 ( .A1(d1stg_sngopa[2]), .A2(n18), .A3(d1stg_dblopa[2]), .A4(
        n17), .Y(n21) );
  OA21X1_RVT U82 ( .A1(div_frac_in2_51), .A2(div_frac_in2_50_0_neq_0), .A3(
        d1stg_dblopa[2]), .Y(n20) );
  OA221X1_RVT U83 ( .A1(n20), .A2(d1stg_sngopa[2]), .A3(n20), .A4(n19), .A5(
        div_exp_in2_exp_neq_ffs), .Y(d1stg_nan_in2) );
  AO21X1_RVT U84 ( .A1(div_exp_in1_exp_neq_ffs), .A2(n21), .A3(d1stg_nan_in2), 
        .Y(d1stg_nan_in) );
  NAND2X0_RVT U85 ( .A1(d1stg_op[6]), .A2(d1stg_op[2]), .Y(n22) );
  NOR3X0_RVT U86 ( .A1(d1stg_op[4]), .A2(d1stg_op[7]), .A3(n22), .Y(n23) );
  AND3X1_RVT U87 ( .A1(d1stg_op[5]), .A2(d1stg_op[3]), .A3(n23), .Y(n26) );
  AND3X1_RVT U88 ( .A1(n26), .A2(d1stg_op[1]), .A3(n24), .Y(n151) );
  AND3X1_RVT U89 ( .A1(d1stg_op[0]), .A2(n26), .A3(n25), .Y(n150) );
  OR2X1_RVT U90 ( .A1(n151), .A2(n150), .Y(\d1stg_opdec[2] ) );
  OA21X1_RVT U91 ( .A1(n27), .A2(d1stg_nan_in), .A3(\d1stg_opdec[2] ), .Y(n36)
         );
  NAND4X0_RVT U92 ( .A1(d1stg_dblopa[1]), .A2(div_exp_in2_exp_neq_ffs), .A3(
        div_frac_in2_50_0_neq_0), .A4(n28), .Y(n124) );
  AND3X1_RVT U93 ( .A1(n36), .A2(d1stg_dblopa[0]), .A3(n124), .Y(n31) );
  NAND3X0_RVT U94 ( .A1(d1stg_dblopa[1]), .A2(div_frac_in2_51), .A3(
        div_exp_in2_exp_neq_ffs), .Y(n86) );
  AND3X1_RVT U95 ( .A1(div_exp_in1_exp_eq_0), .A2(n31), .A3(n86), .Y(
        div_norm_frac_in1_dbl_dnrm) );
  NOR2X0_RVT U96 ( .A1(n29), .A2(n66), .Y(d1stg_2inf_in) );
  NOR2X0_RVT U97 ( .A1(n136), .A2(n135), .Y(d1stg_2zero_in) );
  OA21X1_RVT U98 ( .A1(d1stg_2inf_in), .A2(d1stg_2zero_in), .A3(
        \d1stg_opdec[2] ), .Y(div_norm_qnan) );
  NAND4X0_RVT U99 ( .A1(d1stg_dblopa[1]), .A2(div_exp_in1_exp_neq_ffs), .A3(
        div_frac_in1_50_0_neq_0), .A4(n30), .Y(n126) );
  NAND4X0_RVT U100 ( .A1(d1stg_dblopa[1]), .A2(div_frac_in2_51), .A3(
        div_exp_in2_exp_neq_ffs), .A4(n126), .Y(n33) );
  AND3X1_RVT U101 ( .A1(n31), .A2(n38), .A3(n33), .Y(
        div_norm_frac_in1_dbl_norm) );
  OR2X1_RVT U102 ( .A1(d2stg_infnan_in), .A2(d2stg_zero_in), .Y(n140) );
  INVX1_RVT U103 ( .A(n140), .Y(n32) );
  AND2X1_RVT U104 ( .A1(\d2stg_opdec[2] ), .A2(n32), .Y(n43) );
  NAND2X0_RVT U105 ( .A1(n33), .A2(n124), .Y(n34) );
  AO22X1_RVT U106 ( .A1(d2stg_norm_dbl_in2), .A2(n43), .A3(\d1stg_opdec[2] ), 
        .A4(n34), .Y(div_norm_frac_in2_dbl_norm) );
  AND2X1_RVT U107 ( .A1(n43), .A2(d2stg_denorm_dbl_in2), .Y(
        div_norm_frac_in2_dbl_dnrm) );
  NAND3X0_RVT U108 ( .A1(d5stg_fdivd), .A2(n156), .A3(n141), .Y(n145) );
  INVX1_RVT U109 ( .A(n145), .Y(div_frac_out_shl1_dbl) );
  NAND4X0_RVT U110 ( .A1(div_frac_in2_53_32_neq_0), .A2(
        div_exp_in2_exp_neq_ffs), .A3(d1stg_sngopa[1]), .A4(n35), .Y(n123) );
  AND3X1_RVT U111 ( .A1(n36), .A2(d1stg_sngopa[0]), .A3(n123), .Y(n42) );
  NAND4X0_RVT U112 ( .A1(div_exp_in1_exp_neq_ffs), .A2(
        div_frac_in1_53_32_neq_0), .A3(d1stg_sngopa[1]), .A4(n37), .Y(n125) );
  NAND4X0_RVT U113 ( .A1(div_frac_in2_54), .A2(div_exp_in2_exp_neq_ffs), .A3(
        d1stg_sngopa[1]), .A4(n125), .Y(n40) );
  AND3X1_RVT U114 ( .A1(n42), .A2(n38), .A3(n40), .Y(
        div_norm_frac_in1_sng_norm) );
  NAND2X0_RVT U115 ( .A1(\d5stg_opdec[2] ), .A2(n156), .Y(n107) );
  INVX1_RVT U116 ( .A(div_cnt[0]), .Y(n111) );
  AND2X1_RVT U117 ( .A1(div_expadd2_no_decr_load), .A2(n111), .Y(div_cnt_in[0]) );
  INVX1_RVT U118 ( .A(div_cnt[1]), .Y(n106) );
  INVX1_RVT U119 ( .A(div_cnt[3]), .Y(n54) );
  NAND3X0_RVT U120 ( .A1(div_cnt_in[0]), .A2(n106), .A3(n54), .Y(n39) );
  NOR4X1_RVT U121 ( .A1(div_cnt[4]), .A2(div_cnt[2]), .A3(div_cnt[5]), .A4(n39), .Y(div_bkend_step) );
  NAND2X0_RVT U122 ( .A1(n40), .A2(n123), .Y(n41) );
  AO22X1_RVT U123 ( .A1(d2stg_norm_sng_in2), .A2(n43), .A3(\d1stg_opdec[2] ), 
        .A4(n41), .Y(div_norm_frac_in2_sng_norm) );
  NAND3X0_RVT U124 ( .A1(div_exp_in2_exp_neq_ffs), .A2(div_frac_in2_54), .A3(
        d1stg_sngopa[1]), .Y(n85) );
  AND3X1_RVT U125 ( .A1(div_exp_in1_exp_eq_0), .A2(n42), .A3(n85), .Y(
        div_norm_frac_in1_sng_dnrm) );
  AND2X1_RVT U126 ( .A1(n43), .A2(d2stg_denorm_sng_in2), .Y(
        div_norm_frac_in2_sng_dnrm) );
  NOR4X1_RVT U127 ( .A1(d1stg_div), .A2(d234stg_fdiv), .A3(divs_cnt_lt_23a), 
        .A4(divd_cnt_lt_52a), .Y(n183) );
  AND2X1_RVT U128 ( .A1(n183), .A2(inq_div), .Y(d1stg_div_in) );
  OR4X1_RVT U129 ( .A1(\d1stg_opdec[2] ), .A2(d4stg_fdiv), .A3(d3stg_fdiv), 
        .A4(n43), .Y(div_exp1_expadd1) );
  NOR4X1_RVT U130 ( .A1(d1stg_div), .A2(d234stg_fdiv), .A3(divs_cnt_lt_23), 
        .A4(divd_cnt_lt_52), .Y(d1stg_step) );
  INVX1_RVT U131 ( .A(div_ctl_rst_l), .Y(n148) );
  NAND2X0_RVT U132 ( .A1(div_cnt[5]), .A2(d5stg_fdivd), .Y(n45) );
  AOI222X1_RVT U133 ( .A1(div_cnt[3]), .A2(div_cnt[2]), .A3(div_cnt[3]), .A4(
        n169), .A5(n54), .A6(n45), .Y(n47) );
  NAND2X0_RVT U134 ( .A1(div_cnt[0]), .A2(div_cnt[5]), .Y(n46) );
  NAND3X0_RVT U135 ( .A1(n47), .A2(div_cnt[4]), .A3(n46), .Y(n48) );
  AO221X1_RVT U136 ( .A1(div_cnt[1]), .A2(n75), .A3(n106), .A4(n111), .A5(n48), 
        .Y(n62) );
  NOR4X1_RVT U137 ( .A1(div_exp1[6]), .A2(div_exp1[10]), .A3(div_exp1[9]), 
        .A4(n49), .Y(n173) );
  AOI22X1_RVT U138 ( .A1(n51), .A2(div_exp1[5]), .A3(n80), .A4(div_exp1[4]), 
        .Y(n50) );
  OA221X1_RVT U139 ( .A1(n80), .A2(div_exp1[4]), .A3(n51), .A4(div_exp1[5]), 
        .A5(n50), .Y(n60) );
  INVX1_RVT U140 ( .A(div_exp1[1]), .Y(n170) );
  INVX1_RVT U141 ( .A(div_exp1[0]), .Y(n167) );
  OA22X1_RVT U142 ( .A1(div_cnt[1]), .A2(n170), .A3(div_cnt[0]), .A4(n167), 
        .Y(n52) );
  OA221X1_RVT U143 ( .A1(n111), .A2(div_exp1[0]), .A3(n106), .A4(div_exp1[1]), 
        .A5(n52), .Y(n59) );
  OA22X1_RVT U144 ( .A1(div_cnt[2]), .A2(n165), .A3(div_cnt[3]), .A4(n168), 
        .Y(n53) );
  OA221X1_RVT U145 ( .A1(n75), .A2(div_exp1[2]), .A3(n54), .A4(div_exp1[3]), 
        .A5(n53), .Y(n57) );
  NOR4X1_RVT U146 ( .A1(div_exp1[2]), .A2(div_exp1[5]), .A3(div_exp1[3]), .A4(
        div_exp1[4]), .Y(n55) );
  NAND4X0_RVT U147 ( .A1(n55), .A2(n107), .A3(n170), .A4(n167), .Y(n56) );
  AND4X1_RVT U148 ( .A1(\d5stg_opdec[2] ), .A2(n57), .A3(n56), .A4(n141), .Y(
        n58) );
  NAND4X0_RVT U149 ( .A1(n173), .A2(n60), .A3(n59), .A4(n58), .Y(n61) );
  AND2X1_RVT U150 ( .A1(n62), .A2(n61), .Y(n64) );
  NAND2X0_RVT U151 ( .A1(div_exp1[12]), .A2(div_expadd2_no_decr_load), .Y(n63)
         );
  AND2X1_RVT U152 ( .A1(n64), .A2(n63), .Y(n115) );
  NAND2X0_RVT U153 ( .A1(\d5stg_opdec[2] ), .A2(n115), .Y(d5stg_step) );
  NAND2X0_RVT U154 ( .A1(n65), .A2(n87), .Y(div_cnt_lt_step) );
  NAND2X0_RVT U155 ( .A1(div_sign_out), .A2(div_rnd_mode[1]), .Y(n67) );
  HADDX1_RVT U156 ( .A0(div_rnd_mode[0]), .B0(n67), .SO(d7stg_to_0_inv) );
  NAND3X0_RVT U157 ( .A1(d5stg_fdivs), .A2(n156), .A3(n141), .Y(n144) );
  INVX1_RVT U158 ( .A(n144), .Y(div_frac_out_shl1_sng) );
  INVX1_RVT U159 ( .A(div_bkend_step), .Y(n103) );
  NAND2X0_RVT U160 ( .A1(n142), .A2(n103), .Y(n161) );
  INVX1_RVT U161 ( .A(n161), .Y(div_exp_out_expadd22_inv) );
  NOR4X1_RVT U162 ( .A1(div_exp_out[2]), .A2(div_exp_out[1]), .A3(
        div_exp_out[7]), .A4(div_exp_out[4]), .Y(n70) );
  NOR4X1_RVT U163 ( .A1(div_exp_out[6]), .A2(div_exp_out[5]), .A3(
        div_exp_out[3]), .A4(n68), .Y(n69) );
  AND2X1_RVT U164 ( .A1(n70), .A2(n69), .Y(n128) );
  OR3X2_RVT U165 ( .A1(div_exp_out[12]), .A2(n128), .A3(div_frac_out_54), .Y(
        d6stg_frac_out_nosh) );
  AND2X1_RVT U174 ( .A1(n135), .A2(d1stg_zero_in2), .Y(n73) );
  NOR2X0_RVT U175 ( .A1(d1stg_dblopa[3]), .A2(d1stg_sngopa[3]), .Y(n138) );
  INVX1_RVT U176 ( .A(n138), .Y(n71) );
  NAND2X0_RVT U177 ( .A1(n71), .A2(div_exp_in1_exp_neq_ffs), .Y(n72) );
  AND2X1_RVT U178 ( .A1(n73), .A2(n72), .Y(div_dz_out_in) );
  NAND3X0_RVT U179 ( .A1(div_cnt[0]), .A2(div_cnt[2]), .A3(div_cnt[1]), .Y(
        n105) );
  AND2X1_RVT U180 ( .A1(n105), .A2(div_expadd2_no_decr_load), .Y(n77) );
  AND2X1_RVT U181 ( .A1(div_cnt[0]), .A2(div_cnt[1]), .Y(n108) );
  INVX1_RVT U182 ( .A(n108), .Y(n74) );
  NAND2X0_RVT U183 ( .A1(n75), .A2(n74), .Y(n76) );
  AND2X1_RVT U184 ( .A1(n77), .A2(n76), .Y(div_cnt_in[2]) );
  AND4X1_RVT U185 ( .A1(div_cnt[0]), .A2(div_cnt[2]), .A3(div_cnt[1]), .A4(
        div_cnt[3]), .Y(n78) );
  NAND2X0_RVT U186 ( .A1(div_cnt[4]), .A2(n78), .Y(n104) );
  AND2X1_RVT U187 ( .A1(n104), .A2(div_expadd2_no_decr_load), .Y(n82) );
  NAND2X0_RVT U188 ( .A1(n80), .A2(n79), .Y(n81) );
  AND2X1_RVT U189 ( .A1(n82), .A2(n81), .Y(div_cnt_in[4]) );
  AND2X1_RVT U190 ( .A1(div_exp_in2_exp_eq_0), .A2(d1stg_sngopa[0]), .Y(
        d1stg_denorm_sng_in2) );
  AND2X1_RVT U191 ( .A1(div_exp_in2_exp_eq_0), .A2(d1stg_dblopa[0]), .Y(
        d1stg_denorm_dbl_in2) );
  AND2X1_RVT U192 ( .A1(d1stg_sngopa[0]), .A2(n83), .Y(d1stg_norm_sng_in2) );
  AND2X1_RVT U193 ( .A1(d1stg_dblopa[0]), .A2(n83), .Y(d1stg_norm_dbl_in2) );
  AO22X1_RVT U194 ( .A1(d1stg_dblopa[1]), .A2(div_frac_in1_51), .A3(
        div_frac_in1_54), .A4(d1stg_sngopa[1]), .Y(n84) );
  AND2X1_RVT U195 ( .A1(div_exp_in1_exp_neq_ffs), .A2(n84), .Y(d1stg_qnan_in1)
         );
  NAND2X0_RVT U196 ( .A1(n86), .A2(n85), .Y(d1stg_qnan_in2) );
  AND2X1_RVT U197 ( .A1(d1stg_div_in), .A2(inq_op[7]), .Y(d1stg_op_in[7]) );
  AND2X1_RVT U198 ( .A1(d1stg_div_in), .A2(inq_op[6]), .Y(d1stg_op_in[6]) );
  AND2X1_RVT U199 ( .A1(d1stg_div_in), .A2(inq_op[5]), .Y(d1stg_op_in[5]) );
  AND2X1_RVT U200 ( .A1(d1stg_div_in), .A2(inq_op[4]), .Y(d1stg_op_in[4]) );
  AND2X1_RVT U201 ( .A1(d1stg_div_in), .A2(inq_op[3]), .Y(d1stg_op_in[3]) );
  AND2X1_RVT U202 ( .A1(d1stg_div_in), .A2(inq_op[2]), .Y(d1stg_op_in[2]) );
  AND2X1_RVT U203 ( .A1(inq_op[1]), .A2(d1stg_div_in), .Y(d1stg_op_in[1]) );
  AND2X1_RVT U204 ( .A1(inq_op[0]), .A2(d1stg_div_in), .Y(d1stg_op_in[0]) );
  OA21X1_RVT U207 ( .A1(d4stg_fdiv), .A2(n87), .A3(div_ctl_rst_l), .Y(
        d5stg_fdivb_in) );
  INVX1_RVT U208 ( .A(n115), .Y(n155) );
  AND2X1_RVT U209 ( .A1(d5stg_fdivs), .A2(n155), .Y(d6stg_opdec_in[1]) );
  AND2X1_RVT U210 ( .A1(d5stg_fdivd), .A2(n155), .Y(d6stg_opdec_in[0]) );
  OR2X1_RVT U211 ( .A1(d4stg_fdiv), .A2(d234stg_fdiv_in), .Y(div_exp1_load) );
  OR2X1_RVT U212 ( .A1(\d5stg_opdec[2] ), .A2(d7stg_fdiv), .Y(div_expadd2_cin)
         );
  OR4X1_RVT U213 ( .A1(d6stg_fdiv), .A2(\d8stg_opdec[2] ), .A3(div_exp1_load), 
        .A4(div_expadd2_cin), .Y(div_pipe_active_in) );
  AOI22X1_RVT U214 ( .A1(d2stg_snan_in1), .A2(d2stg_snan_in2), .A3(
        d2stg_nan_in2), .A4(d2stg_qnan_in1), .Y(n88) );
  NAND2X0_RVT U215 ( .A1(d1stg_sign2), .A2(n88), .Y(n93) );
  AND2X1_RVT U216 ( .A1(d1stg_sign1), .A2(d2stg_snan_in2), .Y(n91) );
  INVX1_RVT U217 ( .A(d2stg_snan_in1), .Y(n89) );
  NAND2X0_RVT U218 ( .A1(n89), .A2(d2stg_qnan_in2), .Y(n90) );
  AND2X1_RVT U219 ( .A1(n91), .A2(n90), .Y(n92) );
  HADDX1_RVT U220 ( .A0(n93), .B0(n92), .SO(n94) );
  NOR3X0_RVT U221 ( .A1(d2stg_2inf_in), .A2(d2stg_2zero_in), .A3(n94), .Y(
        d1stg_sign) );
  AND2X1_RVT U222 ( .A1(d1stg_id[2]), .A2(d1stg_id[4]), .Y(n95) );
  AND2X1_RVT U223 ( .A1(div_bkend_step), .A2(d1stg_id[3]), .Y(n99) );
  AO22X1_RVT U224 ( .A1(n95), .A2(n99), .A3(div_id_out[9]), .A4(n103), .Y(
        div_id_out_in[9]) );
  INVX1_RVT U225 ( .A(d1stg_id[2]), .Y(n98) );
  AND2X1_RVT U226 ( .A1(d1stg_id[4]), .A2(n98), .Y(n96) );
  AO22X1_RVT U227 ( .A1(n96), .A2(n99), .A3(div_id_out[8]), .A4(n103), .Y(
        div_id_out_in[8]) );
  NOR2X0_RVT U228 ( .A1(d1stg_id[3]), .A2(n103), .Y(n101) );
  AO22X1_RVT U229 ( .A1(n101), .A2(n95), .A3(div_id_out[7]), .A4(n103), .Y(
        div_id_out_in[7]) );
  AO22X1_RVT U230 ( .A1(n101), .A2(n96), .A3(div_id_out[6]), .A4(n103), .Y(
        div_id_out_in[6]) );
  INVX1_RVT U231 ( .A(d1stg_id[4]), .Y(n97) );
  AND2X1_RVT U232 ( .A1(d1stg_id[2]), .A2(n97), .Y(n100) );
  AO22X1_RVT U233 ( .A1(n100), .A2(n99), .A3(div_id_out[5]), .A4(n103), .Y(
        div_id_out_in[5]) );
  AND2X1_RVT U234 ( .A1(n98), .A2(n97), .Y(n102) );
  AO22X1_RVT U235 ( .A1(n102), .A2(n99), .A3(div_id_out[4]), .A4(n103), .Y(
        div_id_out_in[4]) );
  AO22X1_RVT U236 ( .A1(n100), .A2(n101), .A3(div_id_out[3]), .A4(n103), .Y(
        div_id_out_in[3]) );
  AO22X1_RVT U237 ( .A1(n102), .A2(n101), .A3(div_id_out[2]), .A4(n103), .Y(
        div_id_out_in[2]) );
  AO22X1_RVT U238 ( .A1(div_bkend_step), .A2(d1stg_id[1]), .A3(n103), .A4(
        div_id_out[1]), .Y(div_id_out_in[1]) );
  AO22X1_RVT U239 ( .A1(div_bkend_step), .A2(d1stg_id[0]), .A3(n103), .A4(
        div_id_out[0]), .Y(div_id_out_in[0]) );
  HADDX1_RVT U240 ( .A0(div_cnt[5]), .B0(n104), .SO(n116) );
  NOR2X0_RVT U241 ( .A1(n107), .A2(n116), .Y(div_cnt_in[5]) );
  HADDX1_RVT U242 ( .A0(div_cnt[3]), .B0(n105), .SO(n113) );
  NOR2X0_RVT U243 ( .A1(n107), .A2(n113), .Y(div_cnt_in[3]) );
  OA221X1_RVT U244 ( .A1(div_cnt[0]), .A2(div_cnt[1]), .A3(n111), .A4(n106), 
        .A5(div_expadd2_no_decr_load), .Y(div_cnt_in[1]) );
  NAND2X0_RVT U245 ( .A1(n107), .A2(n146), .Y(div_cnt_step) );
  NAND3X0_RVT U246 ( .A1(div_cnt[2]), .A2(div_cnt[3]), .A3(n108), .Y(n110) );
  NAND3X0_RVT U247 ( .A1(div_cnt[4]), .A2(n110), .A3(n109), .Y(n117) );
  NAND2X0_RVT U248 ( .A1(div_cnt[1]), .A2(n111), .Y(n112) );
  OA221X1_RVT U249 ( .A1(n117), .A2(n113), .A3(n117), .A4(n112), .A5(n116), 
        .Y(n114) );
  OA222X1_RVT U250 ( .A1(d4stg_opdec[1]), .A2(n115), .A3(d4stg_opdec[1]), .A4(
        d5stg_fdivs), .A5(d4stg_opdec[1]), .A6(n114), .Y(divs_cnt_lt_23_in) );
  AND2X1_RVT U251 ( .A1(d5stg_fdivd), .A2(n115), .Y(n121) );
  NAND2X0_RVT U252 ( .A1(n119), .A2(n118), .Y(n120) );
  AND2X1_RVT U253 ( .A1(n121), .A2(n120), .Y(n122) );
  OR2X1_RVT U254 ( .A1(d4stg_opdec[0]), .A2(n122), .Y(divd_cnt_lt_52_in) );
  NAND2X0_RVT U255 ( .A1(n124), .A2(n123), .Y(d1stg_snan_in2) );
  NAND2X0_RVT U256 ( .A1(n126), .A2(n125), .Y(d1stg_snan_in1) );
  OR4X1_RVT U257 ( .A1(d1stg_2inf_in), .A2(d1stg_2zero_in), .A3(d1stg_snan_in1), .A4(d1stg_snan_in2), .Y(div_nv_out_in) );
  AND4X1_RVT U258 ( .A1(n127), .A2(div_of_mask), .A3(n158), .A4(n162), .Y(
        div_of_out_tmp1_in) );
  AND2X1_RVT U259 ( .A1(n129), .A2(n128), .Y(n133) );
  NAND2X0_RVT U260 ( .A1(n131), .A2(n130), .Y(n132) );
  AND2X1_RVT U261 ( .A1(n133), .A2(n132), .Y(n134) );
  OA21X1_RVT U262 ( .A1(div_exp_out[12]), .A2(n134), .A3(div_of_mask), .Y(
        div_uf_out_in) );
  AO21X1_RVT U263 ( .A1(div_of_out_tmp1), .A2(div_out_52_inv), .A3(
        div_of_out_tmp2), .Y(div_exc_out[3]) );
  OR2X1_RVT U264 ( .A1(div_nx_out), .A2(div_exc_out[3]), .Y(div_exc_out[0]) );
  NAND2X0_RVT U265 ( .A1(n136), .A2(n135), .Y(d1stg_zero_in) );
  AO221X1_RVT U266 ( .A1(d1stg_inf_in1), .A2(n138), .A3(d1stg_inf_in1), .A4(
        n137), .A5(div_dz_out_in), .Y(n139) );
  AO22X1_RVT U267 ( .A1(\d2stg_opdec[2] ), .A2(n140), .A3(\d1stg_opdec[2] ), 
        .A4(n139), .Y(div_norm_inf) );
  AND2X1_RVT U268 ( .A1(div_expadd2_no_decr_load), .A2(n141), .Y(
        div_frac_add_in1_add) );
  NAND2X0_RVT U269 ( .A1(n142), .A2(n146), .Y(div_frac_add_in2_load) );
  OR2X1_RVT U270 ( .A1(div_frac_add_in1_add), .A2(div_frac_add_in2_load), .Y(
        div_frac_add_in1_load) );
  AO22X1_RVT U271 ( .A1(d6stg_fdivd), .A2(d6stg_frac_2), .A3(n143), .A4(
        d6stg_frac_31), .Y(d7stg_lsb_in) );
  AO22X1_RVT U272 ( .A1(d6stg_fdivd), .A2(d6stg_frac_1), .A3(n143), .A4(
        d6stg_frac_30), .Y(d7stg_grd_in) );
  AO221X1_RVT U273 ( .A1(d6stg_fdivd), .A2(d6stg_frac_0), .A3(n143), .A4(
        d6stg_frac_29), .A5(div_frac_add_in1_neq_0), .Y(d7stg_stk_in) );
  NAND4X0_RVT U274 ( .A1(n163), .A2(n146), .A3(n145), .A4(n144), .Y(
        div_frac_out_load) );
  NAND2X0_RVT U275 ( .A1(div_ctl_rst_l), .A2(d234stg_fdiv_in), .Y(n147) );
  OA221X1_RVT U276 ( .A1(n183), .A2(d1stg_dblopa[4]), .A3(n152), .A4(inq_op[1]), .A5(n147), .Y(div_expadd1_in1_dbl_in) );
  OA221X1_RVT U277 ( .A1(n183), .A2(d1stg_sngopa[4]), .A3(n152), .A4(inq_op[0]), .A5(n147), .Y(div_expadd1_in1_sng_in) );
  AND2X1_RVT U278 ( .A1(div_expadd1_in2_exp_in2_dbl), .A2(n153), .Y(
        div_exp1_0835) );
  AND2X1_RVT U279 ( .A1(div_expadd1_in2_exp_in2_sng), .A2(n153), .Y(
        div_exp1_0118) );
  AND2X1_RVT U280 ( .A1(\d5stg_opdec[2] ), .A2(n155), .Y(d6stg_opdec_in[2]) );
  OR2X1_RVT U281 ( .A1(d6stg_fdiv), .A2(d6stg_opdec_in[2]), .Y(
        div_expadd2_in1_exp_out_in) );
  AND3X1_RVT U282 ( .A1(d7stg_fdiv), .A2(n158), .A3(n157), .Y(
        div_exp_out_exp_out) );
  NAND2X0_RVT U283 ( .A1(div_exp_out[12]), .A2(d7stg_fdiv), .Y(n159) );
  AO22X1_RVT U284 ( .A1(div_exp_out_exp_out), .A2(n162), .A3(n161), .A4(n159), 
        .Y(div_exp_out_expadd2) );
  AND2X1_RVT U285 ( .A1(d7stg_fdiv), .A2(d7stg_in_of), .Y(div_frac_out_of) );
  NAND2X0_RVT U286 ( .A1(div_exp_out_expadd22_inv), .A2(n163), .Y(
        div_exp_out_load) );
  OA21X1_RVT U287 ( .A1(div_exp1[0]), .A2(d5stg_fdivs), .A3(div_exp1[4]), .Y(
        n172) );
  OA222X1_RVT U288 ( .A1(div_exp1[2]), .A2(d5stg_fdivs), .A3(n165), .A4(
        div_exp1[5]), .A5(n169), .A6(n164), .Y(n166) );
  OA221X1_RVT U289 ( .A1(div_exp1[3]), .A2(n169), .A3(n168), .A4(n167), .A5(
        n166), .Y(n171) );
  AND4X1_RVT U290 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .Y(n174) );
  NOR3X0_RVT U291 ( .A1(n174), .A2(div_frac_out_53), .A3(div_expadd2_12), .Y(
        n154) );
  OA22X1_RVT U292 ( .A1(div_exp_in1_exp_neq_ffs), .A2(div_exp_in2_exp_neq_ffs), 
        .A3(d1stg_dblopa[3]), .A4(d1stg_sngopa[3]), .Y(d1stg_infnan_in) );
  NOR2X0_RVT U293 ( .A1(d1stg_infnan_in), .A2(d1stg_zero_in), .Y(n149) );
endmodule


module clken_buf_5 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_2 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_2 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE11_1 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, net24264, n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE11_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24264), .TE(1'b0) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24264), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24264), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24264), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24264), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24264), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24264), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24264), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24264), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24264), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24264), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24264), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  OR2X1_RVT U15 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_2 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_2 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE13_1 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, net24246,
         n1, n2;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE13_1 clk_gate_q_reg ( .CLK(clk), .EN(n2), 
        .ENCLK(net24246), .TE(1'b0) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24246), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24246), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24246), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24246), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24246), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24246), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24246), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24246), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24246), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24246), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24246), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24246), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24246), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  AND2X1_RVT U15 ( .A1(din[12]), .A2(n1), .Y(N16) );
  OR2X1_RVT U17 ( .A1(se), .A2(en), .Y(n2) );
endmodule


module fpu_div_exp_dp ( inq_in1, inq_in2, d1stg_step, d234stg_fdiv, 
        div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl, 
        div_expadd1_in2_exp_in2_sng, d3stg_fdiv, d4stg_fdiv, div_shl_cnt, 
        div_exp1_expadd1, div_exp1_0835, div_exp1_0118, div_exp1_zero, 
        div_exp1_load, div_expadd2_in1_exp_out, d5stg_fdiva, d5stg_fdivd, 
        d5stg_fdivs, d6stg_fdiv, d7stg_fdiv, div_expadd2_no_decr_inv, 
        div_expadd2_cin, div_exp_out_expadd2, div_exp_out_expadd22_inv, 
        div_exp_out_of, d7stg_to_0_inv, d7stg_fdivd, div_exp_out_exp_out, 
        d7stg_rndup_inv, div_frac_add_52_inv, div_exp_out_load, fdiv_clken_l, 
        rclk, div_exp1, div_expadd2_12, div_exp_out, div_exp_outa, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [5:0] div_shl_cnt;
  output [12:0] div_exp1;
  output [12:0] div_exp_out;
  output [10:0] div_exp_outa;
  input d1stg_step, d234stg_fdiv, div_expadd1_in1_dbl, div_expadd1_in1_sng,
         div_expadd1_in2_exp_in2_dbl, div_expadd1_in2_exp_in2_sng, d3stg_fdiv,
         d4stg_fdiv, div_exp1_expadd1, div_exp1_0835, div_exp1_0118,
         div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out, d5stg_fdiva,
         d5stg_fdivd, d5stg_fdivs, d6stg_fdiv, d7stg_fdiv,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd2,
         div_exp_out_expadd22_inv, div_exp_out_of, d7stg_to_0_inv, d7stg_fdivd,
         div_exp_out_exp_out, d7stg_rndup_inv, div_frac_add_52_inv,
         div_exp_out_load, fdiv_clken_l, rclk, se, si;
  output div_expadd2_12, so;
  wire   clk, \intadd_8/A[8] , \intadd_8/A[7] , \intadd_8/A[6] ,
         \intadd_8/A[5] , \intadd_8/A[4] , \intadd_8/A[3] , \intadd_8/A[2] ,
         \intadd_8/A[1] , \intadd_8/A[0] , \intadd_8/B[8] , \intadd_8/B[7] ,
         \intadd_8/B[6] , \intadd_8/B[5] , \intadd_8/B[4] , \intadd_8/B[3] ,
         \intadd_8/B[2] , \intadd_8/B[1] , \intadd_8/B[0] , \intadd_8/CI ,
         \intadd_8/SUM[8] , \intadd_8/SUM[7] , \intadd_8/SUM[6] ,
         \intadd_8/SUM[5] , \intadd_8/SUM[4] , \intadd_8/SUM[3] ,
         \intadd_8/SUM[2] , \intadd_8/SUM[1] , \intadd_8/SUM[0] ,
         \intadd_8/n9 , \intadd_8/n8 , \intadd_8/n7 , \intadd_8/n6 ,
         \intadd_8/n5 , \intadd_8/n4 , \intadd_8/n3 , \intadd_8/n2 ,
         \intadd_8/n1 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136;
  wire   [10:0] div_exp_in1;
  wire   [10:0] div_exp_in2;
  wire   [12:0] div_exp1_in;
  wire   [12:0] div_exp_out_in;
  assign div_exp_outa[10] = div_exp_out[10];
  assign div_exp_outa[9] = div_exp_out[9];
  assign div_exp_outa[8] = div_exp_out[8];
  assign div_exp_outa[7] = div_exp_out[7];
  assign div_exp_outa[6] = div_exp_out[6];
  assign div_exp_outa[5] = div_exp_out[5];
  assign div_exp_outa[4] = div_exp_out[4];
  assign div_exp_outa[3] = div_exp_out[3];
  assign div_exp_outa[2] = div_exp_out[2];
  assign div_exp_outa[1] = div_exp_out[1];
  assign div_exp_outa[0] = div_exp_out[0];
  assign so = 1'b0;

  clken_buf_5 ckbuf_div_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fdiv_clken_l), 
        .tmb_l(n136) );
  dffe_SIZE11_2 i_div_exp_in1 ( .din(inq_in1), .en(d1stg_step), .clk(clk), .q(
        div_exp_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE11_1 i_div_exp_in2 ( .din(inq_in2), .en(d1stg_step), .clk(clk), .q(
        div_exp_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_2 i_div_exp1 ( .din(div_exp1_in), .en(div_exp1_load), .clk(clk), 
        .q(div_exp1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE13_1 i_div_exp_out ( .din(div_exp_out_in), .en(div_exp_out_load), 
        .clk(clk), .q(div_exp_out), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  FADDX1_RVT \intadd_8/U10  ( .A(\intadd_8/B[0] ), .B(\intadd_8/A[0] ), .CI(
        \intadd_8/CI ), .CO(\intadd_8/n9 ), .S(\intadd_8/SUM[0] ) );
  FADDX1_RVT \intadd_8/U9  ( .A(\intadd_8/B[1] ), .B(\intadd_8/A[1] ), .CI(
        \intadd_8/n9 ), .CO(\intadd_8/n8 ), .S(\intadd_8/SUM[1] ) );
  FADDX1_RVT \intadd_8/U8  ( .A(\intadd_8/B[2] ), .B(\intadd_8/A[2] ), .CI(
        \intadd_8/n8 ), .CO(\intadd_8/n7 ), .S(\intadd_8/SUM[2] ) );
  FADDX1_RVT \intadd_8/U7  ( .A(\intadd_8/B[3] ), .B(\intadd_8/A[3] ), .CI(
        \intadd_8/n7 ), .CO(\intadd_8/n6 ), .S(\intadd_8/SUM[3] ) );
  FADDX1_RVT \intadd_8/U6  ( .A(\intadd_8/B[4] ), .B(\intadd_8/A[4] ), .CI(
        \intadd_8/n6 ), .CO(\intadd_8/n5 ), .S(\intadd_8/SUM[4] ) );
  FADDX1_RVT \intadd_8/U5  ( .A(\intadd_8/B[5] ), .B(\intadd_8/A[5] ), .CI(
        \intadd_8/n5 ), .CO(\intadd_8/n4 ), .S(\intadd_8/SUM[5] ) );
  FADDX1_RVT \intadd_8/U4  ( .A(\intadd_8/B[6] ), .B(\intadd_8/A[6] ), .CI(
        \intadd_8/n4 ), .CO(\intadd_8/n3 ), .S(\intadd_8/SUM[6] ) );
  FADDX1_RVT \intadd_8/U3  ( .A(\intadd_8/B[7] ), .B(\intadd_8/A[7] ), .CI(
        \intadd_8/n3 ), .CO(\intadd_8/n2 ), .S(\intadd_8/SUM[7] ) );
  FADDX1_RVT \intadd_8/U2  ( .A(\intadd_8/B[8] ), .B(\intadd_8/A[8] ), .CI(
        \intadd_8/n2 ), .CO(\intadd_8/n1 ), .S(\intadd_8/SUM[8] ) );
  OR3X1_RVT U1 ( .A1(n97), .A2(n96), .A3(n39), .Y(n40) );
  INVX0_RVT U2 ( .A(n89), .Y(n92) );
  INVX0_RVT U3 ( .A(n77), .Y(n71) );
  INVX0_RVT U4 ( .A(n90), .Y(n91) );
  INVX0_RVT U5 ( .A(div_shl_cnt[4]), .Y(n44) );
  INVX0_RVT U6 ( .A(n98), .Y(n39) );
  INVX1_RVT U7 ( .A(se), .Y(n136) );
  NAND2X0_RVT U8 ( .A1(div_exp_out_expadd22_inv), .A2(div_frac_add_52_inv), 
        .Y(n1) );
  NAND2X0_RVT U9 ( .A1(div_exp_out_expadd2), .A2(n1), .Y(n125) );
  INVX1_RVT U10 ( .A(n125), .Y(n134) );
  INVX1_RVT U11 ( .A(d5stg_fdiva), .Y(n2) );
  NAND2X0_RVT U12 ( .A1(div_expadd2_no_decr_inv), .A2(d6stg_fdiv), .Y(n110) );
  NAND2X0_RVT U13 ( .A1(n2), .A2(n110), .Y(n98) );
  AND2X1_RVT U14 ( .A1(n134), .A2(n98), .Y(n102) );
  AND2X1_RVT U15 ( .A1(n134), .A2(n39), .Y(n101) );
  INVX1_RVT U16 ( .A(div_expadd2_cin), .Y(n131) );
  AOI22X1_RVT U17 ( .A1(d5stg_fdiva), .A2(div_exp1[0]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[0]), .Y(n130) );
  AOI22X1_RVT U18 ( .A1(d5stg_fdiva), .A2(d5stg_fdivs), .A3(
        div_expadd2_no_decr_inv), .A4(d6stg_fdiv), .Y(n129) );
  AOI22X1_RVT U19 ( .A1(d5stg_fdiva), .A2(div_exp1[1]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[1]), .Y(n6) );
  MUX41X1_RVT U20 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n7), .S1(
        n6), .Y(n3) );
  INVX1_RVT U21 ( .A(n3), .Y(n5) );
  INVX1_RVT U22 ( .A(div_exp_out_of), .Y(n127) );
  OA21X1_RVT U23 ( .A1(div_frac_add_52_inv), .A2(d7stg_rndup_inv), .A3(
        div_exp_out_exp_out), .Y(n133) );
  NAND2X0_RVT U24 ( .A1(n133), .A2(div_exp_out[1]), .Y(n4) );
  NAND3X0_RVT U25 ( .A1(n5), .A2(n127), .A3(n4), .Y(div_exp_out_in[1]) );
  AO22X1_RVT U26 ( .A1(d5stg_fdiva), .A2(div_exp1[4]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[4]), .Y(n109) );
  INVX1_RVT U27 ( .A(n109), .Y(n8) );
  AO222X1_RVT U28 ( .A1(n39), .A2(n7), .A3(n39), .A4(n6), .A5(n7), .A6(n6), 
        .Y(n122) );
  AOI22X1_RVT U29 ( .A1(d5stg_fdiva), .A2(div_exp1[2]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[2]), .Y(n121) );
  AOI22X1_RVT U30 ( .A1(d5stg_fdiva), .A2(div_exp1[3]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[3]), .Y(n116) );
  AOI22X1_RVT U31 ( .A1(d5stg_fdiva), .A2(d5stg_fdivd), .A3(
        div_expadd2_no_decr_inv), .A4(d6stg_fdiv), .Y(n115) );
  AO222X1_RVT U32 ( .A1(n8), .A2(n112), .A3(n8), .A4(n110), .A5(n112), .A6(
        n110), .Y(n105) );
  AOI22X1_RVT U33 ( .A1(d5stg_fdiva), .A2(div_exp1[5]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[5]), .Y(n104) );
  AO22X1_RVT U34 ( .A1(d5stg_fdiva), .A2(div_exp1[6]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[6]), .Y(n13) );
  MUX41X1_RVT U35 ( .A1(n101), .A3(n102), .A2(n102), .A4(n101), .S0(n12), .S1(
        n13), .Y(n9) );
  INVX1_RVT U36 ( .A(n9), .Y(n11) );
  NAND2X0_RVT U37 ( .A1(n133), .A2(div_exp_out[6]), .Y(n10) );
  NAND3X0_RVT U38 ( .A1(n11), .A2(n127), .A3(n10), .Y(div_exp_out_in[6]) );
  INVX1_RVT U39 ( .A(n12), .Y(n14) );
  AO222X1_RVT U40 ( .A1(n98), .A2(n14), .A3(n98), .A4(n13), .A5(n14), .A6(n13), 
        .Y(n19) );
  AO22X1_RVT U41 ( .A1(d5stg_fdiva), .A2(div_exp1[7]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[7]), .Y(n18) );
  MUX41X1_RVT U42 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n19), .S1(
        n18), .Y(n15) );
  INVX1_RVT U43 ( .A(n15), .Y(n17) );
  NAND2X0_RVT U44 ( .A1(n133), .A2(div_exp_out[7]), .Y(n16) );
  NAND3X0_RVT U45 ( .A1(n17), .A2(n127), .A3(n16), .Y(div_exp_out_in[7]) );
  AO222X1_RVT U46 ( .A1(n98), .A2(n19), .A3(n98), .A4(n18), .A5(n19), .A6(n18), 
        .Y(n24) );
  AO22X1_RVT U47 ( .A1(d5stg_fdiva), .A2(div_exp1[8]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[8]), .Y(n23) );
  MUX41X1_RVT U48 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n24), .S1(
        n23), .Y(n20) );
  INVX1_RVT U49 ( .A(n20), .Y(n22) );
  NAND2X0_RVT U50 ( .A1(div_exp_out_of), .A2(d7stg_fdivd), .Y(n32) );
  NAND2X0_RVT U51 ( .A1(n133), .A2(div_exp_out[8]), .Y(n21) );
  NAND3X0_RVT U52 ( .A1(n22), .A2(n32), .A3(n21), .Y(div_exp_out_in[8]) );
  AO222X1_RVT U53 ( .A1(n98), .A2(n24), .A3(n98), .A4(n23), .A5(n24), .A6(n23), 
        .Y(n29) );
  AO22X1_RVT U54 ( .A1(d5stg_fdiva), .A2(div_exp1[9]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[9]), .Y(n28) );
  MUX41X1_RVT U55 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n29), .S1(
        n28), .Y(n25) );
  INVX1_RVT U56 ( .A(n25), .Y(n27) );
  NAND2X0_RVT U57 ( .A1(n133), .A2(div_exp_out[9]), .Y(n26) );
  NAND3X0_RVT U58 ( .A1(n27), .A2(n32), .A3(n26), .Y(div_exp_out_in[9]) );
  AO222X1_RVT U59 ( .A1(n98), .A2(n29), .A3(n98), .A4(n28), .A5(n29), .A6(n28), 
        .Y(n97) );
  AO22X1_RVT U60 ( .A1(d5stg_fdiva), .A2(div_exp1[10]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[10]), .Y(n96) );
  MUX41X1_RVT U61 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n97), .S1(
        n96), .Y(n30) );
  INVX1_RVT U62 ( .A(n30), .Y(n33) );
  NAND2X0_RVT U63 ( .A1(n133), .A2(div_exp_out[10]), .Y(n31) );
  NAND3X0_RVT U64 ( .A1(n33), .A2(n32), .A3(n31), .Y(div_exp_out_in[10]) );
  INVX1_RVT U65 ( .A(div_exp1_0835), .Y(n81) );
  INVX1_RVT U66 ( .A(div_exp1_0118), .Y(n80) );
  INVX1_RVT U67 ( .A(\intadd_8/SUM[2] ), .Y(n34) );
  NAND2X0_RVT U68 ( .A1(div_exp1_expadd1), .A2(n34), .Y(n35) );
  NAND3X0_RVT U69 ( .A1(n81), .A2(n80), .A3(n35), .Y(div_exp1_in[4]) );
  INVX1_RVT U70 ( .A(div_expadd1_in1_dbl), .Y(n61) );
  INVX1_RVT U71 ( .A(div_expadd1_in2_exp_in2_sng), .Y(n70) );
  INVX1_RVT U72 ( .A(d3stg_fdiv), .Y(n69) );
  AND2X1_RVT U73 ( .A1(n70), .A2(n69), .Y(n66) );
  AND2X1_RVT U74 ( .A1(n61), .A2(n66), .Y(n38) );
  INVX1_RVT U75 ( .A(div_exp_in2[10]), .Y(n36) );
  NAND2X0_RVT U76 ( .A1(n36), .A2(div_expadd1_in2_exp_in2_dbl), .Y(n37) );
  AND2X1_RVT U77 ( .A1(n38), .A2(n37), .Y(\intadd_8/A[8] ) );
  AOI22X1_RVT U78 ( .A1(d5stg_fdiva), .A2(div_exp1[12]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[12]), .Y(n43) );
  NAND3X0_RVT U79 ( .A1(div_exp_out[11]), .A2(n97), .A3(n96), .Y(n41) );
  AO22X1_RVT U80 ( .A1(d5stg_fdiva), .A2(div_exp1[11]), .A3(
        div_expadd2_in1_exp_out), .A4(div_exp_out[11]), .Y(n99) );
  OA22X1_RVT U81 ( .A1(n98), .A2(n41), .A3(n99), .A4(n40), .Y(n42) );
  HADDX1_RVT U82 ( .A0(n43), .B0(n42), .SO(div_expadd2_12) );
  INVX1_RVT U83 ( .A(div_expadd1_in2_exp_in2_dbl), .Y(n68) );
  OA22X1_RVT U84 ( .A1(div_exp_in2[4]), .A2(n68), .A3(div_exp_in2[7]), .A4(n70), .Y(n46) );
  OAI22X1_RVT U85 ( .A1(n44), .A2(d4stg_fdiv), .A3(div_shl_cnt[4]), .A4(
        d3stg_fdiv), .Y(n45) );
  INVX1_RVT U86 ( .A(div_expadd1_in1_sng), .Y(n64) );
  AND4X1_RVT U87 ( .A1(n46), .A2(n45), .A3(n64), .A4(n61), .Y(\intadd_8/A[2] )
         );
  AOI222X1_RVT U88 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[7]), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[4]), .A5(d234stg_fdiv), .A6(
        div_exp1[4]), .Y(\intadd_8/B[2] ) );
  OA22X1_RVT U89 ( .A1(div_shl_cnt[0]), .A2(n69), .A3(div_exp_in2[3]), .A4(n70), .Y(n49) );
  NAND2X0_RVT U90 ( .A1(d4stg_fdiv), .A2(div_shl_cnt[0]), .Y(n48) );
  OR2X1_RVT U91 ( .A1(div_exp_in2[0]), .A2(n68), .Y(n47) );
  NAND4X0_RVT U92 ( .A1(n49), .A2(n48), .A3(n64), .A4(n47), .Y(n89) );
  AO222X1_RVT U93 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[3]), .A3(
        div_exp_in1[0]), .A4(div_expadd1_in1_dbl), .A5(d234stg_fdiv), .A6(
        div_exp1[0]), .Y(n90) );
  NAND2X0_RVT U94 ( .A1(n89), .A2(n90), .Y(n88) );
  INVX1_RVT U95 ( .A(n88), .Y(n84) );
  OA22X1_RVT U96 ( .A1(div_exp_in2[4]), .A2(n70), .A3(div_shl_cnt[1]), .A4(n69), .Y(n52) );
  NAND2X0_RVT U97 ( .A1(d4stg_fdiv), .A2(div_shl_cnt[1]), .Y(n51) );
  OR2X1_RVT U98 ( .A1(div_exp_in2[1]), .A2(n68), .Y(n50) );
  NAND4X0_RVT U99 ( .A1(n52), .A2(n61), .A3(n51), .A4(n50), .Y(n83) );
  AO222X1_RVT U100 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[4]), .A3(
        d234stg_fdiv), .A4(div_exp1[1]), .A5(div_expadd1_in1_dbl), .A6(
        div_exp_in1[1]), .Y(n85) );
  AOI222X1_RVT U101 ( .A1(n84), .A2(n83), .A3(n84), .A4(n85), .A5(n83), .A6(
        n85), .Y(\intadd_8/A[0] ) );
  OA22X1_RVT U102 ( .A1(div_exp_in2[5]), .A2(n70), .A3(div_shl_cnt[2]), .A4(
        n69), .Y(n55) );
  NAND2X0_RVT U103 ( .A1(d4stg_fdiv), .A2(div_shl_cnt[2]), .Y(n54) );
  OR2X1_RVT U104 ( .A1(div_exp_in2[2]), .A2(n68), .Y(n53) );
  AND4X1_RVT U105 ( .A1(n55), .A2(n61), .A3(n54), .A4(n53), .Y(\intadd_8/B[0] ) );
  AOI222X1_RVT U106 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[5]), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[2]), .A5(d234stg_fdiv), .A6(
        div_exp1[2]), .Y(\intadd_8/CI ) );
  OA22X1_RVT U107 ( .A1(div_exp_in2[6]), .A2(n70), .A3(div_shl_cnt[3]), .A4(
        n69), .Y(n58) );
  NAND2X0_RVT U108 ( .A1(d4stg_fdiv), .A2(div_shl_cnt[3]), .Y(n57) );
  OR2X1_RVT U109 ( .A1(div_exp_in2[3]), .A2(n68), .Y(n56) );
  AND4X1_RVT U110 ( .A1(n58), .A2(n64), .A3(n57), .A4(n56), .Y(\intadd_8/A[1] ) );
  AOI222X1_RVT U111 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[6]), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[3]), .A5(d234stg_fdiv), .A6(
        div_exp1[3]), .Y(\intadd_8/B[1] ) );
  AOI222X1_RVT U112 ( .A1(div_expadd1_in1_sng), .A2(div_exp_in1[8]), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[5]), .A5(d234stg_fdiv), .A6(
        div_exp1[5]), .Y(\intadd_8/A[3] ) );
  OA22X1_RVT U113 ( .A1(div_exp_in2[8]), .A2(n70), .A3(div_shl_cnt[5]), .A4(
        n69), .Y(n62) );
  NAND2X0_RVT U114 ( .A1(d4stg_fdiv), .A2(div_shl_cnt[5]), .Y(n60) );
  OR2X1_RVT U115 ( .A1(div_exp_in2[5]), .A2(n68), .Y(n59) );
  AND4X1_RVT U116 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .Y(\intadd_8/B[3] ) );
  OA22X1_RVT U117 ( .A1(div_exp_in2[6]), .A2(n68), .A3(div_exp_in2[9]), .A4(
        n70), .Y(n63) );
  AND2X1_RVT U118 ( .A1(n63), .A2(n69), .Y(\intadd_8/A[4] ) );
  AOI222X1_RVT U119 ( .A1(div_exp1[6]), .A2(d234stg_fdiv), .A3(
        div_expadd1_in1_sng), .A4(div_exp_in1[9]), .A5(div_expadd1_in1_dbl), 
        .A6(div_exp_in1[6]), .Y(\intadd_8/B[4] ) );
  OA22X1_RVT U120 ( .A1(div_exp_in2[7]), .A2(n68), .A3(div_exp_in2[10]), .A4(
        n70), .Y(n65) );
  AND3X1_RVT U121 ( .A1(n65), .A2(n69), .A3(n64), .Y(\intadd_8/A[5] ) );
  AOI222X1_RVT U122 ( .A1(div_exp1[7]), .A2(d234stg_fdiv), .A3(
        div_expadd1_in1_sng), .A4(div_exp_in1[10]), .A5(div_expadd1_in1_dbl), 
        .A6(div_exp_in1[7]), .Y(\intadd_8/B[5] ) );
  OA21X1_RVT U123 ( .A1(div_exp_in2[8]), .A2(n68), .A3(n66), .Y(
        \intadd_8/A[6] ) );
  AOI22X1_RVT U124 ( .A1(div_exp1[8]), .A2(d234stg_fdiv), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[8]), .Y(\intadd_8/B[6] ) );
  OA21X1_RVT U125 ( .A1(div_exp_in2[9]), .A2(n68), .A3(n66), .Y(
        \intadd_8/A[7] ) );
  AOI22X1_RVT U126 ( .A1(div_exp1[9]), .A2(d234stg_fdiv), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[9]), .Y(\intadd_8/B[7] ) );
  AOI22X1_RVT U128 ( .A1(div_exp1[10]), .A2(d234stg_fdiv), .A3(
        div_expadd1_in1_dbl), .A4(div_exp_in1[10]), .Y(\intadd_8/B[8] ) );
  NAND3X0_RVT U129 ( .A1(n70), .A2(n69), .A3(n68), .Y(n74) );
  NAND2X0_RVT U130 ( .A1(div_exp1[11]), .A2(d234stg_fdiv), .Y(n67) );
  NAND4X0_RVT U131 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .Y(n77) );
  NAND3X0_RVT U132 ( .A1(d234stg_fdiv), .A2(div_exp1[11]), .A3(n74), .Y(n76)
         );
  OA21X1_RVT U133 ( .A1(n71), .A2(\intadd_8/n1 ), .A3(n76), .Y(n73) );
  NAND2X0_RVT U134 ( .A1(d234stg_fdiv), .A2(div_exp1[12]), .Y(n72) );
  FADDX1_RVT U135 ( .A(n74), .B(n73), .CI(n72), .S(n75) );
  AND2X1_RVT U136 ( .A1(div_exp1_expadd1), .A2(n75), .Y(div_exp1_in[12]) );
  NAND2X0_RVT U137 ( .A1(n77), .A2(n76), .Y(n78) );
  HADDX1_RVT U138 ( .A0(\intadd_8/n1 ), .B0(n78), .SO(n79) );
  AO21X1_RVT U139 ( .A1(div_exp1_expadd1), .A2(n79), .A3(div_exp1_0835), .Y(
        div_exp1_in[11]) );
  INVX1_RVT U140 ( .A(div_exp1_expadd1), .Y(n82) );
  NOR2X0_RVT U141 ( .A1(\intadd_8/SUM[8] ), .A2(n82), .Y(div_exp1_in[10]) );
  NOR2X0_RVT U142 ( .A1(\intadd_8/SUM[7] ), .A2(n82), .Y(div_exp1_in[9]) );
  OAI21X1_RVT U143 ( .A1(\intadd_8/SUM[6] ), .A2(n82), .A3(n80), .Y(
        div_exp1_in[8]) );
  NOR2X0_RVT U144 ( .A1(\intadd_8/SUM[5] ), .A2(n82), .Y(div_exp1_in[7]) );
  NOR2X0_RVT U145 ( .A1(\intadd_8/SUM[4] ), .A2(n82), .Y(div_exp1_in[6]) );
  OAI21X1_RVT U146 ( .A1(\intadd_8/SUM[3] ), .A2(n82), .A3(n81), .Y(
        div_exp1_in[5]) );
  OAI21X1_RVT U147 ( .A1(\intadd_8/SUM[1] ), .A2(n82), .A3(n80), .Y(
        div_exp1_in[3]) );
  OAI21X1_RVT U148 ( .A1(\intadd_8/SUM[0] ), .A2(n82), .A3(n81), .Y(
        div_exp1_in[2]) );
  HADDX1_RVT U149 ( .A0(n84), .B0(n83), .SO(n86) );
  HADDX1_RVT U150 ( .A0(n86), .B0(n85), .SO(n87) );
  AND2X1_RVT U151 ( .A1(n87), .A2(div_exp1_expadd1), .Y(div_exp1_in[1]) );
  AND2X1_RVT U152 ( .A1(n88), .A2(div_exp1_expadd1), .Y(n94) );
  NAND2X0_RVT U153 ( .A1(n92), .A2(n91), .Y(n93) );
  AND2X1_RVT U154 ( .A1(n94), .A2(n93), .Y(n95) );
  OR2X1_RVT U155 ( .A1(div_exp1_0835), .A2(n95), .Y(div_exp1_in[0]) );
  AO22X1_RVT U156 ( .A1(n134), .A2(div_expadd2_12), .A3(n133), .A4(
        div_exp_out[12]), .Y(div_exp_out_in[12]) );
  AO222X1_RVT U157 ( .A1(n98), .A2(n97), .A3(n98), .A4(n96), .A5(n97), .A6(n96), .Y(n100) );
  MUX41X1_RVT U158 ( .A1(n102), .A3(n101), .A2(n101), .A4(n102), .S0(n100), 
        .S1(n99), .Y(n103) );
  AO21X1_RVT U159 ( .A1(div_exp_out[11]), .A2(n133), .A3(n103), .Y(
        div_exp_out_in[11]) );
  FADDX1_RVT U160 ( .A(n129), .B(n105), .CI(n104), .CO(n12), .S(n107) );
  INVX1_RVT U161 ( .A(n133), .Y(n124) );
  INVX1_RVT U162 ( .A(div_exp_out[5]), .Y(n106) );
  OA22X1_RVT U163 ( .A1(n107), .A2(n125), .A3(n124), .A4(n106), .Y(n108) );
  NAND2X0_RVT U164 ( .A1(n108), .A2(n127), .Y(div_exp_out_in[5]) );
  HADDX1_RVT U165 ( .A0(n110), .B0(n109), .SO(n111) );
  HADDX1_RVT U166 ( .A0(n112), .B0(n111), .SO(n113) );
  AO22X1_RVT U167 ( .A1(n134), .A2(n113), .A3(n133), .A4(div_exp_out[4]), .Y(
        n114) );
  OR2X1_RVT U168 ( .A1(div_exp_out_of), .A2(n114), .Y(div_exp_out_in[4]) );
  FADDX1_RVT U169 ( .A(n117), .B(n116), .CI(n115), .CO(n112), .S(n119) );
  INVX1_RVT U170 ( .A(div_exp_out[3]), .Y(n118) );
  OA22X1_RVT U171 ( .A1(n119), .A2(n125), .A3(n124), .A4(n118), .Y(n120) );
  NAND2X0_RVT U172 ( .A1(n120), .A2(n127), .Y(div_exp_out_in[3]) );
  FADDX1_RVT U173 ( .A(n129), .B(n122), .CI(n121), .CO(n117), .S(n126) );
  INVX1_RVT U174 ( .A(div_exp_out[2]), .Y(n123) );
  OA22X1_RVT U175 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .Y(n128) );
  NAND2X0_RVT U176 ( .A1(n128), .A2(n127), .Y(div_exp_out_in[2]) );
  FADDX1_RVT U177 ( .A(n131), .B(n130), .CI(n129), .CO(n7), .S(n132) );
  INVX1_RVT U178 ( .A(n132), .Y(n135) );
  AO222X1_RVT U179 ( .A1(n135), .A2(n134), .A3(div_exp_out_of), .A4(
        d7stg_to_0_inv), .A5(n133), .A6(div_exp_out[0]), .Y(div_exp_out_in[0])
         );
endmodule


module clken_buf_4 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N1, clken, n2;

  LATCHX1_RVT clken_reg ( .CLK(n2), .D(N1), .Q(clken) );
  NAND2X0_RVT U2 ( .A1(tmb_l), .A2(enb_l), .Y(N1) );
  AND2X1_RVT U3 ( .A1(rclk), .A2(clken), .Y(clk) );
  INVX0_RVT U4 ( .A(rclk), .Y(n2) );
endmodule


module fpu_cnt_lead0_lvl4_1 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX1_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_24_eq_0), .A2(n1), .Y(lead0_32b_3) );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl4_2 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_31_16_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_31_16_eq_0), .A2(din_15_0_eq_0), .Y(din_31_0_eq_0)
         );
  AO22X1_RVT U3 ( .A1(din_31_16_eq_0), .A2(din_15_8_eq_0), .A3(n1), .A4(
        din_31_24_eq_0), .Y(lead0_32b_3) );
  AO22X1_RVT U4 ( .A1(din_31_16_eq_0), .A2(lead0_16b_2_lo), .A3(n1), .A4(
        lead0_16b_2_hi), .Y(lead0_32b_2) );
  AO22X1_RVT U5 ( .A1(din_31_16_eq_0), .A2(lead0_16b_1_lo), .A3(n1), .A4(
        lead0_16b_1_hi), .Y(lead0_32b_1) );
  AO22X1_RVT U6 ( .A1(din_31_16_eq_0), .A2(lead0_16b_0_lo), .A3(n1), .A4(
        lead0_16b_0_hi), .Y(lead0_32b_0) );
endmodule


module fpu_cnt_lead0_lvl3_1 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_2 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl3_3 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_15_8_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_15_8_eq_0), .A2(din_7_0_eq_0), .Y(din_15_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_15_8_eq_0), .A2(din_7_4_eq_0), .A3(n1), .A4(
        din_15_12_eq_0), .Y(lead0_16b_2) );
  AO22X1_RVT U4 ( .A1(din_15_8_eq_0), .A2(lead0_8b_1_lo), .A3(n1), .A4(
        lead0_8b_1_hi), .Y(lead0_16b_1) );
  AO22X1_RVT U5 ( .A1(din_15_8_eq_0), .A2(lead0_8b_0_lo), .A3(n1), .A4(
        lead0_8b_0_hi), .Y(lead0_16b_0) );
endmodule


module fpu_cnt_lead0_lvl1_1 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_2 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_3 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_4 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_5 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_6 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_7 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_8 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_9 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_10 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_11 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_12 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl1_13 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din[2]), .Y(n1) );
  AOI21X1_RVT U2 ( .A1(din[1]), .A2(n1), .A3(din[3]), .Y(lead0_4b_0) );
  NOR4X1_RVT U3 ( .A1(din[3]), .A2(din[2]), .A3(din[1]), .A4(din[0]), .Y(
        din_3_0_eq_0) );
  NOR2X0_RVT U4 ( .A1(din[3]), .A2(din[2]), .Y(din_3_2_eq_0) );
endmodule


module fpu_cnt_lead0_lvl2_1 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_2 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_3 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_4 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_5 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_lvl2_6 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   n1;

  INVX0_RVT U1 ( .A(din_7_4_eq_0), .Y(n1) );
  AND2X1_RVT U2 ( .A1(din_7_4_eq_0), .A2(din_3_0_eq_0), .Y(din_7_0_eq_0) );
  AO22X1_RVT U3 ( .A1(din_7_4_eq_0), .A2(din_3_2_eq_0), .A3(n1), .A4(
        din_7_6_eq_0), .Y(lead0_8b_1) );
  AO22X1_RVT U4 ( .A1(din_7_4_eq_0), .A2(lead0_4b_0_lo), .A3(n1), .A4(
        lead0_4b_0_hi), .Y(lead0_8b_0) );
endmodule


module fpu_cnt_lead0_53b_1 ( din, lead0 );
  input [52:0] din;
  output [5:0] lead0;
  wire   din_52_49_eq_0, din_52_51_eq_0, lead0_52_49_0, din_48_45_eq_0,
         din_48_47_eq_0, lead0_48_45_0, din_44_41_eq_0, din_44_43_eq_0,
         lead0_44_41_0, din_40_37_eq_0, din_40_39_eq_0, lead0_40_37_0,
         din_36_33_eq_0, din_36_35_eq_0, lead0_36_33_0, din_32_29_eq_0,
         din_32_31_eq_0, lead0_32_29_0, din_28_25_eq_0, din_28_27_eq_0,
         lead0_28_25_0, din_24_21_eq_0, din_24_23_eq_0, lead0_24_21_0,
         din_20_17_eq_0, din_20_19_eq_0, lead0_20_17_0, din_16_13_eq_0,
         din_16_15_eq_0, lead0_16_13_0, din_12_9_eq_0, din_12_11_eq_0,
         lead0_12_9_0, din_8_5_eq_0, din_8_7_eq_0, lead0_8_5_0, din_4_1_eq_0,
         din_4_3_eq_0, lead0_4_1_0, din_52_45_eq_0, lead0_52_45_1,
         lead0_52_45_0, din_44_37_eq_0, lead0_44_37_1, lead0_44_37_0,
         din_36_29_eq_0, lead0_36_29_1, lead0_36_29_0, din_28_21_eq_0,
         lead0_28_21_1, lead0_28_21_0, din_20_13_eq_0, lead0_20_13_1,
         lead0_20_13_0, din_12_5_eq_0, lead0_12_5_1, lead0_12_5_0, lead0_4_0_1,
         lead0_4_0_0, din_52_37_eq_0, lead0_52_37_2, lead0_52_37_1,
         lead0_52_37_0, din_36_21_eq_0, lead0_36_21_2, lead0_36_21_1,
         lead0_36_21_0, din_20_5_eq_0, lead0_20_5_2, lead0_20_5_1,
         lead0_20_5_0, lead0_52_21_3, lead0_52_21_2, lead0_52_21_1,
         lead0_52_21_0, lead0_20_0_3, lead0_20_0_2, lead0_20_0_1, lead0_20_0_0,
         n1, n2, n3;

  fpu_cnt_lead0_lvl1_13 i_fpu_cnt_lead0_lvl1_52_49 ( .din(din[52:49]), 
        .din_3_0_eq_0(din_52_49_eq_0), .din_3_2_eq_0(din_52_51_eq_0), 
        .lead0_4b_0(lead0_52_49_0) );
  fpu_cnt_lead0_lvl1_12 i_fpu_cnt_lead0_lvl1_48_45 ( .din(din[48:45]), 
        .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(din_48_47_eq_0), 
        .lead0_4b_0(lead0_48_45_0) );
  fpu_cnt_lead0_lvl1_11 i_fpu_cnt_lead0_lvl1_44_41 ( .din(din[44:41]), 
        .din_3_0_eq_0(din_44_41_eq_0), .din_3_2_eq_0(din_44_43_eq_0), 
        .lead0_4b_0(lead0_44_41_0) );
  fpu_cnt_lead0_lvl1_10 i_fpu_cnt_lead0_lvl1_40_37 ( .din(din[40:37]), 
        .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(din_40_39_eq_0), 
        .lead0_4b_0(lead0_40_37_0) );
  fpu_cnt_lead0_lvl1_9 i_fpu_cnt_lead0_lvl1_36_33 ( .din(din[36:33]), 
        .din_3_0_eq_0(din_36_33_eq_0), .din_3_2_eq_0(din_36_35_eq_0), 
        .lead0_4b_0(lead0_36_33_0) );
  fpu_cnt_lead0_lvl1_8 i_fpu_cnt_lead0_lvl1_32_29 ( .din(din[32:29]), 
        .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(din_32_31_eq_0), 
        .lead0_4b_0(lead0_32_29_0) );
  fpu_cnt_lead0_lvl1_7 i_fpu_cnt_lead0_lvl1_28_25 ( .din(din[28:25]), 
        .din_3_0_eq_0(din_28_25_eq_0), .din_3_2_eq_0(din_28_27_eq_0), 
        .lead0_4b_0(lead0_28_25_0) );
  fpu_cnt_lead0_lvl1_6 i_fpu_cnt_lead0_lvl1_24_21 ( .din(din[24:21]), 
        .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(din_24_23_eq_0), 
        .lead0_4b_0(lead0_24_21_0) );
  fpu_cnt_lead0_lvl1_5 i_fpu_cnt_lead0_lvl1_20_17 ( .din(din[20:17]), 
        .din_3_0_eq_0(din_20_17_eq_0), .din_3_2_eq_0(din_20_19_eq_0), 
        .lead0_4b_0(lead0_20_17_0) );
  fpu_cnt_lead0_lvl1_4 i_fpu_cnt_lead0_lvl1_16_13 ( .din(din[16:13]), 
        .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(din_16_15_eq_0), 
        .lead0_4b_0(lead0_16_13_0) );
  fpu_cnt_lead0_lvl1_3 i_fpu_cnt_lead0_lvl1_12_9 ( .din(din[12:9]), 
        .din_3_0_eq_0(din_12_9_eq_0), .din_3_2_eq_0(din_12_11_eq_0), 
        .lead0_4b_0(lead0_12_9_0) );
  fpu_cnt_lead0_lvl1_2 i_fpu_cnt_lead0_lvl1_8_5 ( .din(din[8:5]), 
        .din_3_0_eq_0(din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0(
        lead0_8_5_0) );
  fpu_cnt_lead0_lvl1_1 i_fpu_cnt_lead0_lvl1_4_1 ( .din(din[4:1]), 
        .din_3_0_eq_0(din_4_1_eq_0), .din_3_2_eq_0(din_4_3_eq_0), .lead0_4b_0(
        lead0_4_1_0) );
  fpu_cnt_lead0_lvl2_6 i_fpu_cnt_lead0_lvl2_52_45 ( .din_7_4_eq_0(
        din_52_49_eq_0), .din_7_6_eq_0(din_52_51_eq_0), .lead0_4b_0_hi(
        lead0_52_49_0), .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(
        din_48_47_eq_0), .lead0_4b_0_lo(lead0_48_45_0), .din_7_0_eq_0(
        din_52_45_eq_0), .lead0_8b_1(lead0_52_45_1), .lead0_8b_0(lead0_52_45_0) );
  fpu_cnt_lead0_lvl2_5 i_fpu_cnt_lead0_lvl2_44_37 ( .din_7_4_eq_0(
        din_44_41_eq_0), .din_7_6_eq_0(din_44_43_eq_0), .lead0_4b_0_hi(
        lead0_44_41_0), .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(
        din_40_39_eq_0), .lead0_4b_0_lo(lead0_40_37_0), .din_7_0_eq_0(
        din_44_37_eq_0), .lead0_8b_1(lead0_44_37_1), .lead0_8b_0(lead0_44_37_0) );
  fpu_cnt_lead0_lvl2_4 i_fpu_cnt_lead0_lvl2_36_29 ( .din_7_4_eq_0(
        din_36_33_eq_0), .din_7_6_eq_0(din_36_35_eq_0), .lead0_4b_0_hi(
        lead0_36_33_0), .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(
        din_32_31_eq_0), .lead0_4b_0_lo(lead0_32_29_0), .din_7_0_eq_0(
        din_36_29_eq_0), .lead0_8b_1(lead0_36_29_1), .lead0_8b_0(lead0_36_29_0) );
  fpu_cnt_lead0_lvl2_3 i_fpu_cnt_lead0_lvl2_28_21 ( .din_7_4_eq_0(
        din_28_25_eq_0), .din_7_6_eq_0(din_28_27_eq_0), .lead0_4b_0_hi(
        lead0_28_25_0), .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(
        din_24_23_eq_0), .lead0_4b_0_lo(lead0_24_21_0), .din_7_0_eq_0(
        din_28_21_eq_0), .lead0_8b_1(lead0_28_21_1), .lead0_8b_0(lead0_28_21_0) );
  fpu_cnt_lead0_lvl2_2 i_fpu_cnt_lead0_lvl2_20_13 ( .din_7_4_eq_0(
        din_20_17_eq_0), .din_7_6_eq_0(din_20_19_eq_0), .lead0_4b_0_hi(
        lead0_20_17_0), .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(
        din_16_15_eq_0), .lead0_4b_0_lo(lead0_16_13_0), .din_7_0_eq_0(
        din_20_13_eq_0), .lead0_8b_1(lead0_20_13_1), .lead0_8b_0(lead0_20_13_0) );
  fpu_cnt_lead0_lvl2_1 i_fpu_cnt_lead0_lvl2_12_5 ( .din_7_4_eq_0(din_12_9_eq_0), .din_7_6_eq_0(din_12_11_eq_0), .lead0_4b_0_hi(lead0_12_9_0), .din_3_0_eq_0(
        din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0_lo(lead0_8_5_0), .din_7_0_eq_0(din_12_5_eq_0), .lead0_8b_1(lead0_12_5_1), .lead0_8b_0(
        lead0_12_5_0) );
  fpu_cnt_lead0_lvl3_3 i_fpu_cnt_lead0_lvl3_52_37 ( .din_15_8_eq_0(
        din_52_45_eq_0), .din_15_12_eq_0(din_52_49_eq_0), .lead0_8b_1_hi(
        lead0_52_45_1), .lead0_8b_0_hi(lead0_52_45_0), .din_7_0_eq_0(
        din_44_37_eq_0), .din_7_4_eq_0(din_44_41_eq_0), .lead0_8b_1_lo(
        lead0_44_37_1), .lead0_8b_0_lo(lead0_44_37_0), .din_15_0_eq_0(
        din_52_37_eq_0), .lead0_16b_2(lead0_52_37_2), .lead0_16b_1(
        lead0_52_37_1), .lead0_16b_0(lead0_52_37_0) );
  fpu_cnt_lead0_lvl3_2 i_fpu_cnt_lead0_lvl3_36_21 ( .din_15_8_eq_0(
        din_36_29_eq_0), .din_15_12_eq_0(din_36_33_eq_0), .lead0_8b_1_hi(
        lead0_36_29_1), .lead0_8b_0_hi(lead0_36_29_0), .din_7_0_eq_0(
        din_28_21_eq_0), .din_7_4_eq_0(din_28_25_eq_0), .lead0_8b_1_lo(
        lead0_28_21_1), .lead0_8b_0_lo(lead0_28_21_0), .din_15_0_eq_0(
        din_36_21_eq_0), .lead0_16b_2(lead0_36_21_2), .lead0_16b_1(
        lead0_36_21_1), .lead0_16b_0(lead0_36_21_0) );
  fpu_cnt_lead0_lvl3_1 i_fpu_cnt_lead0_lvl3_20_5 ( .din_15_8_eq_0(
        din_20_13_eq_0), .din_15_12_eq_0(din_20_17_eq_0), .lead0_8b_1_hi(
        lead0_20_13_1), .lead0_8b_0_hi(lead0_20_13_0), .din_7_0_eq_0(
        din_12_5_eq_0), .din_7_4_eq_0(din_12_9_eq_0), .lead0_8b_1_lo(
        lead0_12_5_1), .lead0_8b_0_lo(lead0_12_5_0), .din_15_0_eq_0(
        din_20_5_eq_0), .lead0_16b_2(lead0_20_5_2), .lead0_16b_1(lead0_20_5_1), 
        .lead0_16b_0(lead0_20_5_0) );
  fpu_cnt_lead0_lvl4_2 i_fpu_cnt_lead0_lvl4_52_21 ( .din_31_16_eq_0(
        din_52_37_eq_0), .din_31_24_eq_0(din_52_45_eq_0), .lead0_16b_2_hi(
        lead0_52_37_2), .lead0_16b_1_hi(lead0_52_37_1), .lead0_16b_0_hi(
        lead0_52_37_0), .din_15_0_eq_0(din_36_21_eq_0), .din_15_8_eq_0(
        din_36_29_eq_0), .lead0_16b_2_lo(lead0_36_21_2), .lead0_16b_1_lo(
        lead0_36_21_1), .lead0_16b_0_lo(lead0_36_21_0), .din_31_0_eq_0(
        lead0[5]), .lead0_32b_3(lead0_52_21_3), .lead0_32b_2(lead0_52_21_2), 
        .lead0_32b_1(lead0_52_21_1), .lead0_32b_0(lead0_52_21_0) );
  fpu_cnt_lead0_lvl4_1 i_fpu_cnt_lead0_lvl4_20_0 ( .din_31_16_eq_0(
        din_20_5_eq_0), .din_31_24_eq_0(din_20_13_eq_0), .lead0_16b_2_hi(
        lead0_20_5_2), .lead0_16b_1_hi(lead0_20_5_1), .lead0_16b_0_hi(
        lead0_20_5_0), .din_15_0_eq_0(1'b0), .din_15_8_eq_0(1'b0), 
        .lead0_16b_2_lo(din_4_1_eq_0), .lead0_16b_1_lo(lead0_4_0_1), 
        .lead0_16b_0_lo(lead0_4_0_0), .lead0_32b_3(lead0_20_0_3), 
        .lead0_32b_2(lead0_20_0_2), .lead0_32b_1(lead0_20_0_1), .lead0_32b_0(
        lead0_20_0_0) );
  INVX0_RVT U2 ( .A(din[0]), .Y(n2) );
  INVX1_RVT U4 ( .A(din_4_1_eq_0), .Y(n1) );
  AND2X1_RVT U5 ( .A1(din_4_3_eq_0), .A2(n1), .Y(lead0_4_0_1) );
  AO22X1_RVT U6 ( .A1(din_4_1_eq_0), .A2(n2), .A3(n1), .A4(lead0_4_1_0), .Y(
        lead0_4_0_0) );
  INVX1_RVT U7 ( .A(lead0[5]), .Y(n3) );
  AO22X1_RVT U8 ( .A1(lead0[5]), .A2(din_20_5_eq_0), .A3(n3), .A4(
        din_52_37_eq_0), .Y(lead0[4]) );
  AO22X1_RVT U9 ( .A1(lead0[5]), .A2(lead0_20_0_3), .A3(n3), .A4(lead0_52_21_3), .Y(lead0[3]) );
  AO22X1_RVT U10 ( .A1(lead0[5]), .A2(lead0_20_0_2), .A3(n3), .A4(
        lead0_52_21_2), .Y(lead0[2]) );
  AO22X1_RVT U11 ( .A1(lead0[5]), .A2(lead0_20_0_1), .A3(n3), .A4(
        lead0_52_21_1), .Y(lead0[1]) );
  AO22X1_RVT U12 ( .A1(lead0[5]), .A2(lead0_20_0_0), .A3(n3), .A4(
        lead0_52_21_0), .Y(lead0[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_7 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_7 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n5), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n5), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n5), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n5), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n5), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n5), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_6 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_6 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n5), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n5), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n5), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n5), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n5), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n5), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module dff_SIZE53_0 ( din, clk, se, si, so, \q[52]_BAR , \q[51]_BAR , 
        \q[50]_BAR , \q[49]_BAR , \q[48]_BAR , \q[47]_BAR , \q[46]_BAR , 
        \q[45]_BAR , \q[44]_BAR , \q[43]_BAR , \q[42]_BAR , \q[41]_BAR , 
        \q[40]_BAR , \q[39]_BAR , \q[38]_BAR , \q[37]_BAR , \q[36]_BAR , 
        \q[35]_BAR , \q[34]_BAR , \q[33]_BAR , \q[32]_BAR , \q[31]_BAR , 
        \q[30]_BAR , \q[29]_BAR , \q[28]_BAR , \q[27]_BAR , \q[26]_BAR , 
        \q[25]_BAR , \q[24]_BAR , \q[23]_BAR , \q[22]_BAR , \q[21]_BAR , 
        \q[20]_BAR , \q[19]_BAR , \q[18]_BAR , \q[17]_BAR , \q[16]_BAR , 
        \q[15]_BAR , \q[14]_BAR , \q[13]_BAR , \q[12]_BAR , \q[11]_BAR , 
        \q[10]_BAR , \q[9]_BAR , \q[8]_BAR , \q[7]_BAR , \q[6]_BAR , 
        \q[5]_BAR , \q[4]_BAR , \q[3]_BAR , \q[2]_BAR , \q[1]_BAR , \q[0]_BAR 
 );
  input [52:0] din;
  input [52:0] si;
  output [52:0] so;
  input clk, se;
  output \q[52]_BAR , \q[51]_BAR , \q[50]_BAR , \q[49]_BAR , \q[48]_BAR ,
         \q[47]_BAR , \q[46]_BAR , \q[45]_BAR , \q[44]_BAR , \q[43]_BAR ,
         \q[42]_BAR , \q[41]_BAR , \q[40]_BAR , \q[39]_BAR , \q[38]_BAR ,
         \q[37]_BAR , \q[36]_BAR , \q[35]_BAR , \q[34]_BAR , \q[33]_BAR ,
         \q[32]_BAR , \q[31]_BAR , \q[30]_BAR , \q[29]_BAR , \q[28]_BAR ,
         \q[27]_BAR , \q[26]_BAR , \q[25]_BAR , \q[24]_BAR , \q[23]_BAR ,
         \q[22]_BAR , \q[21]_BAR , \q[20]_BAR , \q[19]_BAR , \q[18]_BAR ,
         \q[17]_BAR , \q[16]_BAR , \q[15]_BAR , \q[14]_BAR , \q[13]_BAR ,
         \q[12]_BAR , \q[11]_BAR , \q[10]_BAR , \q[9]_BAR , \q[8]_BAR ,
         \q[7]_BAR , \q[6]_BAR , \q[5]_BAR , \q[4]_BAR , \q[3]_BAR ,
         \q[2]_BAR , \q[1]_BAR , \q[0]_BAR ;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N54, N55, n1, n2, n3;

  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .QN(\q[52]_BAR ) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .QN(\q[51]_BAR ) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .QN(\q[45]_BAR ) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .QN(\q[44]_BAR ) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .QN(\q[43]_BAR ) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .QN(\q[42]_BAR ) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .QN(\q[41]_BAR ) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .QN(\q[40]_BAR ) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .QN(\q[39]_BAR ) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .QN(\q[38]_BAR ) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .QN(\q[37]_BAR ) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .QN(\q[36]_BAR ) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .QN(\q[35]_BAR ) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .QN(\q[34]_BAR ) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .QN(\q[32]_BAR ) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .QN(\q[31]_BAR ) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .QN(\q[30]_BAR ) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .QN(\q[29]_BAR ) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .QN(\q[28]_BAR ) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .QN(\q[27]_BAR ) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .QN(\q[26]_BAR ) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .QN(\q[25]_BAR ) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .QN(\q[24]_BAR ) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .QN(\q[23]_BAR ) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .QN(\q[22]_BAR ) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .QN(\q[21]_BAR ) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .QN(\q[20]_BAR ) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .QN(\q[19]_BAR ) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .QN(\q[18]_BAR ) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .QN(\q[17]_BAR ) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .QN(\q[16]_BAR ) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .QN(\q[15]_BAR ) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .QN(\q[14]_BAR ) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .QN(\q[13]_BAR ) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .QN(\q[12]_BAR ) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .QN(\q[11]_BAR ) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .QN(\q[10]_BAR ) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .QN(\q[9]_BAR ) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .QN(\q[8]_BAR ) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .QN(\q[7]_BAR ) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .QN(\q[6]_BAR ) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .QN(\q[5]_BAR ) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .QN(\q[4]_BAR ) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .QN(\q[3]_BAR ) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .QN(\q[2]_BAR ) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .QN(\q[1]_BAR ) );
  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\q[0]_BAR ) );
  DFFSSRX1_RVT \q_reg[33]  ( .D(1'b0), .SETB(se), .RSTB(din[33]), .CLK(clk), 
        .QN(\q[33]_BAR ) );
  DFFSSRX1_RVT \q_reg[50]  ( .D(1'b0), .SETB(se), .RSTB(din[50]), .CLK(clk), 
        .QN(\q[50]_BAR ) );
  DFFSSRX1_RVT \q_reg[49]  ( .D(1'b0), .SETB(se), .RSTB(din[49]), .CLK(clk), 
        .QN(\q[49]_BAR ) );
  DFFSSRX1_RVT \q_reg[48]  ( .D(1'b0), .SETB(se), .RSTB(din[48]), .CLK(clk), 
        .QN(\q[48]_BAR ) );
  DFFSSRX1_RVT \q_reg[47]  ( .D(1'b0), .SETB(se), .RSTB(din[47]), .CLK(clk), 
        .QN(\q[47]_BAR ) );
  DFFSSRX1_RVT \q_reg[46]  ( .D(1'b0), .SETB(se), .RSTB(din[46]), .CLK(clk), 
        .QN(\q[46]_BAR ) );
  INVX1_RVT U10 ( .A(se), .Y(n1) );
  AND2X1_RVT U11 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U12 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U13 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U14 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U15 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U16 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U17 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U18 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U19 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U20 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U21 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U22 ( .A(se), .Y(n2) );
  AND2X1_RVT U23 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U24 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U25 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U26 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U27 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U28 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U29 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U30 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U31 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U32 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U33 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U34 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U35 ( .A(se), .Y(n3) );
  AND2X1_RVT U36 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U37 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U38 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U39 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U40 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U41 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U42 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U43 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U44 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U45 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U46 ( .A1(din[35]), .A2(n3), .Y(N38) );
  AND2X1_RVT U47 ( .A1(din[36]), .A2(n3), .Y(N39) );
  AND2X1_RVT U48 ( .A1(din[37]), .A2(n1), .Y(N40) );
  AND2X1_RVT U49 ( .A1(din[38]), .A2(n2), .Y(N41) );
  AND2X1_RVT U50 ( .A1(din[39]), .A2(n3), .Y(N42) );
  AND2X1_RVT U51 ( .A1(din[40]), .A2(n1), .Y(N43) );
  AND2X1_RVT U52 ( .A1(din[41]), .A2(n2), .Y(N44) );
  AND2X1_RVT U53 ( .A1(din[42]), .A2(n3), .Y(N45) );
  AND2X1_RVT U54 ( .A1(din[43]), .A2(n1), .Y(N46) );
  AND2X1_RVT U55 ( .A1(din[44]), .A2(n2), .Y(N47) );
  AND2X1_RVT U56 ( .A1(din[45]), .A2(n3), .Y(N48) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n1), .Y(N54) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N55) );
endmodule


module dff_SIZE12 ( din, clk, q, se, si, so );
  input [11:0] din;
  output [11:0] q;
  input [11:0] si;
  output [11:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, n1;
  assign q[5] = q[11];
  assign q[4] = q[10];
  assign q[3] = q[9];
  assign q[1] = q[7];
  assign q[0] = q[6];
  assign q[8] = q[2];

  DFFX1_RVT \q_reg[11]  ( .D(N8), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N7), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N6), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[7]  ( .D(N4), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N3), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
endmodule


module dff_SIZE53_1 ( din, clk, q, se, si, so );
  input [52:0] din;
  output [52:0] q;
  input [52:0] si;
  output [52:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, n1, n2, n3, n4;

  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  AND2X1_RVT U55 ( .A1(din[48]), .A2(n4), .Y(N51) );
  AND2X1_RVT U56 ( .A1(din[49]), .A2(n4), .Y(N52) );
  AND2X1_RVT U57 ( .A1(din[50]), .A2(n4), .Y(N53) );
  AND2X1_RVT U58 ( .A1(din[51]), .A2(n4), .Y(N54) );
  AND2X1_RVT U59 ( .A1(din[52]), .A2(n4), .Y(N55) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_5 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, net24228, n1, n2,
         n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_5 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  OR2X1_RVT U60 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_4 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, net24228, n1,
         n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_4 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  OR2X1_RVT U61 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_3 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_3 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_2 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_2 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n5), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n5), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n5), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n5), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n5), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n5), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module dffe_SIZE55_1 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, net24228,
         n1, n2, n4, n5, n6;

  SNPS_CLOCK_GATE_HIGH_dffe_SIZE55_1 clk_gate_q_reg ( .CLK(clk), .EN(n6), 
        .ENCLK(net24228), .TE(1'b0) );
  DFFX1_RVT \q_reg[54]  ( .D(N58), .CLK(net24228), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N57), .CLK(net24228), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N56), .CLK(net24228), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N55), .CLK(net24228), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N54), .CLK(net24228), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N53), .CLK(net24228), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N52), .CLK(net24228), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N51), .CLK(net24228), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N50), .CLK(net24228), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N49), .CLK(net24228), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N48), .CLK(net24228), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N47), .CLK(net24228), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N46), .CLK(net24228), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N45), .CLK(net24228), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N44), .CLK(net24228), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N43), .CLK(net24228), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N42), .CLK(net24228), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N41), .CLK(net24228), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N40), .CLK(net24228), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N39), .CLK(net24228), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N38), .CLK(net24228), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N37), .CLK(net24228), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N36), .CLK(net24228), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N35), .CLK(net24228), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N34), .CLK(net24228), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N33), .CLK(net24228), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N32), .CLK(net24228), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N31), .CLK(net24228), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N30), .CLK(net24228), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N29), .CLK(net24228), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N28), .CLK(net24228), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N27), .CLK(net24228), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N26), .CLK(net24228), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N25), .CLK(net24228), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N24), .CLK(net24228), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N23), .CLK(net24228), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N22), .CLK(net24228), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N21), .CLK(net24228), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N20), .CLK(net24228), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N19), .CLK(net24228), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N18), .CLK(net24228), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N17), .CLK(net24228), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N16), .CLK(net24228), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N15), .CLK(net24228), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N14), .CLK(net24228), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N13), .CLK(net24228), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N12), .CLK(net24228), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N11), .CLK(net24228), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N10), .CLK(net24228), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N9), .CLK(net24228), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N8), .CLK(net24228), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N7), .CLK(net24228), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N6), .CLK(net24228), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N5), .CLK(net24228), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N4), .CLK(net24228), .Q(q[0]) );
  INVX1_RVT U2 ( .A(se), .Y(n1) );
  AND2X1_RVT U3 ( .A1(din[0]), .A2(n1), .Y(N4) );
  AND2X1_RVT U4 ( .A1(din[1]), .A2(n1), .Y(N5) );
  AND2X1_RVT U5 ( .A1(din[2]), .A2(n1), .Y(N6) );
  AND2X1_RVT U6 ( .A1(din[3]), .A2(n1), .Y(N7) );
  AND2X1_RVT U7 ( .A1(din[4]), .A2(n1), .Y(N8) );
  AND2X1_RVT U8 ( .A1(din[5]), .A2(n1), .Y(N9) );
  AND2X1_RVT U9 ( .A1(din[6]), .A2(n1), .Y(N10) );
  AND2X1_RVT U10 ( .A1(din[7]), .A2(n1), .Y(N11) );
  AND2X1_RVT U11 ( .A1(din[8]), .A2(n1), .Y(N12) );
  AND2X1_RVT U12 ( .A1(din[9]), .A2(n1), .Y(N13) );
  AND2X1_RVT U13 ( .A1(din[10]), .A2(n1), .Y(N14) );
  AND2X1_RVT U14 ( .A1(din[11]), .A2(n1), .Y(N15) );
  INVX1_RVT U15 ( .A(se), .Y(n2) );
  AND2X1_RVT U16 ( .A1(din[12]), .A2(n2), .Y(N16) );
  AND2X1_RVT U17 ( .A1(din[13]), .A2(n2), .Y(N17) );
  AND2X1_RVT U18 ( .A1(din[14]), .A2(n2), .Y(N18) );
  AND2X1_RVT U19 ( .A1(din[15]), .A2(n2), .Y(N19) );
  AND2X1_RVT U20 ( .A1(din[16]), .A2(n2), .Y(N20) );
  AND2X1_RVT U21 ( .A1(din[17]), .A2(n2), .Y(N21) );
  AND2X1_RVT U22 ( .A1(din[18]), .A2(n2), .Y(N22) );
  AND2X1_RVT U23 ( .A1(din[19]), .A2(n2), .Y(N23) );
  AND2X1_RVT U24 ( .A1(din[20]), .A2(n2), .Y(N24) );
  AND2X1_RVT U25 ( .A1(din[21]), .A2(n2), .Y(N25) );
  AND2X1_RVT U26 ( .A1(din[22]), .A2(n2), .Y(N26) );
  AND2X1_RVT U27 ( .A1(din[23]), .A2(n2), .Y(N27) );
  INVX1_RVT U28 ( .A(se), .Y(n4) );
  AND2X1_RVT U29 ( .A1(din[24]), .A2(n4), .Y(N28) );
  AND2X1_RVT U30 ( .A1(din[25]), .A2(n4), .Y(N29) );
  AND2X1_RVT U31 ( .A1(din[26]), .A2(n4), .Y(N30) );
  AND2X1_RVT U32 ( .A1(din[27]), .A2(n4), .Y(N31) );
  AND2X1_RVT U33 ( .A1(din[28]), .A2(n4), .Y(N32) );
  AND2X1_RVT U34 ( .A1(din[29]), .A2(n4), .Y(N33) );
  AND2X1_RVT U35 ( .A1(din[30]), .A2(n4), .Y(N34) );
  AND2X1_RVT U36 ( .A1(din[31]), .A2(n4), .Y(N35) );
  AND2X1_RVT U37 ( .A1(din[32]), .A2(n4), .Y(N36) );
  AND2X1_RVT U38 ( .A1(din[33]), .A2(n4), .Y(N37) );
  AND2X1_RVT U39 ( .A1(din[34]), .A2(n4), .Y(N38) );
  AND2X1_RVT U40 ( .A1(din[35]), .A2(n4), .Y(N39) );
  INVX1_RVT U41 ( .A(se), .Y(n5) );
  AND2X1_RVT U42 ( .A1(din[36]), .A2(n5), .Y(N40) );
  AND2X1_RVT U43 ( .A1(din[37]), .A2(n5), .Y(N41) );
  AND2X1_RVT U44 ( .A1(din[38]), .A2(n5), .Y(N42) );
  AND2X1_RVT U45 ( .A1(din[39]), .A2(n5), .Y(N43) );
  AND2X1_RVT U46 ( .A1(din[40]), .A2(n5), .Y(N44) );
  AND2X1_RVT U47 ( .A1(din[41]), .A2(n5), .Y(N45) );
  AND2X1_RVT U48 ( .A1(din[42]), .A2(n5), .Y(N46) );
  AND2X1_RVT U49 ( .A1(din[43]), .A2(n5), .Y(N47) );
  AND2X1_RVT U50 ( .A1(din[44]), .A2(n5), .Y(N48) );
  AND2X1_RVT U51 ( .A1(din[45]), .A2(n5), .Y(N49) );
  AND2X1_RVT U52 ( .A1(din[46]), .A2(n5), .Y(N50) );
  AND2X1_RVT U53 ( .A1(din[47]), .A2(n5), .Y(N51) );
  AND2X1_RVT U54 ( .A1(din[48]), .A2(n1), .Y(N52) );
  AND2X1_RVT U55 ( .A1(din[49]), .A2(n2), .Y(N53) );
  AND2X1_RVT U56 ( .A1(din[50]), .A2(n4), .Y(N54) );
  AND2X1_RVT U57 ( .A1(din[51]), .A2(n5), .Y(N55) );
  AND2X1_RVT U58 ( .A1(din[52]), .A2(n1), .Y(N56) );
  AND2X1_RVT U59 ( .A1(din[53]), .A2(n2), .Y(N57) );
  AND2X1_RVT U60 ( .A1(din[54]), .A2(n4), .Y(N58) );
  OR2X1_RVT U62 ( .A1(se), .A2(en), .Y(n6) );
endmodule


module fpu_div_frac_dp ( inq_in1, inq_in2, d1stg_step, 
        div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm, 
        div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm, 
        div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm, 
        div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf, 
        div_norm_qnan, d1stg_dblop, div_norm_zero, d1stg_snan_dbl_in1, 
        d1stg_snan_sng_in1, d1stg_snan_dbl_in2, d1stg_snan_sng_in2, d3stg_fdiv, 
        d6stg_fdiv, d6stg_fdivd, d6stg_fdivs, div_frac_add_in2_load, 
        d6stg_frac_out_shl1, d6stg_frac_out_nosh, d4stg_fdiv, 
        div_frac_add_in1_add, div_frac_add_in1_load, d5stg_fdivb, 
        div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl, 
        div_frac_out_shl1_sng, div_frac_out_of, d7stg_to_0, div_frac_out_load, 
        fdiv_clken_l, rclk, div_shl_cnt, d6stg_frac_0, d6stg_frac_1, 
        d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, d6stg_frac_31, 
        div_frac_add_in1_neq_0, div_frac_add_52_inv, div_frac_add_52_inva, 
        div_frac_out_54_53, div_frac_outa, se, si, so );
  input [54:0] inq_in1;
  input [54:0] inq_in2;
  output [5:0] div_shl_cnt;
  output [1:0] div_frac_out_54_53;
  output [51:0] div_frac_outa;
  input d1stg_step, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm,
         div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm,
         div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm,
         div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf,
         div_norm_qnan, d1stg_dblop, div_norm_zero, d1stg_snan_dbl_in1,
         d1stg_snan_sng_in1, d1stg_snan_dbl_in2, d1stg_snan_sng_in2,
         d3stg_fdiv, d6stg_fdiv, d6stg_fdivd, d6stg_fdivs,
         div_frac_add_in2_load, d6stg_frac_out_shl1, d6stg_frac_out_nosh,
         d4stg_fdiv, div_frac_add_in1_add, div_frac_add_in1_load, d5stg_fdivb,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, d7stg_to_0, div_frac_out_load,
         fdiv_clken_l, rclk, se, si;
  output d6stg_frac_0, d6stg_frac_1, d6stg_frac_2, d6stg_frac_29,
         d6stg_frac_30, d6stg_frac_31, div_frac_add_in1_neq_0,
         div_frac_add_52_inv, div_frac_add_52_inva, so;
  wire   clk, \div_frac_out[52] , n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, div_frac_add_52_inva, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1028;
  wire   [54:0] div_frac_in1;
  wire   [54:0] div_frac_in2;
  wire   [52:0] div_norm_inv;
  wire   [5:0] div_lead0;
  wire   [5:0] div_shl_cnta;
  wire   [52:0] div_shl_data;
  wire   [105:53] div_shl_tmp;
  wire   [54:0] div_shl_save;
  wire   [52:0] div_frac_add_in2_in;
  wire   [54:0] div_frac_add_in2;
  wire   [54:0] div_frac_add_in1;
  wire   [54:0] div_frac_add_in1_in;
  wire   [54:0] div_frac_add_in1a;
  wire   [54:0] div_frac_out_in;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign so = 1'b0;
  assign div_frac_add_52_inv = div_frac_add_52_inva;

  clken_buf_4 ckbuf_div_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fdiv_clken_l), 
        .tmb_l(n1028) );
  dffe_SIZE55_7 i_div_frac_in1 ( .din(inq_in1), .en(d1stg_step), .clk(clk), 
        .q(div_frac_in1), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE55_6 i_div_frac_in2 ( .din(inq_in2), .en(d1stg_step), .clk(clk), 
        .q(div_frac_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dff_SIZE53_0 i_div_norm_inv ( .din({n703, n702, n701, n700, n699, n698, n697, 
        n696, n695, n694, n693, n692, n691, n690, n689, n688, n687, n686, n685, 
        n684, n683, n682, n681, n680, n679, n678, n677, n676, n675, n674, n673, 
        n672, n671, n670, n669, n668, n667, n666, n665, n664, n663, n662, n661, 
        n660, n659, n658, n657, n656, n655, n654, n653, n652, n651}), .clk(clk), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\q[52]_BAR (
        div_norm_inv[52]), .\q[51]_BAR (div_norm_inv[51]), .\q[50]_BAR (
        div_norm_inv[50]), .\q[49]_BAR (div_norm_inv[49]), .\q[48]_BAR (
        div_norm_inv[48]), .\q[47]_BAR (div_norm_inv[47]), .\q[46]_BAR (
        div_norm_inv[46]), .\q[45]_BAR (div_norm_inv[45]), .\q[44]_BAR (
        div_norm_inv[44]), .\q[43]_BAR (div_norm_inv[43]), .\q[42]_BAR (
        div_norm_inv[42]), .\q[41]_BAR (div_norm_inv[41]), .\q[40]_BAR (
        div_norm_inv[40]), .\q[39]_BAR (div_norm_inv[39]), .\q[38]_BAR (
        div_norm_inv[38]), .\q[37]_BAR (div_norm_inv[37]), .\q[36]_BAR (
        div_norm_inv[36]), .\q[35]_BAR (div_norm_inv[35]), .\q[34]_BAR (
        div_norm_inv[34]), .\q[33]_BAR (div_norm_inv[33]), .\q[32]_BAR (
        div_norm_inv[32]), .\q[31]_BAR (div_norm_inv[31]), .\q[30]_BAR (
        div_norm_inv[30]), .\q[29]_BAR (div_norm_inv[29]), .\q[28]_BAR (
        div_norm_inv[28]), .\q[27]_BAR (div_norm_inv[27]), .\q[26]_BAR (
        div_norm_inv[26]), .\q[25]_BAR (div_norm_inv[25]), .\q[24]_BAR (
        div_norm_inv[24]), .\q[23]_BAR (div_norm_inv[23]), .\q[22]_BAR (
        div_norm_inv[22]), .\q[21]_BAR (div_norm_inv[21]), .\q[20]_BAR (
        div_norm_inv[20]), .\q[19]_BAR (div_norm_inv[19]), .\q[18]_BAR (
        div_norm_inv[18]), .\q[17]_BAR (div_norm_inv[17]), .\q[16]_BAR (
        div_norm_inv[16]), .\q[15]_BAR (div_norm_inv[15]), .\q[14]_BAR (
        div_norm_inv[14]), .\q[13]_BAR (div_norm_inv[13]), .\q[12]_BAR (
        div_norm_inv[12]), .\q[11]_BAR (div_norm_inv[11]), .\q[10]_BAR (
        div_norm_inv[10]), .\q[9]_BAR (div_norm_inv[9]), .\q[8]_BAR (
        div_norm_inv[8]), .\q[7]_BAR (div_norm_inv[7]), .\q[6]_BAR (
        div_norm_inv[6]), .\q[5]_BAR (div_norm_inv[5]), .\q[4]_BAR (
        div_norm_inv[4]), .\q[3]_BAR (div_norm_inv[3]), .\q[2]_BAR (
        div_norm_inv[2]), .\q[1]_BAR (div_norm_inv[1]), .\q[0]_BAR (
        div_norm_inv[0]) );
  fpu_cnt_lead0_53b_1 i_div_lead0 ( .din(div_norm_inv), .lead0(div_lead0) );
  dff_SIZE12 i_dstg_xtra_regs ( .din({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        div_lead0}), .clk(clk), .q({div_shl_cnta, div_shl_cnt}), .se(se), .si(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dff_SIZE53_1 i_div_shl_data ( .din(div_norm_inv), .clk(clk), .q(div_shl_data), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_5 i_div_shl_save ( .din({1'b0, 1'b0, div_shl_tmp}), .en(
        d3stg_fdiv), .clk(clk), .q({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, div_shl_save[52:0]}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_4 i_div_frac_add_in2 ( .din({1'b0, d4stg_fdiv, 
        div_frac_add_in2_in}), .en(div_frac_add_in2_load), .clk(clk), .q(
        div_frac_add_in2), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dffe_SIZE55_3 i_div_frac_add_in1 ( .din(div_frac_add_in1_in), .en(
        div_frac_add_in1_load), .clk(clk), .q(div_frac_add_in1), .se(se), .si(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_2 i_div_frac_add_in1a ( .din(div_frac_add_in1_in), .en(
        div_frac_add_in1_load), .clk(clk), .q(div_frac_add_in1a), .se(se), 
        .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dffe_SIZE55_1 i_div_frac_out ( .din(div_frac_out_in), .en(div_frac_out_load), 
        .clk(clk), .q({div_frac_out_54_53, \div_frac_out[52] , div_frac_outa}), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  OR3X1_RVT U2 ( .A1(n48), .A2(n47), .A3(n46), .Y(div_shl_tmp[98]) );
  INVX0_RVT U3 ( .A(div_shl_tmp[82]), .Y(n741) );
  INVX0_RVT U4 ( .A(n606), .Y(n522) );
  INVX0_RVT U5 ( .A(n640), .Y(n571) );
  INVX0_RVT U6 ( .A(n636), .Y(n574) );
  INVX0_RVT U7 ( .A(n709), .Y(n712) );
  INVX0_RVT U8 ( .A(n635), .Y(n637) );
  INVX0_RVT U9 ( .A(n618), .Y(n620) );
  INVX0_RVT U10 ( .A(n601), .Y(n603) );
  INVX0_RVT U11 ( .A(n599), .Y(n515) );
  INVX0_RVT U12 ( .A(n716), .Y(n585) );
  INVX0_RVT U13 ( .A(n711), .Y(n588) );
  INVX0_RVT U14 ( .A(n623), .Y(n558) );
  INVX0_RVT U15 ( .A(n619), .Y(n561) );
  INVX0_RVT U16 ( .A(n786), .Y(div_shl_tmp[53]) );
  INVX0_RVT U17 ( .A(div_norm_qnan), .Y(n50) );
  INVX0_RVT U18 ( .A(n736), .Y(n722) );
  AOI22X1_RVT U19 ( .A1(d4stg_fdiv), .A2(div_shl_save[14]), .A3(n795), .A4(
        n270), .Y(n1) );
  AOI22X1_RVT U20 ( .A1(d4stg_fdiv), .A2(div_shl_save[15]), .A3(n795), .A4(
        n273), .Y(n2) );
  AOI22X1_RVT U21 ( .A1(d4stg_fdiv), .A2(div_shl_save[16]), .A3(n795), .A4(
        n276), .Y(n3) );
  AOI22X1_RVT U22 ( .A1(d4stg_fdiv), .A2(div_shl_save[17]), .A3(n795), .A4(
        n279), .Y(n4) );
  AOI22X1_RVT U23 ( .A1(d4stg_fdiv), .A2(div_shl_save[18]), .A3(n795), .A4(
        n282), .Y(n5) );
  AOI22X1_RVT U24 ( .A1(d4stg_fdiv), .A2(div_shl_save[19]), .A3(n795), .A4(
        n285), .Y(n6) );
  AOI22X1_RVT U25 ( .A1(d4stg_fdiv), .A2(div_shl_save[20]), .A3(n795), .A4(
        n288), .Y(n7) );
  AOI22X1_RVT U26 ( .A1(d4stg_fdiv), .A2(div_shl_save[21]), .A3(n795), .A4(
        n291), .Y(n8) );
  AOI22X1_RVT U27 ( .A1(d4stg_fdiv), .A2(div_shl_save[22]), .A3(n795), .A4(
        n294), .Y(n9) );
  AOI22X1_RVT U28 ( .A1(d4stg_fdiv), .A2(div_shl_save[23]), .A3(n795), .A4(
        n297), .Y(n10) );
  AOI22X1_RVT U29 ( .A1(d4stg_fdiv), .A2(div_shl_save[24]), .A3(n795), .A4(
        n300), .Y(n11) );
  AOI22X1_RVT U30 ( .A1(d4stg_fdiv), .A2(div_shl_save[25]), .A3(n795), .A4(
        n303), .Y(n12) );
  AOI22X1_RVT U31 ( .A1(d4stg_fdiv), .A2(div_shl_save[26]), .A3(n795), .A4(
        n307), .Y(n13) );
  NAND2X0_RVT U32 ( .A1(d7stg_to_0), .A2(div_frac_out_of), .Y(n14) );
  INVX1_RVT U33 ( .A(n401), .Y(div_frac_add_52_inva) );
  INVX1_RVT U34 ( .A(se), .Y(n1028) );
  INVX1_RVT U35 ( .A(div_shl_cnta[0]), .Y(n16) );
  INVX1_RVT U36 ( .A(div_shl_cnta[1]), .Y(n15) );
  AND2X1_RVT U37 ( .A1(n16), .A2(n15), .Y(n408) );
  INVX1_RVT U38 ( .A(div_shl_cnta[2]), .Y(n521) );
  AND3X1_RVT U39 ( .A1(n408), .A2(div_shl_data[0]), .A3(n521), .Y(n607) );
  INVX1_RVT U40 ( .A(div_shl_cnta[5]), .Y(n775) );
  INVX1_RVT U41 ( .A(div_shl_cnta[4]), .Y(n774) );
  NAND2X0_RVT U42 ( .A1(n775), .A2(n774), .Y(n759) );
  INVX1_RVT U43 ( .A(n759), .Y(n25) );
  INVX1_RVT U44 ( .A(div_shl_cnta[3]), .Y(n779) );
  NAND3X0_RVT U45 ( .A1(n607), .A2(n25), .A3(n779), .Y(n786) );
  NAND2X0_RVT U46 ( .A1(div_shl_cnta[4]), .A2(n775), .Y(n758) );
  INVX1_RVT U47 ( .A(n758), .Y(n752) );
  AND2X1_RVT U48 ( .A1(div_shl_cnta[0]), .A2(n15), .Y(n425) );
  AO22X1_RVT U49 ( .A1(n408), .A2(div_shl_data[9]), .A3(n425), .A4(
        div_shl_data[8]), .Y(n18) );
  AND2X1_RVT U50 ( .A1(div_shl_cnta[0]), .A2(div_shl_cnta[1]), .Y(n22) );
  AND2X1_RVT U51 ( .A1(div_shl_cnta[1]), .A2(n16), .Y(n506) );
  AO22X1_RVT U52 ( .A1(n22), .A2(div_shl_data[6]), .A3(n506), .A4(
        div_shl_data[7]), .Y(n17) );
  OR2X1_RVT U53 ( .A1(n18), .A2(n17), .Y(n707) );
  NAND2X0_RVT U54 ( .A1(div_shl_cnta[2]), .A2(n779), .Y(n604) );
  INVX1_RVT U55 ( .A(n604), .Y(n715) );
  AO22X1_RVT U56 ( .A1(n408), .A2(div_shl_data[13]), .A3(n425), .A4(
        div_shl_data[12]), .Y(n20) );
  AO22X1_RVT U57 ( .A1(n22), .A2(div_shl_data[10]), .A3(n506), .A4(
        div_shl_data[11]), .Y(n19) );
  OR2X1_RVT U58 ( .A1(n20), .A2(n19), .Y(n709) );
  NAND2X0_RVT U59 ( .A1(n779), .A2(n521), .Y(n710) );
  INVX1_RVT U60 ( .A(n710), .Y(n21) );
  AO22X1_RVT U61 ( .A1(n408), .A2(div_shl_data[1]), .A3(div_shl_data[0]), .A4(
        n425), .Y(n784) );
  AO22X1_RVT U62 ( .A1(n408), .A2(div_shl_data[5]), .A3(n425), .A4(
        div_shl_data[4]), .Y(n24) );
  AO22X1_RVT U63 ( .A1(n22), .A2(div_shl_data[2]), .A3(n506), .A4(
        div_shl_data[3]), .Y(n23) );
  OR2X1_RVT U64 ( .A1(n24), .A2(n23), .Y(n501) );
  AO22X1_RVT U65 ( .A1(div_shl_cnta[2]), .A2(n784), .A3(n521), .A4(n501), .Y(
        n780) );
  AO222X1_RVT U66 ( .A1(n707), .A2(n715), .A3(n709), .A4(n21), .A5(n780), .A6(
        div_shl_cnta[3]), .Y(n769) );
  AO22X1_RVT U67 ( .A1(n408), .A2(div_shl_data[25]), .A3(n425), .A4(
        div_shl_data[24]), .Y(n27) );
  AO22X1_RVT U68 ( .A1(n22), .A2(div_shl_data[22]), .A3(n506), .A4(
        div_shl_data[23]), .Y(n26) );
  NOR2X0_RVT U69 ( .A1(n27), .A2(n26), .Y(n647) );
  AO22X1_RVT U70 ( .A1(n408), .A2(div_shl_data[29]), .A3(n425), .A4(
        div_shl_data[28]), .Y(n29) );
  AO22X1_RVT U71 ( .A1(n22), .A2(div_shl_data[26]), .A3(n506), .A4(
        div_shl_data[27]), .Y(n28) );
  NOR2X0_RVT U72 ( .A1(n29), .A2(n28), .Y(n649) );
  OA22X1_RVT U73 ( .A1(n647), .A2(n604), .A3(n649), .A4(n710), .Y(n36) );
  AO22X1_RVT U74 ( .A1(n408), .A2(div_shl_data[17]), .A3(n425), .A4(
        div_shl_data[16]), .Y(n31) );
  AO22X1_RVT U75 ( .A1(n22), .A2(div_shl_data[14]), .A3(n506), .A4(
        div_shl_data[15]), .Y(n30) );
  OR2X1_RVT U76 ( .A1(n31), .A2(n30), .Y(n716) );
  NAND2X0_RVT U77 ( .A1(div_shl_cnta[3]), .A2(div_shl_cnta[2]), .Y(n537) );
  AO22X1_RVT U78 ( .A1(n408), .A2(div_shl_data[21]), .A3(n425), .A4(
        div_shl_data[20]), .Y(n33) );
  AO22X1_RVT U79 ( .A1(n22), .A2(div_shl_data[18]), .A3(n506), .A4(
        div_shl_data[19]), .Y(n32) );
  NOR2X0_RVT U80 ( .A1(n33), .A2(n32), .Y(n711) );
  NAND2X0_RVT U81 ( .A1(div_shl_cnta[3]), .A2(n521), .Y(n34) );
  OA22X1_RVT U82 ( .A1(n585), .A2(n537), .A3(n711), .A4(n34), .Y(n35) );
  NAND2X0_RVT U83 ( .A1(n36), .A2(n35), .Y(n45) );
  AO22X1_RVT U84 ( .A1(n752), .A2(n769), .A3(n25), .A4(n45), .Y(
        div_shl_tmp[82]) );
  INVX1_RVT U85 ( .A(n34), .Y(n592) );
  NAND2X0_RVT U86 ( .A1(n592), .A2(n25), .Y(n648) );
  AO22X1_RVT U87 ( .A1(n408), .A2(div_shl_data[37]), .A3(n425), .A4(
        div_shl_data[36]), .Y(n38) );
  AO22X1_RVT U88 ( .A1(n22), .A2(div_shl_data[34]), .A3(n506), .A4(
        div_shl_data[35]), .Y(n37) );
  OR2X1_RVT U89 ( .A1(n38), .A2(n37), .Y(n582) );
  INVX1_RVT U90 ( .A(n582), .Y(n706) );
  INVX1_RVT U91 ( .A(n537), .Y(n708) );
  NAND2X0_RVT U92 ( .A1(n708), .A2(n25), .Y(n646) );
  AO22X1_RVT U93 ( .A1(n408), .A2(div_shl_data[33]), .A3(n425), .A4(
        div_shl_data[32]), .Y(n40) );
  AO22X1_RVT U94 ( .A1(n22), .A2(div_shl_data[30]), .A3(n506), .A4(
        div_shl_data[31]), .Y(n39) );
  NOR2X0_RVT U95 ( .A1(n40), .A2(n39), .Y(n704) );
  OAI22X1_RVT U96 ( .A1(n648), .A2(n706), .A3(n646), .A4(n704), .Y(n48) );
  NAND2X0_RVT U97 ( .A1(n715), .A2(n25), .Y(n650) );
  INVX1_RVT U98 ( .A(n650), .Y(n583) );
  AO22X1_RVT U99 ( .A1(n408), .A2(div_shl_data[41]), .A3(n425), .A4(
        div_shl_data[40]), .Y(n42) );
  AO22X1_RVT U100 ( .A1(n22), .A2(div_shl_data[38]), .A3(n506), .A4(
        div_shl_data[39]), .Y(n41) );
  OR2X1_RVT U101 ( .A1(n42), .A2(n41), .Y(n584) );
  NAND2X0_RVT U102 ( .A1(n21), .A2(n25), .Y(n705) );
  INVX1_RVT U103 ( .A(n705), .Y(n785) );
  AO22X1_RVT U104 ( .A1(n408), .A2(div_shl_data[45]), .A3(n425), .A4(
        div_shl_data[44]), .Y(n44) );
  AO22X1_RVT U105 ( .A1(n22), .A2(div_shl_data[42]), .A3(n506), .A4(
        div_shl_data[43]), .Y(n43) );
  OR2X1_RVT U106 ( .A1(n44), .A2(n43), .Y(n505) );
  AO22X1_RVT U107 ( .A1(n583), .A2(n584), .A3(n785), .A4(n505), .Y(n47) );
  NAND2X0_RVT U108 ( .A1(div_shl_cnta[5]), .A2(n774), .Y(n736) );
  AO22X1_RVT U109 ( .A1(n752), .A2(n45), .A3(n722), .A4(n769), .Y(n46) );
  AOI22X1_RVT U117 ( .A1(div_norm_frac_in2_sng_norm), .A2(div_frac_in2[32]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[29]), .Y(n51) );
  NAND2X0_RVT U118 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[29]), 
        .Y(n49) );
  AND3X1_RVT U119 ( .A1(n51), .A2(n50), .A3(n49), .Y(n54) );
  AOI22X1_RVT U120 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[28]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[32]), .Y(n53) );
  NAND2X0_RVT U121 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[28]), 
        .Y(n52) );
  AND3X1_RVT U122 ( .A1(n54), .A2(n53), .A3(n52), .Y(n680) );
  FADDX1_RVT U123 ( .A(div_frac_add_in1a[0]), .B(div_frac_add_in2[0]), .CI(
        d5stg_fdivb), .CO(n59), .S(n218) );
  FADDX1_RVT U124 ( .A(div_frac_add_in1a[52]), .B(div_frac_add_in2[52]), .CI(
        n55), .CO(n211), .S(n401) );
  FADDX1_RVT U125 ( .A(div_frac_add_in2[54]), .B(div_frac_add_in1a[54]), .CI(
        n56), .S(n217) );
  INVX1_RVT U126 ( .A(n217), .Y(n403) );
  AOI22X1_RVT U127 ( .A1(div_frac_out_add), .A2(n218), .A3(
        div_frac_out_shl1_dbl), .A4(n403), .Y(n58) );
  NAND2X0_RVT U128 ( .A1(div_frac_add_in1[0]), .A2(div_frac_out_add_in1), .Y(
        n57) );
  NAND3X0_RVT U129 ( .A1(n58), .A2(n14), .A3(n57), .Y(div_frac_out_in[0]) );
  FADDX1_RVT U130 ( .A(div_frac_add_in1a[1]), .B(div_frac_add_in2[1]), .CI(n59), .CO(n62), .S(n222) );
  AOI22X1_RVT U131 ( .A1(n222), .A2(div_frac_out_add), .A3(
        div_frac_out_shl1_dbl), .A4(div_frac_outa[0]), .Y(n61) );
  NAND2X0_RVT U132 ( .A1(div_frac_add_in1[1]), .A2(div_frac_out_add_in1), .Y(
        n60) );
  NAND3X0_RVT U133 ( .A1(n61), .A2(n14), .A3(n60), .Y(div_frac_out_in[1]) );
  FADDX1_RVT U134 ( .A(div_frac_add_in1a[2]), .B(div_frac_add_in2[2]), .CI(n62), .CO(n65), .S(n226) );
  AOI22X1_RVT U135 ( .A1(n226), .A2(div_frac_out_add), .A3(
        div_frac_out_shl1_dbl), .A4(div_frac_outa[1]), .Y(n64) );
  NAND2X0_RVT U136 ( .A1(div_frac_add_in1[2]), .A2(div_frac_out_add_in1), .Y(
        n63) );
  NAND3X0_RVT U137 ( .A1(n64), .A2(n14), .A3(n63), .Y(div_frac_out_in[2]) );
  FADDX1_RVT U138 ( .A(div_frac_add_in1a[3]), .B(div_frac_add_in2[3]), .CI(n65), .CO(n68), .S(n230) );
  AOI22X1_RVT U139 ( .A1(n230), .A2(div_frac_out_add), .A3(div_frac_outa[2]), 
        .A4(div_frac_out_shl1_dbl), .Y(n67) );
  NAND2X0_RVT U140 ( .A1(div_frac_add_in1[3]), .A2(div_frac_out_add_in1), .Y(
        n66) );
  NAND3X0_RVT U141 ( .A1(n67), .A2(n14), .A3(n66), .Y(div_frac_out_in[3]) );
  FADDX1_RVT U142 ( .A(div_frac_add_in1a[4]), .B(div_frac_add_in2[4]), .CI(n68), .CO(n71), .S(n234) );
  AOI22X1_RVT U143 ( .A1(n234), .A2(div_frac_out_add), .A3(div_frac_outa[3]), 
        .A4(div_frac_out_shl1_dbl), .Y(n70) );
  NAND2X0_RVT U144 ( .A1(div_frac_add_in1[4]), .A2(div_frac_out_add_in1), .Y(
        n69) );
  NAND3X0_RVT U145 ( .A1(n70), .A2(n14), .A3(n69), .Y(div_frac_out_in[4]) );
  FADDX1_RVT U146 ( .A(div_frac_add_in1a[5]), .B(div_frac_add_in2[5]), .CI(n71), .CO(n74), .S(n238) );
  AOI22X1_RVT U147 ( .A1(n238), .A2(div_frac_out_add), .A3(div_frac_outa[4]), 
        .A4(div_frac_out_shl1_dbl), .Y(n73) );
  NAND2X0_RVT U148 ( .A1(div_frac_add_in1[5]), .A2(div_frac_out_add_in1), .Y(
        n72) );
  NAND3X0_RVT U149 ( .A1(n73), .A2(n14), .A3(n72), .Y(div_frac_out_in[5]) );
  FADDX1_RVT U150 ( .A(div_frac_add_in1a[6]), .B(div_frac_add_in2[6]), .CI(n74), .CO(n77), .S(n242) );
  AOI22X1_RVT U151 ( .A1(n242), .A2(div_frac_out_add), .A3(div_frac_outa[5]), 
        .A4(div_frac_out_shl1_dbl), .Y(n76) );
  NAND2X0_RVT U152 ( .A1(div_frac_add_in1[6]), .A2(div_frac_out_add_in1), .Y(
        n75) );
  NAND3X0_RVT U153 ( .A1(n76), .A2(n14), .A3(n75), .Y(div_frac_out_in[6]) );
  FADDX1_RVT U154 ( .A(div_frac_add_in1a[7]), .B(div_frac_add_in2[7]), .CI(n77), .CO(n80), .S(n246) );
  AOI22X1_RVT U155 ( .A1(n246), .A2(div_frac_out_add), .A3(div_frac_outa[6]), 
        .A4(div_frac_out_shl1_dbl), .Y(n79) );
  NAND2X0_RVT U156 ( .A1(div_frac_add_in1[7]), .A2(div_frac_out_add_in1), .Y(
        n78) );
  NAND3X0_RVT U157 ( .A1(n79), .A2(n14), .A3(n78), .Y(div_frac_out_in[7]) );
  FADDX1_RVT U158 ( .A(div_frac_add_in1a[8]), .B(div_frac_add_in2[8]), .CI(n80), .CO(n83), .S(n250) );
  AOI22X1_RVT U159 ( .A1(n250), .A2(div_frac_out_add), .A3(div_frac_outa[7]), 
        .A4(div_frac_out_shl1_dbl), .Y(n82) );
  NAND2X0_RVT U160 ( .A1(div_frac_add_in1[8]), .A2(div_frac_out_add_in1), .Y(
        n81) );
  NAND3X0_RVT U161 ( .A1(n82), .A2(n14), .A3(n81), .Y(div_frac_out_in[8]) );
  FADDX1_RVT U162 ( .A(div_frac_add_in1a[9]), .B(div_frac_add_in2[9]), .CI(n83), .CO(n86), .S(n254) );
  AOI22X1_RVT U163 ( .A1(n254), .A2(div_frac_out_add), .A3(div_frac_outa[8]), 
        .A4(div_frac_out_shl1_dbl), .Y(n85) );
  NAND2X0_RVT U164 ( .A1(div_frac_add_in1[9]), .A2(div_frac_out_add_in1), .Y(
        n84) );
  NAND3X0_RVT U165 ( .A1(n85), .A2(n14), .A3(n84), .Y(div_frac_out_in[9]) );
  FADDX1_RVT U166 ( .A(div_frac_add_in1a[10]), .B(div_frac_add_in2[10]), .CI(
        n86), .CO(n89), .S(n258) );
  AOI22X1_RVT U167 ( .A1(n258), .A2(div_frac_out_add), .A3(div_frac_outa[9]), 
        .A4(div_frac_out_shl1_dbl), .Y(n88) );
  NAND2X0_RVT U168 ( .A1(div_frac_add_in1[10]), .A2(div_frac_out_add_in1), .Y(
        n87) );
  NAND3X0_RVT U169 ( .A1(n88), .A2(n14), .A3(n87), .Y(div_frac_out_in[10]) );
  FADDX1_RVT U170 ( .A(div_frac_add_in1a[11]), .B(div_frac_add_in2[11]), .CI(
        n89), .CO(n92), .S(n262) );
  AOI22X1_RVT U171 ( .A1(n262), .A2(div_frac_out_add), .A3(div_frac_outa[10]), 
        .A4(div_frac_out_shl1_dbl), .Y(n91) );
  NAND2X0_RVT U172 ( .A1(div_frac_add_in1[11]), .A2(div_frac_out_add_in1), .Y(
        n90) );
  NAND3X0_RVT U173 ( .A1(n91), .A2(n14), .A3(n90), .Y(div_frac_out_in[11]) );
  FADDX1_RVT U174 ( .A(div_frac_add_in1a[12]), .B(div_frac_add_in2[12]), .CI(
        n92), .CO(n95), .S(n266) );
  AOI22X1_RVT U175 ( .A1(n266), .A2(div_frac_out_add), .A3(div_frac_outa[11]), 
        .A4(div_frac_out_shl1_dbl), .Y(n94) );
  NAND2X0_RVT U176 ( .A1(div_frac_add_in1[12]), .A2(div_frac_out_add_in1), .Y(
        n93) );
  NAND3X0_RVT U177 ( .A1(n94), .A2(n14), .A3(n93), .Y(div_frac_out_in[12]) );
  FADDX1_RVT U178 ( .A(div_frac_add_in1a[13]), .B(div_frac_add_in2[13]), .CI(
        n95), .CO(n98), .S(n270) );
  AOI22X1_RVT U179 ( .A1(n270), .A2(div_frac_out_add), .A3(div_frac_outa[12]), 
        .A4(div_frac_out_shl1_dbl), .Y(n97) );
  NAND2X0_RVT U180 ( .A1(div_frac_add_in1[13]), .A2(div_frac_out_add_in1), .Y(
        n96) );
  NAND3X0_RVT U181 ( .A1(n97), .A2(n14), .A3(n96), .Y(div_frac_out_in[13]) );
  FADDX1_RVT U182 ( .A(div_frac_add_in1a[14]), .B(div_frac_add_in2[14]), .CI(
        n98), .CO(n101), .S(n273) );
  AOI22X1_RVT U183 ( .A1(n273), .A2(div_frac_out_add), .A3(div_frac_outa[13]), 
        .A4(div_frac_out_shl1_dbl), .Y(n100) );
  NAND2X0_RVT U184 ( .A1(div_frac_add_in1[14]), .A2(div_frac_out_add_in1), .Y(
        n99) );
  NAND3X0_RVT U185 ( .A1(n100), .A2(n14), .A3(n99), .Y(div_frac_out_in[14]) );
  FADDX1_RVT U186 ( .A(div_frac_add_in1a[15]), .B(div_frac_add_in2[15]), .CI(
        n101), .CO(n104), .S(n276) );
  AOI22X1_RVT U187 ( .A1(n276), .A2(div_frac_out_add), .A3(div_frac_outa[14]), 
        .A4(div_frac_out_shl1_dbl), .Y(n103) );
  NAND2X0_RVT U188 ( .A1(div_frac_add_in1[15]), .A2(div_frac_out_add_in1), .Y(
        n102) );
  NAND3X0_RVT U189 ( .A1(n103), .A2(n14), .A3(n102), .Y(div_frac_out_in[15])
         );
  FADDX1_RVT U190 ( .A(div_frac_add_in1a[16]), .B(div_frac_add_in2[16]), .CI(
        n104), .CO(n107), .S(n279) );
  AOI22X1_RVT U191 ( .A1(n279), .A2(div_frac_out_add), .A3(div_frac_outa[15]), 
        .A4(div_frac_out_shl1_dbl), .Y(n106) );
  NAND2X0_RVT U192 ( .A1(div_frac_add_in1[16]), .A2(div_frac_out_add_in1), .Y(
        n105) );
  NAND3X0_RVT U193 ( .A1(n106), .A2(n14), .A3(n105), .Y(div_frac_out_in[16])
         );
  FADDX1_RVT U194 ( .A(div_frac_add_in1a[17]), .B(div_frac_add_in2[17]), .CI(
        n107), .CO(n110), .S(n282) );
  AOI22X1_RVT U195 ( .A1(n282), .A2(div_frac_out_add), .A3(div_frac_outa[16]), 
        .A4(div_frac_out_shl1_dbl), .Y(n109) );
  NAND2X0_RVT U196 ( .A1(div_frac_add_in1[17]), .A2(div_frac_out_add_in1), .Y(
        n108) );
  NAND3X0_RVT U197 ( .A1(n109), .A2(n14), .A3(n108), .Y(div_frac_out_in[17])
         );
  FADDX1_RVT U198 ( .A(div_frac_add_in1a[18]), .B(div_frac_add_in2[18]), .CI(
        n110), .CO(n113), .S(n285) );
  AOI22X1_RVT U199 ( .A1(n285), .A2(div_frac_out_add), .A3(div_frac_outa[17]), 
        .A4(div_frac_out_shl1_dbl), .Y(n112) );
  NAND2X0_RVT U200 ( .A1(div_frac_add_in1[18]), .A2(div_frac_out_add_in1), .Y(
        n111) );
  NAND3X0_RVT U201 ( .A1(n112), .A2(n14), .A3(n111), .Y(div_frac_out_in[18])
         );
  FADDX1_RVT U202 ( .A(div_frac_add_in1a[19]), .B(div_frac_add_in2[19]), .CI(
        n113), .CO(n116), .S(n288) );
  AOI22X1_RVT U203 ( .A1(n288), .A2(div_frac_out_add), .A3(div_frac_outa[18]), 
        .A4(div_frac_out_shl1_dbl), .Y(n115) );
  NAND2X0_RVT U204 ( .A1(div_frac_add_in1[19]), .A2(div_frac_out_add_in1), .Y(
        n114) );
  NAND3X0_RVT U205 ( .A1(n115), .A2(n14), .A3(n114), .Y(div_frac_out_in[19])
         );
  FADDX1_RVT U206 ( .A(div_frac_add_in1a[20]), .B(div_frac_add_in2[20]), .CI(
        n116), .CO(n119), .S(n291) );
  AOI22X1_RVT U207 ( .A1(n291), .A2(div_frac_out_add), .A3(div_frac_outa[19]), 
        .A4(div_frac_out_shl1_dbl), .Y(n118) );
  NAND2X0_RVT U208 ( .A1(div_frac_add_in1[20]), .A2(div_frac_out_add_in1), .Y(
        n117) );
  NAND3X0_RVT U209 ( .A1(n118), .A2(n14), .A3(n117), .Y(div_frac_out_in[20])
         );
  FADDX1_RVT U210 ( .A(div_frac_add_in1a[21]), .B(div_frac_add_in2[21]), .CI(
        n119), .CO(n122), .S(n294) );
  AOI22X1_RVT U211 ( .A1(n294), .A2(div_frac_out_add), .A3(div_frac_outa[20]), 
        .A4(div_frac_out_shl1_dbl), .Y(n121) );
  NAND2X0_RVT U212 ( .A1(div_frac_add_in1[21]), .A2(div_frac_out_add_in1), .Y(
        n120) );
  NAND3X0_RVT U213 ( .A1(n121), .A2(n14), .A3(n120), .Y(div_frac_out_in[21])
         );
  FADDX1_RVT U214 ( .A(div_frac_add_in1a[22]), .B(div_frac_add_in2[22]), .CI(
        n122), .CO(n125), .S(n297) );
  AOI22X1_RVT U215 ( .A1(n297), .A2(div_frac_out_add), .A3(div_frac_outa[21]), 
        .A4(div_frac_out_shl1_dbl), .Y(n124) );
  NAND2X0_RVT U216 ( .A1(div_frac_add_in1[22]), .A2(div_frac_out_add_in1), .Y(
        n123) );
  NAND3X0_RVT U217 ( .A1(n124), .A2(n14), .A3(n123), .Y(div_frac_out_in[22])
         );
  FADDX1_RVT U218 ( .A(div_frac_add_in1a[23]), .B(div_frac_add_in2[23]), .CI(
        n125), .CO(n128), .S(n300) );
  AOI22X1_RVT U219 ( .A1(n300), .A2(div_frac_out_add), .A3(div_frac_outa[22]), 
        .A4(div_frac_out_shl1_dbl), .Y(n127) );
  NAND2X0_RVT U220 ( .A1(div_frac_add_in1[23]), .A2(div_frac_out_add_in1), .Y(
        n126) );
  NAND3X0_RVT U221 ( .A1(n127), .A2(n14), .A3(n126), .Y(div_frac_out_in[23])
         );
  FADDX1_RVT U222 ( .A(div_frac_add_in1a[24]), .B(div_frac_add_in2[24]), .CI(
        n128), .CO(n131), .S(n303) );
  AOI22X1_RVT U223 ( .A1(n303), .A2(div_frac_out_add), .A3(div_frac_outa[23]), 
        .A4(div_frac_out_shl1_dbl), .Y(n130) );
  NAND2X0_RVT U224 ( .A1(div_frac_add_in1[24]), .A2(div_frac_out_add_in1), .Y(
        n129) );
  NAND3X0_RVT U225 ( .A1(n130), .A2(n14), .A3(n129), .Y(div_frac_out_in[24])
         );
  FADDX1_RVT U226 ( .A(div_frac_add_in1a[25]), .B(div_frac_add_in2[25]), .CI(
        n131), .CO(n134), .S(n307) );
  AOI22X1_RVT U227 ( .A1(n307), .A2(div_frac_out_add), .A3(div_frac_outa[24]), 
        .A4(div_frac_out_shl1_dbl), .Y(n133) );
  NAND2X0_RVT U228 ( .A1(div_frac_add_in1[25]), .A2(div_frac_out_add_in1), .Y(
        n132) );
  NAND3X0_RVT U229 ( .A1(n133), .A2(n14), .A3(n132), .Y(div_frac_out_in[25])
         );
  FADDX1_RVT U230 ( .A(div_frac_add_in1a[26]), .B(div_frac_add_in2[26]), .CI(
        n134), .CO(n137), .S(n794) );
  AOI22X1_RVT U231 ( .A1(div_frac_outa[25]), .A2(div_frac_out_shl1_dbl), .A3(
        n794), .A4(div_frac_out_add), .Y(n136) );
  NAND2X0_RVT U232 ( .A1(div_frac_add_in1[26]), .A2(div_frac_out_add_in1), .Y(
        n135) );
  NAND3X0_RVT U233 ( .A1(n136), .A2(n14), .A3(n135), .Y(div_frac_out_in[26])
         );
  FADDX1_RVT U234 ( .A(div_frac_add_in1a[27]), .B(div_frac_add_in2[27]), .CI(
        n137), .CO(n140), .S(n791) );
  AOI22X1_RVT U235 ( .A1(div_frac_outa[26]), .A2(div_frac_out_shl1_dbl), .A3(
        n791), .A4(div_frac_out_add), .Y(n139) );
  NAND2X0_RVT U236 ( .A1(div_frac_add_in1[27]), .A2(div_frac_out_add_in1), .Y(
        n138) );
  NAND3X0_RVT U237 ( .A1(n139), .A2(n14), .A3(n138), .Y(div_frac_out_in[27])
         );
  FADDX1_RVT U238 ( .A(div_frac_add_in1a[28]), .B(div_frac_add_in2[28]), .CI(
        n140), .CO(n311), .S(n788) );
  AOI22X1_RVT U239 ( .A1(div_frac_outa[27]), .A2(div_frac_out_shl1_dbl), .A3(
        n788), .A4(div_frac_out_add), .Y(n142) );
  NAND2X0_RVT U240 ( .A1(div_frac_add_in1[28]), .A2(div_frac_out_add_in1), .Y(
        n141) );
  NAND3X0_RVT U241 ( .A1(n142), .A2(n14), .A3(n141), .Y(div_frac_out_in[28])
         );
  FADDX1_RVT U242 ( .A(div_frac_add_in1a[30]), .B(div_frac_add_in2[30]), .CI(
        n143), .CO(n146), .S(n315) );
  OR2X1_RVT U243 ( .A1(div_frac_out_shl1_dbl), .A2(div_frac_out_shl1_sng), .Y(
        n214) );
  AOI22X1_RVT U244 ( .A1(n315), .A2(div_frac_out_add), .A3(div_frac_outa[29]), 
        .A4(n214), .Y(n145) );
  NAND2X0_RVT U245 ( .A1(div_frac_add_in1[30]), .A2(div_frac_out_add_in1), .Y(
        n144) );
  NAND3X0_RVT U246 ( .A1(n145), .A2(n14), .A3(n144), .Y(div_frac_out_in[30])
         );
  FADDX1_RVT U247 ( .A(div_frac_add_in1a[31]), .B(div_frac_add_in2[31]), .CI(
        n146), .CO(n149), .S(n319) );
  AOI22X1_RVT U248 ( .A1(n319), .A2(div_frac_out_add), .A3(div_frac_outa[30]), 
        .A4(n214), .Y(n148) );
  NAND2X0_RVT U249 ( .A1(div_frac_add_in1[31]), .A2(div_frac_out_add_in1), .Y(
        n147) );
  NAND3X0_RVT U250 ( .A1(n148), .A2(n14), .A3(n147), .Y(div_frac_out_in[31])
         );
  FADDX1_RVT U251 ( .A(div_frac_add_in1a[32]), .B(div_frac_add_in2[32]), .CI(
        n149), .CO(n152), .S(n323) );
  AOI22X1_RVT U252 ( .A1(n323), .A2(div_frac_out_add), .A3(div_frac_outa[31]), 
        .A4(n214), .Y(n151) );
  NAND2X0_RVT U253 ( .A1(div_frac_add_in1[32]), .A2(div_frac_out_add_in1), .Y(
        n150) );
  NAND3X0_RVT U254 ( .A1(n151), .A2(n14), .A3(n150), .Y(div_frac_out_in[32])
         );
  FADDX1_RVT U255 ( .A(div_frac_add_in1a[33]), .B(div_frac_add_in2[33]), .CI(
        n152), .CO(n155), .S(n327) );
  AOI22X1_RVT U256 ( .A1(n327), .A2(div_frac_out_add), .A3(div_frac_outa[32]), 
        .A4(n214), .Y(n154) );
  NAND2X0_RVT U257 ( .A1(div_frac_add_in1[33]), .A2(div_frac_out_add_in1), .Y(
        n153) );
  NAND3X0_RVT U258 ( .A1(n154), .A2(n14), .A3(n153), .Y(div_frac_out_in[33])
         );
  FADDX1_RVT U259 ( .A(div_frac_add_in1a[34]), .B(div_frac_add_in2[34]), .CI(
        n155), .CO(n158), .S(n331) );
  AOI22X1_RVT U260 ( .A1(n331), .A2(div_frac_out_add), .A3(div_frac_outa[33]), 
        .A4(n214), .Y(n157) );
  NAND2X0_RVT U261 ( .A1(div_frac_add_in1[34]), .A2(div_frac_out_add_in1), .Y(
        n156) );
  NAND3X0_RVT U262 ( .A1(n157), .A2(n14), .A3(n156), .Y(div_frac_out_in[34])
         );
  FADDX1_RVT U263 ( .A(div_frac_add_in1a[35]), .B(div_frac_add_in2[35]), .CI(
        n158), .CO(n161), .S(n335) );
  AOI22X1_RVT U264 ( .A1(n335), .A2(div_frac_out_add), .A3(div_frac_outa[34]), 
        .A4(n214), .Y(n160) );
  NAND2X0_RVT U265 ( .A1(div_frac_add_in1[35]), .A2(div_frac_out_add_in1), .Y(
        n159) );
  NAND3X0_RVT U266 ( .A1(n160), .A2(n14), .A3(n159), .Y(div_frac_out_in[35])
         );
  FADDX1_RVT U267 ( .A(div_frac_add_in1a[36]), .B(div_frac_add_in2[36]), .CI(
        n161), .CO(n164), .S(n339) );
  AOI22X1_RVT U268 ( .A1(n339), .A2(div_frac_out_add), .A3(div_frac_outa[35]), 
        .A4(n214), .Y(n163) );
  NAND2X0_RVT U269 ( .A1(div_frac_add_in1[36]), .A2(div_frac_out_add_in1), .Y(
        n162) );
  NAND3X0_RVT U270 ( .A1(n163), .A2(n14), .A3(n162), .Y(div_frac_out_in[36])
         );
  FADDX1_RVT U271 ( .A(div_frac_add_in1a[37]), .B(div_frac_add_in2[37]), .CI(
        n164), .CO(n167), .S(n343) );
  AOI22X1_RVT U272 ( .A1(n343), .A2(div_frac_out_add), .A3(div_frac_outa[36]), 
        .A4(n214), .Y(n166) );
  NAND2X0_RVT U273 ( .A1(div_frac_add_in1[37]), .A2(div_frac_out_add_in1), .Y(
        n165) );
  NAND3X0_RVT U274 ( .A1(n166), .A2(n14), .A3(n165), .Y(div_frac_out_in[37])
         );
  FADDX1_RVT U275 ( .A(div_frac_add_in1a[38]), .B(div_frac_add_in2[38]), .CI(
        n167), .CO(n170), .S(n347) );
  AOI22X1_RVT U276 ( .A1(n347), .A2(div_frac_out_add), .A3(div_frac_outa[37]), 
        .A4(n214), .Y(n169) );
  NAND2X0_RVT U277 ( .A1(div_frac_add_in1[38]), .A2(div_frac_out_add_in1), .Y(
        n168) );
  NAND3X0_RVT U278 ( .A1(n169), .A2(n14), .A3(n168), .Y(div_frac_out_in[38])
         );
  FADDX1_RVT U279 ( .A(div_frac_add_in1a[39]), .B(div_frac_add_in2[39]), .CI(
        n170), .CO(n173), .S(n351) );
  AOI22X1_RVT U280 ( .A1(n351), .A2(div_frac_out_add), .A3(div_frac_outa[38]), 
        .A4(n214), .Y(n172) );
  NAND2X0_RVT U281 ( .A1(div_frac_add_in1[39]), .A2(div_frac_out_add_in1), .Y(
        n171) );
  NAND3X0_RVT U282 ( .A1(n172), .A2(n14), .A3(n171), .Y(div_frac_out_in[39])
         );
  FADDX1_RVT U283 ( .A(div_frac_add_in1a[40]), .B(div_frac_add_in2[40]), .CI(
        n173), .CO(n176), .S(n355) );
  AOI22X1_RVT U284 ( .A1(n355), .A2(div_frac_out_add), .A3(div_frac_outa[39]), 
        .A4(n214), .Y(n175) );
  NAND2X0_RVT U285 ( .A1(div_frac_add_in1[40]), .A2(div_frac_out_add_in1), .Y(
        n174) );
  NAND3X0_RVT U286 ( .A1(n175), .A2(n14), .A3(n174), .Y(div_frac_out_in[40])
         );
  FADDX1_RVT U287 ( .A(div_frac_add_in1a[41]), .B(div_frac_add_in2[41]), .CI(
        n176), .CO(n179), .S(n359) );
  AOI22X1_RVT U288 ( .A1(n359), .A2(div_frac_out_add), .A3(div_frac_outa[40]), 
        .A4(n214), .Y(n178) );
  NAND2X0_RVT U289 ( .A1(div_frac_add_in1[41]), .A2(div_frac_out_add_in1), .Y(
        n177) );
  NAND3X0_RVT U290 ( .A1(n178), .A2(n14), .A3(n177), .Y(div_frac_out_in[41])
         );
  FADDX1_RVT U291 ( .A(div_frac_add_in1a[42]), .B(div_frac_add_in2[42]), .CI(
        n179), .CO(n182), .S(n363) );
  AOI22X1_RVT U292 ( .A1(n363), .A2(div_frac_out_add), .A3(div_frac_outa[41]), 
        .A4(n214), .Y(n181) );
  NAND2X0_RVT U293 ( .A1(div_frac_add_in1[42]), .A2(div_frac_out_add_in1), .Y(
        n180) );
  NAND3X0_RVT U294 ( .A1(n181), .A2(n14), .A3(n180), .Y(div_frac_out_in[42])
         );
  FADDX1_RVT U295 ( .A(div_frac_add_in1a[43]), .B(div_frac_add_in2[43]), .CI(
        n182), .CO(n185), .S(n367) );
  AOI22X1_RVT U296 ( .A1(n367), .A2(div_frac_out_add), .A3(div_frac_outa[42]), 
        .A4(n214), .Y(n184) );
  NAND2X0_RVT U297 ( .A1(div_frac_add_in1[43]), .A2(div_frac_out_add_in1), .Y(
        n183) );
  NAND3X0_RVT U298 ( .A1(n184), .A2(n14), .A3(n183), .Y(div_frac_out_in[43])
         );
  FADDX1_RVT U299 ( .A(div_frac_add_in1a[44]), .B(div_frac_add_in2[44]), .CI(
        n185), .CO(n188), .S(n371) );
  AOI22X1_RVT U300 ( .A1(n371), .A2(div_frac_out_add), .A3(div_frac_outa[43]), 
        .A4(n214), .Y(n187) );
  NAND2X0_RVT U301 ( .A1(div_frac_add_in1[44]), .A2(div_frac_out_add_in1), .Y(
        n186) );
  NAND3X0_RVT U302 ( .A1(n187), .A2(n14), .A3(n186), .Y(div_frac_out_in[44])
         );
  FADDX1_RVT U303 ( .A(div_frac_add_in1a[45]), .B(div_frac_add_in2[45]), .CI(
        n188), .CO(n191), .S(n375) );
  AOI22X1_RVT U304 ( .A1(n375), .A2(div_frac_out_add), .A3(div_frac_outa[44]), 
        .A4(n214), .Y(n190) );
  NAND2X0_RVT U305 ( .A1(div_frac_add_in1[45]), .A2(div_frac_out_add_in1), .Y(
        n189) );
  NAND3X0_RVT U306 ( .A1(n190), .A2(n14), .A3(n189), .Y(div_frac_out_in[45])
         );
  FADDX1_RVT U307 ( .A(div_frac_add_in1a[46]), .B(div_frac_add_in2[46]), .CI(
        n191), .CO(n194), .S(n379) );
  AOI22X1_RVT U308 ( .A1(n379), .A2(div_frac_out_add), .A3(div_frac_outa[45]), 
        .A4(n214), .Y(n193) );
  NAND2X0_RVT U309 ( .A1(div_frac_add_in1[46]), .A2(div_frac_out_add_in1), .Y(
        n192) );
  NAND3X0_RVT U310 ( .A1(n193), .A2(n14), .A3(n192), .Y(div_frac_out_in[46])
         );
  FADDX1_RVT U311 ( .A(div_frac_add_in1a[47]), .B(div_frac_add_in2[47]), .CI(
        n194), .CO(n197), .S(n383) );
  AOI22X1_RVT U312 ( .A1(n383), .A2(div_frac_out_add), .A3(div_frac_outa[46]), 
        .A4(n214), .Y(n196) );
  NAND2X0_RVT U313 ( .A1(div_frac_add_in1[47]), .A2(div_frac_out_add_in1), .Y(
        n195) );
  NAND3X0_RVT U314 ( .A1(n196), .A2(n14), .A3(n195), .Y(div_frac_out_in[47])
         );
  FADDX1_RVT U315 ( .A(div_frac_add_in1a[48]), .B(div_frac_add_in2[48]), .CI(
        n197), .CO(n200), .S(n387) );
  AOI22X1_RVT U316 ( .A1(n387), .A2(div_frac_out_add), .A3(div_frac_outa[47]), 
        .A4(n214), .Y(n199) );
  NAND2X0_RVT U317 ( .A1(div_frac_add_in1[48]), .A2(div_frac_out_add_in1), .Y(
        n198) );
  NAND3X0_RVT U318 ( .A1(n199), .A2(n14), .A3(n198), .Y(div_frac_out_in[48])
         );
  FADDX1_RVT U319 ( .A(div_frac_add_in1a[49]), .B(div_frac_add_in2[49]), .CI(
        n200), .CO(n203), .S(n391) );
  AOI22X1_RVT U320 ( .A1(n391), .A2(div_frac_out_add), .A3(div_frac_outa[48]), 
        .A4(n214), .Y(n202) );
  NAND2X0_RVT U321 ( .A1(div_frac_add_in1[49]), .A2(div_frac_out_add_in1), .Y(
        n201) );
  NAND3X0_RVT U322 ( .A1(n202), .A2(n14), .A3(n201), .Y(div_frac_out_in[49])
         );
  FADDX1_RVT U323 ( .A(div_frac_add_in1a[50]), .B(div_frac_add_in2[50]), .CI(
        n203), .CO(n206), .S(n397) );
  AOI22X1_RVT U324 ( .A1(n397), .A2(div_frac_out_add), .A3(div_frac_outa[49]), 
        .A4(n214), .Y(n205) );
  NAND2X0_RVT U325 ( .A1(div_frac_add_in1[50]), .A2(div_frac_out_add_in1), .Y(
        n204) );
  NAND3X0_RVT U326 ( .A1(n205), .A2(n14), .A3(n204), .Y(div_frac_out_in[50])
         );
  FADDX1_RVT U327 ( .A(div_frac_add_in1a[51]), .B(div_frac_add_in2[51]), .CI(
        n206), .CO(n55), .S(n787) );
  AOI22X1_RVT U328 ( .A1(div_frac_outa[50]), .A2(n214), .A3(div_frac_out_add), 
        .A4(n787), .Y(n208) );
  NAND2X0_RVT U329 ( .A1(div_frac_add_in1[51]), .A2(div_frac_out_add_in1), .Y(
        n207) );
  NAND3X0_RVT U330 ( .A1(n208), .A2(n14), .A3(n207), .Y(div_frac_out_in[51])
         );
  AOI22X1_RVT U331 ( .A1(div_frac_outa[51]), .A2(n214), .A3(div_frac_out_add), 
        .A4(n401), .Y(n210) );
  NAND2X0_RVT U332 ( .A1(div_frac_add_in1[52]), .A2(div_frac_out_add_in1), .Y(
        n209) );
  NAND3X0_RVT U333 ( .A1(n210), .A2(n14), .A3(n209), .Y(div_frac_out_in[52])
         );
  FADDX1_RVT U334 ( .A(div_frac_add_in1a[53]), .B(div_frac_add_in2[53]), .CI(
        n211), .CO(n56), .S(n402) );
  AOI22X1_RVT U335 ( .A1(\div_frac_out[52] ), .A2(n214), .A3(div_frac_out_add), 
        .A4(n402), .Y(n213) );
  NAND2X0_RVT U336 ( .A1(div_frac_add_in1[53]), .A2(div_frac_out_add_in1), .Y(
        n212) );
  NAND3X0_RVT U337 ( .A1(n213), .A2(n14), .A3(n212), .Y(div_frac_out_in[53])
         );
  AOI22X1_RVT U338 ( .A1(n217), .A2(div_frac_out_add), .A3(
        div_frac_out_54_53[0]), .A4(n214), .Y(n216) );
  NAND2X0_RVT U339 ( .A1(div_frac_add_in1[54]), .A2(div_frac_out_add_in1), .Y(
        n215) );
  NAND3X0_RVT U340 ( .A1(n216), .A2(n14), .A3(n215), .Y(div_frac_out_in[54])
         );
  AND2X2_RVT U341 ( .A1(div_frac_add_in1_add), .A2(n217), .Y(n796) );
  INVX1_RVT U342 ( .A(d6stg_frac_out_nosh), .Y(n799) );
  AND2X1_RVT U343 ( .A1(d6stg_fdiv), .A2(n799), .Y(n395) );
  AND2X1_RVT U344 ( .A1(d6stg_fdivd), .A2(n395), .Y(n306) );
  AOI22X1_RVT U345 ( .A1(div_frac_add_in1[0]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[2]), .Y(n221) );
  AND2X2_RVT U346 ( .A1(div_frac_add_in1_add), .A2(n403), .Y(n795) );
  AOI22X1_RVT U347 ( .A1(d4stg_fdiv), .A2(div_shl_save[1]), .A3(n795), .A4(
        n218), .Y(n220) );
  AND2X1_RVT U348 ( .A1(d6stg_fdiv), .A2(d6stg_frac_out_nosh), .Y(n396) );
  AND2X1_RVT U349 ( .A1(d6stg_fdivd), .A2(n396), .Y(n308) );
  NAND2X0_RVT U350 ( .A1(n308), .A2(div_frac_outa[3]), .Y(n219) );
  NAND3X0_RVT U351 ( .A1(n221), .A2(n220), .A3(n219), .Y(
        div_frac_add_in1_in[1]) );
  AOI22X1_RVT U352 ( .A1(div_frac_add_in1[1]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[3]), .Y(n225) );
  AOI22X1_RVT U353 ( .A1(d4stg_fdiv), .A2(div_shl_save[2]), .A3(n795), .A4(
        n222), .Y(n224) );
  NAND2X0_RVT U354 ( .A1(n308), .A2(div_frac_outa[4]), .Y(n223) );
  NAND3X0_RVT U355 ( .A1(n225), .A2(n224), .A3(n223), .Y(
        div_frac_add_in1_in[2]) );
  AOI22X1_RVT U356 ( .A1(div_frac_add_in1[2]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[4]), .Y(n229) );
  AOI22X1_RVT U357 ( .A1(d4stg_fdiv), .A2(div_shl_save[3]), .A3(n795), .A4(
        n226), .Y(n228) );
  NAND2X0_RVT U358 ( .A1(n308), .A2(div_frac_outa[5]), .Y(n227) );
  NAND3X0_RVT U359 ( .A1(n229), .A2(n228), .A3(n227), .Y(
        div_frac_add_in1_in[3]) );
  AOI22X1_RVT U360 ( .A1(div_frac_add_in1[3]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[5]), .Y(n233) );
  AOI22X1_RVT U361 ( .A1(d4stg_fdiv), .A2(div_shl_save[4]), .A3(n795), .A4(
        n230), .Y(n232) );
  NAND2X0_RVT U362 ( .A1(n308), .A2(div_frac_outa[6]), .Y(n231) );
  NAND3X0_RVT U363 ( .A1(n233), .A2(n232), .A3(n231), .Y(
        div_frac_add_in1_in[4]) );
  AOI22X1_RVT U364 ( .A1(div_frac_add_in1[4]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[6]), .Y(n237) );
  AOI22X1_RVT U365 ( .A1(d4stg_fdiv), .A2(div_shl_save[5]), .A3(n795), .A4(
        n234), .Y(n236) );
  NAND2X0_RVT U366 ( .A1(n308), .A2(div_frac_outa[7]), .Y(n235) );
  NAND3X0_RVT U367 ( .A1(n237), .A2(n236), .A3(n235), .Y(
        div_frac_add_in1_in[5]) );
  AOI22X1_RVT U368 ( .A1(div_frac_add_in1[5]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[7]), .Y(n241) );
  AOI22X1_RVT U369 ( .A1(d4stg_fdiv), .A2(div_shl_save[6]), .A3(n795), .A4(
        n238), .Y(n240) );
  NAND2X0_RVT U370 ( .A1(n308), .A2(div_frac_outa[8]), .Y(n239) );
  NAND3X0_RVT U371 ( .A1(n241), .A2(n240), .A3(n239), .Y(
        div_frac_add_in1_in[6]) );
  AOI22X1_RVT U372 ( .A1(div_frac_add_in1[6]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[8]), .Y(n245) );
  AOI22X1_RVT U373 ( .A1(d4stg_fdiv), .A2(div_shl_save[7]), .A3(n795), .A4(
        n242), .Y(n244) );
  NAND2X0_RVT U374 ( .A1(n308), .A2(div_frac_outa[9]), .Y(n243) );
  NAND3X0_RVT U375 ( .A1(n245), .A2(n244), .A3(n243), .Y(
        div_frac_add_in1_in[7]) );
  AOI22X1_RVT U376 ( .A1(div_frac_add_in1[7]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[9]), .Y(n249) );
  AOI22X1_RVT U377 ( .A1(d4stg_fdiv), .A2(div_shl_save[8]), .A3(n795), .A4(
        n246), .Y(n248) );
  NAND2X0_RVT U378 ( .A1(n308), .A2(div_frac_outa[10]), .Y(n247) );
  NAND3X0_RVT U379 ( .A1(n249), .A2(n248), .A3(n247), .Y(
        div_frac_add_in1_in[8]) );
  AOI22X1_RVT U380 ( .A1(div_frac_add_in1[8]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[10]), .Y(n253) );
  AOI22X1_RVT U381 ( .A1(d4stg_fdiv), .A2(div_shl_save[9]), .A3(n795), .A4(
        n250), .Y(n252) );
  NAND2X0_RVT U382 ( .A1(n308), .A2(div_frac_outa[11]), .Y(n251) );
  NAND3X0_RVT U383 ( .A1(n253), .A2(n252), .A3(n251), .Y(
        div_frac_add_in1_in[9]) );
  AOI22X1_RVT U384 ( .A1(div_frac_add_in1[9]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[11]), .Y(n257) );
  AOI22X1_RVT U385 ( .A1(d4stg_fdiv), .A2(div_shl_save[10]), .A3(n795), .A4(
        n254), .Y(n256) );
  NAND2X0_RVT U386 ( .A1(n308), .A2(div_frac_outa[12]), .Y(n255) );
  NAND3X0_RVT U387 ( .A1(n257), .A2(n256), .A3(n255), .Y(
        div_frac_add_in1_in[10]) );
  AOI22X1_RVT U388 ( .A1(div_frac_add_in1[10]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[12]), .Y(n261) );
  AOI22X1_RVT U389 ( .A1(d4stg_fdiv), .A2(div_shl_save[11]), .A3(n795), .A4(
        n258), .Y(n260) );
  NAND2X0_RVT U390 ( .A1(n308), .A2(div_frac_outa[13]), .Y(n259) );
  NAND3X0_RVT U391 ( .A1(n261), .A2(n260), .A3(n259), .Y(
        div_frac_add_in1_in[11]) );
  AOI22X1_RVT U392 ( .A1(div_frac_add_in1[11]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[13]), .Y(n265) );
  AOI22X1_RVT U393 ( .A1(d4stg_fdiv), .A2(div_shl_save[12]), .A3(n795), .A4(
        n262), .Y(n264) );
  NAND2X0_RVT U394 ( .A1(n308), .A2(div_frac_outa[14]), .Y(n263) );
  NAND3X0_RVT U395 ( .A1(n265), .A2(n264), .A3(n263), .Y(
        div_frac_add_in1_in[12]) );
  AOI22X1_RVT U396 ( .A1(div_frac_add_in1[12]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[14]), .Y(n269) );
  AOI22X1_RVT U397 ( .A1(d4stg_fdiv), .A2(div_shl_save[13]), .A3(n795), .A4(
        n266), .Y(n268) );
  NAND2X0_RVT U398 ( .A1(n308), .A2(div_frac_outa[15]), .Y(n267) );
  NAND3X0_RVT U399 ( .A1(n269), .A2(n268), .A3(n267), .Y(
        div_frac_add_in1_in[13]) );
  AOI22X1_RVT U400 ( .A1(div_frac_add_in1[13]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[15]), .Y(n272) );
  NAND2X0_RVT U401 ( .A1(n308), .A2(div_frac_outa[16]), .Y(n271) );
  NAND3X0_RVT U402 ( .A1(n272), .A2(n1), .A3(n271), .Y(div_frac_add_in1_in[14]) );
  AOI22X1_RVT U403 ( .A1(div_frac_add_in1[14]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[16]), .Y(n275) );
  NAND2X0_RVT U404 ( .A1(n308), .A2(div_frac_outa[17]), .Y(n274) );
  NAND3X0_RVT U405 ( .A1(n275), .A2(n2), .A3(n274), .Y(div_frac_add_in1_in[15]) );
  AOI22X1_RVT U406 ( .A1(div_frac_add_in1[15]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[17]), .Y(n278) );
  NAND2X0_RVT U407 ( .A1(n308), .A2(div_frac_outa[18]), .Y(n277) );
  NAND3X0_RVT U408 ( .A1(n278), .A2(n3), .A3(n277), .Y(div_frac_add_in1_in[16]) );
  AOI22X1_RVT U409 ( .A1(div_frac_add_in1[16]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[18]), .Y(n281) );
  NAND2X0_RVT U410 ( .A1(n308), .A2(div_frac_outa[19]), .Y(n280) );
  NAND3X0_RVT U411 ( .A1(n281), .A2(n4), .A3(n280), .Y(div_frac_add_in1_in[17]) );
  AOI22X1_RVT U412 ( .A1(div_frac_add_in1[17]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[19]), .Y(n284) );
  NAND2X0_RVT U413 ( .A1(n308), .A2(div_frac_outa[20]), .Y(n283) );
  NAND3X0_RVT U414 ( .A1(n284), .A2(n5), .A3(n283), .Y(div_frac_add_in1_in[18]) );
  AOI22X1_RVT U415 ( .A1(div_frac_add_in1[18]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[20]), .Y(n287) );
  NAND2X0_RVT U416 ( .A1(n308), .A2(div_frac_outa[21]), .Y(n286) );
  NAND3X0_RVT U417 ( .A1(n287), .A2(n6), .A3(n286), .Y(div_frac_add_in1_in[19]) );
  AOI22X1_RVT U418 ( .A1(div_frac_add_in1[19]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[21]), .Y(n290) );
  NAND2X0_RVT U419 ( .A1(n308), .A2(div_frac_outa[22]), .Y(n289) );
  NAND3X0_RVT U420 ( .A1(n290), .A2(n7), .A3(n289), .Y(div_frac_add_in1_in[20]) );
  AOI22X1_RVT U421 ( .A1(div_frac_add_in1[20]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[22]), .Y(n293) );
  NAND2X0_RVT U422 ( .A1(n308), .A2(div_frac_outa[23]), .Y(n292) );
  NAND3X0_RVT U423 ( .A1(n293), .A2(n8), .A3(n292), .Y(div_frac_add_in1_in[21]) );
  AOI22X1_RVT U424 ( .A1(div_frac_add_in1[21]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[23]), .Y(n296) );
  NAND2X0_RVT U425 ( .A1(n308), .A2(div_frac_outa[24]), .Y(n295) );
  NAND3X0_RVT U426 ( .A1(n296), .A2(n9), .A3(n295), .Y(div_frac_add_in1_in[22]) );
  AOI22X1_RVT U427 ( .A1(div_frac_add_in1[22]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[24]), .Y(n299) );
  NAND2X0_RVT U428 ( .A1(n308), .A2(div_frac_outa[25]), .Y(n298) );
  NAND3X0_RVT U429 ( .A1(n299), .A2(n10), .A3(n298), .Y(
        div_frac_add_in1_in[23]) );
  AOI22X1_RVT U430 ( .A1(div_frac_add_in1[23]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[25]), .Y(n302) );
  NAND2X0_RVT U431 ( .A1(n308), .A2(div_frac_outa[26]), .Y(n301) );
  NAND3X0_RVT U432 ( .A1(n302), .A2(n11), .A3(n301), .Y(
        div_frac_add_in1_in[24]) );
  AOI22X1_RVT U433 ( .A1(div_frac_add_in1[24]), .A2(n796), .A3(n306), .A4(
        div_frac_outa[26]), .Y(n305) );
  NAND2X0_RVT U434 ( .A1(n308), .A2(div_frac_outa[27]), .Y(n304) );
  NAND3X0_RVT U435 ( .A1(n305), .A2(n12), .A3(n304), .Y(
        div_frac_add_in1_in[25]) );
  AOI22X1_RVT U436 ( .A1(div_frac_add_in1[25]), .A2(n796), .A3(
        div_frac_outa[27]), .A4(n306), .Y(n310) );
  NAND2X0_RVT U437 ( .A1(div_frac_outa[28]), .A2(n308), .Y(n309) );
  NAND3X0_RVT U438 ( .A1(n310), .A2(n13), .A3(n309), .Y(
        div_frac_add_in1_in[26]) );
  AOI22X1_RVT U439 ( .A1(n396), .A2(div_frac_outa[32]), .A3(n395), .A4(
        div_frac_outa[31]), .Y(n314) );
  AOI22X1_RVT U440 ( .A1(d4stg_fdiv), .A2(div_shl_save[30]), .A3(
        div_frac_add_in1[29]), .A4(n796), .Y(n313) );
  FADDX1_RVT U441 ( .A(div_frac_add_in1a[29]), .B(div_frac_add_in2[29]), .CI(
        n311), .CO(n143), .S(n407) );
  NAND2X0_RVT U442 ( .A1(n795), .A2(n407), .Y(n312) );
  NAND3X0_RVT U443 ( .A1(n314), .A2(n313), .A3(n312), .Y(
        div_frac_add_in1_in[30]) );
  AOI22X1_RVT U444 ( .A1(n396), .A2(div_frac_outa[33]), .A3(n395), .A4(
        div_frac_outa[32]), .Y(n318) );
  AOI22X1_RVT U445 ( .A1(d4stg_fdiv), .A2(div_shl_save[31]), .A3(
        div_frac_add_in1[30]), .A4(n796), .Y(n317) );
  NAND2X0_RVT U446 ( .A1(n795), .A2(n315), .Y(n316) );
  NAND3X0_RVT U447 ( .A1(n318), .A2(n317), .A3(n316), .Y(
        div_frac_add_in1_in[31]) );
  AOI22X1_RVT U448 ( .A1(n396), .A2(div_frac_outa[34]), .A3(n395), .A4(
        div_frac_outa[33]), .Y(n322) );
  AOI22X1_RVT U449 ( .A1(d4stg_fdiv), .A2(div_shl_save[32]), .A3(
        div_frac_add_in1[31]), .A4(n796), .Y(n321) );
  NAND2X0_RVT U450 ( .A1(n795), .A2(n319), .Y(n320) );
  NAND3X0_RVT U451 ( .A1(n322), .A2(n321), .A3(n320), .Y(
        div_frac_add_in1_in[32]) );
  AOI22X1_RVT U452 ( .A1(n396), .A2(div_frac_outa[35]), .A3(n395), .A4(
        div_frac_outa[34]), .Y(n326) );
  AOI22X1_RVT U453 ( .A1(d4stg_fdiv), .A2(div_shl_save[33]), .A3(
        div_frac_add_in1[32]), .A4(n796), .Y(n325) );
  NAND2X0_RVT U454 ( .A1(n795), .A2(n323), .Y(n324) );
  NAND3X0_RVT U455 ( .A1(n326), .A2(n325), .A3(n324), .Y(
        div_frac_add_in1_in[33]) );
  AOI22X1_RVT U456 ( .A1(n396), .A2(div_frac_outa[36]), .A3(n395), .A4(
        div_frac_outa[35]), .Y(n330) );
  AOI22X1_RVT U457 ( .A1(d4stg_fdiv), .A2(div_shl_save[34]), .A3(
        div_frac_add_in1[33]), .A4(n796), .Y(n329) );
  NAND2X0_RVT U458 ( .A1(n795), .A2(n327), .Y(n328) );
  NAND3X0_RVT U459 ( .A1(n330), .A2(n329), .A3(n328), .Y(
        div_frac_add_in1_in[34]) );
  AOI22X1_RVT U460 ( .A1(n396), .A2(div_frac_outa[37]), .A3(n395), .A4(
        div_frac_outa[36]), .Y(n334) );
  AOI22X1_RVT U461 ( .A1(d4stg_fdiv), .A2(div_shl_save[35]), .A3(
        div_frac_add_in1[34]), .A4(n796), .Y(n333) );
  NAND2X0_RVT U462 ( .A1(n795), .A2(n331), .Y(n332) );
  NAND3X0_RVT U463 ( .A1(n334), .A2(n333), .A3(n332), .Y(
        div_frac_add_in1_in[35]) );
  AOI22X1_RVT U464 ( .A1(n396), .A2(div_frac_outa[38]), .A3(n395), .A4(
        div_frac_outa[37]), .Y(n338) );
  AOI22X1_RVT U465 ( .A1(d4stg_fdiv), .A2(div_shl_save[36]), .A3(
        div_frac_add_in1[35]), .A4(n796), .Y(n337) );
  NAND2X0_RVT U466 ( .A1(n795), .A2(n335), .Y(n336) );
  NAND3X0_RVT U467 ( .A1(n338), .A2(n337), .A3(n336), .Y(
        div_frac_add_in1_in[36]) );
  AOI22X1_RVT U468 ( .A1(n396), .A2(div_frac_outa[39]), .A3(n395), .A4(
        div_frac_outa[38]), .Y(n342) );
  AOI22X1_RVT U469 ( .A1(d4stg_fdiv), .A2(div_shl_save[37]), .A3(
        div_frac_add_in1[36]), .A4(n796), .Y(n341) );
  NAND2X0_RVT U470 ( .A1(n795), .A2(n339), .Y(n340) );
  NAND3X0_RVT U471 ( .A1(n342), .A2(n341), .A3(n340), .Y(
        div_frac_add_in1_in[37]) );
  AOI22X1_RVT U472 ( .A1(n396), .A2(div_frac_outa[40]), .A3(n395), .A4(
        div_frac_outa[39]), .Y(n346) );
  AOI22X1_RVT U473 ( .A1(d4stg_fdiv), .A2(div_shl_save[38]), .A3(
        div_frac_add_in1[37]), .A4(n796), .Y(n345) );
  NAND2X0_RVT U474 ( .A1(n795), .A2(n343), .Y(n344) );
  NAND3X0_RVT U475 ( .A1(n346), .A2(n345), .A3(n344), .Y(
        div_frac_add_in1_in[38]) );
  AOI22X1_RVT U476 ( .A1(n396), .A2(div_frac_outa[41]), .A3(n395), .A4(
        div_frac_outa[40]), .Y(n350) );
  AOI22X1_RVT U477 ( .A1(d4stg_fdiv), .A2(div_shl_save[39]), .A3(
        div_frac_add_in1[38]), .A4(n796), .Y(n349) );
  NAND2X0_RVT U478 ( .A1(n795), .A2(n347), .Y(n348) );
  NAND3X0_RVT U479 ( .A1(n350), .A2(n349), .A3(n348), .Y(
        div_frac_add_in1_in[39]) );
  AOI22X1_RVT U480 ( .A1(n396), .A2(div_frac_outa[42]), .A3(n395), .A4(
        div_frac_outa[41]), .Y(n354) );
  AOI22X1_RVT U481 ( .A1(d4stg_fdiv), .A2(div_shl_save[40]), .A3(
        div_frac_add_in1[39]), .A4(n796), .Y(n353) );
  NAND2X0_RVT U482 ( .A1(n795), .A2(n351), .Y(n352) );
  NAND3X0_RVT U483 ( .A1(n354), .A2(n353), .A3(n352), .Y(
        div_frac_add_in1_in[40]) );
  AOI22X1_RVT U484 ( .A1(n396), .A2(div_frac_outa[43]), .A3(n395), .A4(
        div_frac_outa[42]), .Y(n358) );
  AOI22X1_RVT U485 ( .A1(d4stg_fdiv), .A2(div_shl_save[41]), .A3(
        div_frac_add_in1[40]), .A4(n796), .Y(n357) );
  NAND2X0_RVT U486 ( .A1(n795), .A2(n355), .Y(n356) );
  NAND3X0_RVT U487 ( .A1(n358), .A2(n357), .A3(n356), .Y(
        div_frac_add_in1_in[41]) );
  AOI22X1_RVT U488 ( .A1(n396), .A2(div_frac_outa[44]), .A3(n395), .A4(
        div_frac_outa[43]), .Y(n362) );
  AOI22X1_RVT U489 ( .A1(d4stg_fdiv), .A2(div_shl_save[42]), .A3(
        div_frac_add_in1[41]), .A4(n796), .Y(n361) );
  NAND2X0_RVT U490 ( .A1(n795), .A2(n359), .Y(n360) );
  NAND3X0_RVT U491 ( .A1(n362), .A2(n361), .A3(n360), .Y(
        div_frac_add_in1_in[42]) );
  AOI22X1_RVT U492 ( .A1(n396), .A2(div_frac_outa[45]), .A3(n395), .A4(
        div_frac_outa[44]), .Y(n366) );
  AOI22X1_RVT U493 ( .A1(d4stg_fdiv), .A2(div_shl_save[43]), .A3(
        div_frac_add_in1[42]), .A4(n796), .Y(n365) );
  NAND2X0_RVT U494 ( .A1(n795), .A2(n363), .Y(n364) );
  NAND3X0_RVT U495 ( .A1(n366), .A2(n365), .A3(n364), .Y(
        div_frac_add_in1_in[43]) );
  AOI22X1_RVT U496 ( .A1(n396), .A2(div_frac_outa[46]), .A3(n395), .A4(
        div_frac_outa[45]), .Y(n370) );
  AOI22X1_RVT U497 ( .A1(d4stg_fdiv), .A2(div_shl_save[44]), .A3(
        div_frac_add_in1[43]), .A4(n796), .Y(n369) );
  NAND2X0_RVT U498 ( .A1(n795), .A2(n367), .Y(n368) );
  NAND3X0_RVT U499 ( .A1(n370), .A2(n369), .A3(n368), .Y(
        div_frac_add_in1_in[44]) );
  AOI22X1_RVT U500 ( .A1(n396), .A2(div_frac_outa[47]), .A3(n395), .A4(
        div_frac_outa[46]), .Y(n374) );
  AOI22X1_RVT U501 ( .A1(d4stg_fdiv), .A2(div_shl_save[45]), .A3(
        div_frac_add_in1[44]), .A4(n796), .Y(n373) );
  NAND2X0_RVT U502 ( .A1(n795), .A2(n371), .Y(n372) );
  NAND3X0_RVT U503 ( .A1(n374), .A2(n373), .A3(n372), .Y(
        div_frac_add_in1_in[45]) );
  AOI22X1_RVT U504 ( .A1(n396), .A2(div_frac_outa[48]), .A3(n395), .A4(
        div_frac_outa[47]), .Y(n378) );
  AOI22X1_RVT U505 ( .A1(d4stg_fdiv), .A2(div_shl_save[46]), .A3(
        div_frac_add_in1[45]), .A4(n796), .Y(n377) );
  NAND2X0_RVT U506 ( .A1(n795), .A2(n375), .Y(n376) );
  NAND3X0_RVT U507 ( .A1(n378), .A2(n377), .A3(n376), .Y(
        div_frac_add_in1_in[46]) );
  AOI22X1_RVT U508 ( .A1(n396), .A2(div_frac_outa[49]), .A3(n395), .A4(
        div_frac_outa[48]), .Y(n382) );
  AOI22X1_RVT U509 ( .A1(d4stg_fdiv), .A2(div_shl_save[47]), .A3(
        div_frac_add_in1[46]), .A4(n796), .Y(n381) );
  NAND2X0_RVT U510 ( .A1(n795), .A2(n379), .Y(n380) );
  NAND3X0_RVT U511 ( .A1(n382), .A2(n381), .A3(n380), .Y(
        div_frac_add_in1_in[47]) );
  AOI22X1_RVT U512 ( .A1(n396), .A2(div_frac_outa[50]), .A3(n395), .A4(
        div_frac_outa[49]), .Y(n386) );
  AOI22X1_RVT U513 ( .A1(d4stg_fdiv), .A2(div_shl_save[48]), .A3(
        div_frac_add_in1[47]), .A4(n796), .Y(n385) );
  NAND2X0_RVT U514 ( .A1(n795), .A2(n383), .Y(n384) );
  NAND3X0_RVT U515 ( .A1(n386), .A2(n385), .A3(n384), .Y(
        div_frac_add_in1_in[48]) );
  AOI22X1_RVT U516 ( .A1(n396), .A2(div_frac_outa[51]), .A3(n395), .A4(
        div_frac_outa[50]), .Y(n390) );
  AOI22X1_RVT U517 ( .A1(d4stg_fdiv), .A2(div_shl_save[49]), .A3(
        div_frac_add_in1[48]), .A4(n796), .Y(n389) );
  NAND2X0_RVT U518 ( .A1(n795), .A2(n387), .Y(n388) );
  NAND3X0_RVT U519 ( .A1(n390), .A2(n389), .A3(n388), .Y(
        div_frac_add_in1_in[49]) );
  AOI22X1_RVT U520 ( .A1(n396), .A2(\div_frac_out[52] ), .A3(n395), .A4(
        div_frac_outa[51]), .Y(n394) );
  AOI22X1_RVT U521 ( .A1(d4stg_fdiv), .A2(div_shl_save[50]), .A3(
        div_frac_add_in1[49]), .A4(n796), .Y(n393) );
  NAND2X0_RVT U522 ( .A1(n795), .A2(n391), .Y(n392) );
  NAND3X0_RVT U523 ( .A1(n394), .A2(n393), .A3(n392), .Y(
        div_frac_add_in1_in[50]) );
  AOI22X1_RVT U524 ( .A1(div_frac_out_54_53[0]), .A2(n396), .A3(
        \div_frac_out[52] ), .A4(n395), .Y(n400) );
  AOI22X1_RVT U525 ( .A1(d4stg_fdiv), .A2(div_shl_save[51]), .A3(
        div_frac_add_in1[50]), .A4(n796), .Y(n399) );
  NAND2X0_RVT U526 ( .A1(n795), .A2(n397), .Y(n398) );
  NAND3X0_RVT U527 ( .A1(n400), .A2(n399), .A3(n398), .Y(
        div_frac_add_in1_in[51]) );
  AO22X1_RVT U528 ( .A1(div_frac_add_in1[52]), .A2(n796), .A3(n795), .A4(n401), 
        .Y(div_frac_add_in1_in[53]) );
  AO22X1_RVT U529 ( .A1(div_frac_add_in1[53]), .A2(n796), .A3(n795), .A4(n402), 
        .Y(div_frac_add_in1_in[54]) );
  AOI22X1_RVT U530 ( .A1(div_frac_out_shl1_dbl), .A2(div_frac_outa[28]), .A3(
        div_frac_out_shl1_sng), .A4(n403), .Y(n405) );
  NAND2X0_RVT U531 ( .A1(div_frac_add_in1[29]), .A2(div_frac_out_add_in1), .Y(
        n404) );
  NAND3X0_RVT U532 ( .A1(n405), .A2(n14), .A3(n404), .Y(n406) );
  AO21X1_RVT U533 ( .A1(n407), .A2(div_frac_out_add), .A3(n406), .Y(
        div_frac_out_in[29]) );
  AO22X1_RVT U534 ( .A1(n408), .A2(div_shl_data[4]), .A3(n425), .A4(
        div_shl_data[3]), .Y(n410) );
  AO22X1_RVT U535 ( .A1(div_shl_data[1]), .A2(n22), .A3(n506), .A4(
        div_shl_data[2]), .Y(n409) );
  OR2X1_RVT U536 ( .A1(n410), .A2(n409), .Y(n519) );
  OA222X1_RVT U537 ( .A1(n521), .A2(n408), .A3(n521), .A4(div_shl_data[0]), 
        .A5(div_shl_cnta[2]), .A6(n519), .Y(n551) );
  AND2X1_RVT U538 ( .A1(n551), .A2(n779), .Y(n781) );
  AO22X1_RVT U539 ( .A1(n408), .A2(div_shl_data[16]), .A3(n425), .A4(
        div_shl_data[15]), .Y(n412) );
  AO22X1_RVT U540 ( .A1(n22), .A2(div_shl_data[13]), .A3(n506), .A4(
        div_shl_data[14]), .Y(n411) );
  OR2X1_RVT U541 ( .A1(n412), .A2(n411), .Y(n547) );
  AO22X1_RVT U542 ( .A1(n408), .A2(div_shl_data[20]), .A3(n425), .A4(
        div_shl_data[19]), .Y(n414) );
  AO22X1_RVT U543 ( .A1(n22), .A2(div_shl_data[17]), .A3(n506), .A4(
        div_shl_data[18]), .Y(n413) );
  OR2X1_RVT U544 ( .A1(n414), .A2(n413), .Y(n601) );
  AO22X1_RVT U545 ( .A1(n408), .A2(div_shl_data[8]), .A3(n425), .A4(
        div_shl_data[7]), .Y(n416) );
  AO22X1_RVT U546 ( .A1(n22), .A2(div_shl_data[5]), .A3(n506), .A4(
        div_shl_data[6]), .Y(n415) );
  OR2X1_RVT U547 ( .A1(n416), .A2(n415), .Y(n518) );
  AO22X1_RVT U548 ( .A1(n408), .A2(div_shl_data[12]), .A3(n425), .A4(
        div_shl_data[11]), .Y(n418) );
  AO22X1_RVT U549 ( .A1(n22), .A2(div_shl_data[9]), .A3(n506), .A4(
        div_shl_data[10]), .Y(n417) );
  OR2X1_RVT U550 ( .A1(n418), .A2(n417), .Y(n520) );
  AO22X1_RVT U551 ( .A1(div_shl_cnta[2]), .A2(n518), .A3(n521), .A4(n520), .Y(
        n550) );
  AO222X1_RVT U552 ( .A1(n547), .A2(n715), .A3(n601), .A4(n21), .A5(n550), 
        .A6(div_shl_cnta[3]), .Y(n723) );
  AO22X1_RVT U553 ( .A1(div_shl_cnta[4]), .A2(n781), .A3(n774), .A4(n723), .Y(
        n762) );
  AO22X1_RVT U554 ( .A1(n408), .A2(div_shl_data[32]), .A3(n425), .A4(
        div_shl_data[31]), .Y(n420) );
  AO22X1_RVT U555 ( .A1(n22), .A2(div_shl_data[29]), .A3(n506), .A4(
        div_shl_data[30]), .Y(n419) );
  NOR2X0_RVT U556 ( .A1(n420), .A2(n419), .Y(n600) );
  AO22X1_RVT U557 ( .A1(n408), .A2(div_shl_data[36]), .A3(n425), .A4(
        div_shl_data[35]), .Y(n422) );
  AO22X1_RVT U558 ( .A1(n22), .A2(div_shl_data[33]), .A3(n506), .A4(
        div_shl_data[34]), .Y(n421) );
  NOR2X0_RVT U559 ( .A1(n422), .A2(n421), .Y(n597) );
  OA22X1_RVT U560 ( .A1(n600), .A2(n604), .A3(n597), .A4(n710), .Y(n429) );
  AO22X1_RVT U561 ( .A1(n408), .A2(div_shl_data[24]), .A3(n425), .A4(
        div_shl_data[23]), .Y(n424) );
  AO22X1_RVT U562 ( .A1(n22), .A2(div_shl_data[21]), .A3(n506), .A4(
        div_shl_data[22]), .Y(n423) );
  NOR2X0_RVT U563 ( .A1(n424), .A2(n423), .Y(n602) );
  AO22X1_RVT U564 ( .A1(n408), .A2(div_shl_data[28]), .A3(n425), .A4(
        div_shl_data[27]), .Y(n427) );
  AO22X1_RVT U565 ( .A1(n22), .A2(div_shl_data[25]), .A3(n506), .A4(
        div_shl_data[26]), .Y(n426) );
  NOR2X0_RVT U566 ( .A1(n427), .A2(n426), .Y(n599) );
  OA22X1_RVT U567 ( .A1(n602), .A2(n537), .A3(n599), .A4(n34), .Y(n428) );
  NAND2X0_RVT U568 ( .A1(n429), .A2(n428), .Y(n724) );
  AO22X1_RVT U569 ( .A1(n408), .A2(div_shl_data[40]), .A3(n425), .A4(
        div_shl_data[39]), .Y(n431) );
  AO22X1_RVT U570 ( .A1(n22), .A2(div_shl_data[37]), .A3(n506), .A4(
        div_shl_data[38]), .Y(n430) );
  OR2X1_RVT U571 ( .A1(n431), .A2(n430), .Y(n543) );
  AO22X1_RVT U572 ( .A1(n408), .A2(div_shl_data[44]), .A3(n425), .A4(
        div_shl_data[43]), .Y(n433) );
  AO22X1_RVT U573 ( .A1(n22), .A2(div_shl_data[41]), .A3(n506), .A4(
        div_shl_data[42]), .Y(n432) );
  OR2X1_RVT U574 ( .A1(n433), .A2(n432), .Y(n544) );
  AO22X1_RVT U575 ( .A1(n408), .A2(div_shl_data[48]), .A3(n425), .A4(
        div_shl_data[47]), .Y(n435) );
  AO22X1_RVT U576 ( .A1(n22), .A2(div_shl_data[45]), .A3(n506), .A4(
        div_shl_data[46]), .Y(n434) );
  OR2X1_RVT U577 ( .A1(n435), .A2(n434), .Y(n512) );
  AO222X1_RVT U578 ( .A1(n543), .A2(n708), .A3(n544), .A4(n592), .A5(n512), 
        .A6(n715), .Y(n439) );
  AO22X1_RVT U579 ( .A1(n408), .A2(div_shl_data[52]), .A3(n425), .A4(
        div_shl_data[51]), .Y(n437) );
  AO22X1_RVT U580 ( .A1(n22), .A2(div_shl_data[49]), .A3(n506), .A4(
        div_shl_data[50]), .Y(n436) );
  AND2X1_RVT U581 ( .A1(n21), .A2(n774), .Y(n725) );
  OA21X1_RVT U582 ( .A1(n437), .A2(n436), .A3(n725), .Y(n438) );
  AO221X1_RVT U583 ( .A1(div_shl_cnta[4]), .A2(n724), .A3(n774), .A4(n439), 
        .A5(n438), .Y(n440) );
  AO22X1_RVT U584 ( .A1(div_shl_cnta[5]), .A2(n762), .A3(n775), .A4(n440), .Y(
        div_shl_tmp[105]) );
  NOR2X0_RVT U585 ( .A1(div_shl_tmp[105]), .A2(n761), .Y(
        div_frac_add_in2_in[52]) );
  AND2X1_RVT U586 ( .A1(div_shl_cnta[4]), .A2(n21), .Y(n502) );
  AO22X1_RVT U587 ( .A1(n408), .A2(div_shl_data[3]), .A3(div_shl_data[2]), 
        .A4(n425), .Y(n442) );
  AO22X1_RVT U588 ( .A1(div_shl_data[0]), .A2(n22), .A3(div_shl_data[1]), .A4(
        n506), .Y(n441) );
  OR2X1_RVT U589 ( .A1(n442), .A2(n441), .Y(n782) );
  AO22X1_RVT U590 ( .A1(n408), .A2(div_shl_data[15]), .A3(n425), .A4(
        div_shl_data[14]), .Y(n444) );
  AO22X1_RVT U591 ( .A1(n22), .A2(div_shl_data[12]), .A3(n506), .A4(
        div_shl_data[13]), .Y(n443) );
  OR2X1_RVT U592 ( .A1(n444), .A2(n443), .Y(n618) );
  AO22X1_RVT U593 ( .A1(n408), .A2(div_shl_data[19]), .A3(n425), .A4(
        div_shl_data[18]), .Y(n446) );
  AO22X1_RVT U594 ( .A1(n22), .A2(div_shl_data[16]), .A3(n506), .A4(
        div_shl_data[17]), .Y(n445) );
  OR2X1_RVT U595 ( .A1(n446), .A2(n445), .Y(n623) );
  AO22X1_RVT U596 ( .A1(n408), .A2(div_shl_data[7]), .A3(n425), .A4(
        div_shl_data[6]), .Y(n448) );
  AO22X1_RVT U597 ( .A1(n22), .A2(div_shl_data[4]), .A3(n506), .A4(
        div_shl_data[5]), .Y(n447) );
  OR2X1_RVT U598 ( .A1(n448), .A2(n447), .Y(n616) );
  AO22X1_RVT U599 ( .A1(n408), .A2(div_shl_data[11]), .A3(n425), .A4(
        div_shl_data[10]), .Y(n450) );
  AO22X1_RVT U600 ( .A1(n22), .A2(div_shl_data[8]), .A3(n506), .A4(
        div_shl_data[9]), .Y(n449) );
  OR2X1_RVT U601 ( .A1(n450), .A2(n449), .Y(n617) );
  AO22X1_RVT U602 ( .A1(div_shl_cnta[2]), .A2(n616), .A3(n521), .A4(n617), .Y(
        n564) );
  AO222X1_RVT U603 ( .A1(n618), .A2(n715), .A3(n623), .A4(n21), .A5(n564), 
        .A6(div_shl_cnta[3]), .Y(n727) );
  AO22X1_RVT U604 ( .A1(n502), .A2(n782), .A3(n774), .A4(n727), .Y(n763) );
  AO22X1_RVT U605 ( .A1(n408), .A2(div_shl_data[31]), .A3(n425), .A4(
        div_shl_data[30]), .Y(n452) );
  AO22X1_RVT U606 ( .A1(n22), .A2(div_shl_data[28]), .A3(n506), .A4(
        div_shl_data[29]), .Y(n451) );
  NOR2X0_RVT U607 ( .A1(n452), .A2(n451), .Y(n613) );
  AO22X1_RVT U608 ( .A1(n408), .A2(div_shl_data[35]), .A3(n425), .A4(
        div_shl_data[34]), .Y(n454) );
  AO22X1_RVT U609 ( .A1(n22), .A2(div_shl_data[32]), .A3(n506), .A4(
        div_shl_data[33]), .Y(n453) );
  NOR2X0_RVT U610 ( .A1(n454), .A2(n453), .Y(n614) );
  OA22X1_RVT U611 ( .A1(n613), .A2(n604), .A3(n614), .A4(n710), .Y(n460) );
  AO22X1_RVT U612 ( .A1(n408), .A2(div_shl_data[23]), .A3(n425), .A4(
        div_shl_data[22]), .Y(n456) );
  AO22X1_RVT U613 ( .A1(n22), .A2(div_shl_data[20]), .A3(n506), .A4(
        div_shl_data[21]), .Y(n455) );
  NOR2X0_RVT U614 ( .A1(n456), .A2(n455), .Y(n619) );
  AO22X1_RVT U615 ( .A1(n408), .A2(div_shl_data[27]), .A3(n425), .A4(
        div_shl_data[26]), .Y(n458) );
  AO22X1_RVT U616 ( .A1(n22), .A2(div_shl_data[24]), .A3(n506), .A4(
        div_shl_data[25]), .Y(n457) );
  NOR2X0_RVT U617 ( .A1(n458), .A2(n457), .Y(n612) );
  OA22X1_RVT U618 ( .A1(n619), .A2(n537), .A3(n612), .A4(n34), .Y(n459) );
  NAND2X0_RVT U619 ( .A1(n460), .A2(n459), .Y(n726) );
  AO22X1_RVT U620 ( .A1(n408), .A2(div_shl_data[39]), .A3(n425), .A4(
        div_shl_data[38]), .Y(n462) );
  AO22X1_RVT U621 ( .A1(n22), .A2(div_shl_data[36]), .A3(n506), .A4(
        div_shl_data[37]), .Y(n461) );
  OR2X1_RVT U622 ( .A1(n462), .A2(n461), .Y(n556) );
  AO22X1_RVT U623 ( .A1(n408), .A2(div_shl_data[43]), .A3(n425), .A4(
        div_shl_data[42]), .Y(n464) );
  AO22X1_RVT U624 ( .A1(n22), .A2(div_shl_data[40]), .A3(n506), .A4(
        div_shl_data[41]), .Y(n463) );
  OR2X1_RVT U625 ( .A1(n464), .A2(n463), .Y(n557) );
  AO22X1_RVT U626 ( .A1(n408), .A2(div_shl_data[47]), .A3(n425), .A4(
        div_shl_data[46]), .Y(n466) );
  AO22X1_RVT U627 ( .A1(n22), .A2(div_shl_data[44]), .A3(n506), .A4(
        div_shl_data[45]), .Y(n465) );
  OR2X1_RVT U628 ( .A1(n466), .A2(n465), .Y(n526) );
  AO222X1_RVT U629 ( .A1(n556), .A2(n708), .A3(n557), .A4(n592), .A5(n526), 
        .A6(n715), .Y(n470) );
  AO22X1_RVT U630 ( .A1(n408), .A2(div_shl_data[51]), .A3(n425), .A4(
        div_shl_data[50]), .Y(n468) );
  AO22X1_RVT U631 ( .A1(n22), .A2(div_shl_data[48]), .A3(n506), .A4(
        div_shl_data[49]), .Y(n467) );
  OA21X1_RVT U632 ( .A1(n468), .A2(n467), .A3(n725), .Y(n469) );
  AO221X1_RVT U633 ( .A1(div_shl_cnta[4]), .A2(n726), .A3(n774), .A4(n470), 
        .A5(n469), .Y(n471) );
  AO22X1_RVT U634 ( .A1(div_shl_cnta[5]), .A2(n763), .A3(n775), .A4(n471), .Y(
        div_shl_tmp[104]) );
  NOR2X0_RVT U635 ( .A1(div_shl_tmp[104]), .A2(n761), .Y(
        div_frac_add_in2_in[51]) );
  AO222X1_RVT U636 ( .A1(n408), .A2(div_shl_data[2]), .A3(div_shl_data[1]), 
        .A4(n425), .A5(div_shl_data[0]), .A6(n506), .Y(n783) );
  AO22X1_RVT U637 ( .A1(n408), .A2(div_shl_data[14]), .A3(n425), .A4(
        div_shl_data[13]), .Y(n473) );
  AO22X1_RVT U638 ( .A1(n22), .A2(div_shl_data[11]), .A3(n506), .A4(
        div_shl_data[12]), .Y(n472) );
  OR2X1_RVT U639 ( .A1(n473), .A2(n472), .Y(n635) );
  AO22X1_RVT U640 ( .A1(n408), .A2(div_shl_data[18]), .A3(n425), .A4(
        div_shl_data[17]), .Y(n475) );
  AO22X1_RVT U641 ( .A1(n22), .A2(div_shl_data[15]), .A3(n506), .A4(
        div_shl_data[16]), .Y(n474) );
  OR2X1_RVT U642 ( .A1(n475), .A2(n474), .Y(n640) );
  AO22X1_RVT U643 ( .A1(n408), .A2(div_shl_data[6]), .A3(n425), .A4(
        div_shl_data[5]), .Y(n477) );
  AO22X1_RVT U644 ( .A1(n22), .A2(div_shl_data[3]), .A3(n506), .A4(
        div_shl_data[4]), .Y(n476) );
  OR2X1_RVT U645 ( .A1(n477), .A2(n476), .Y(n633) );
  AO22X1_RVT U646 ( .A1(n408), .A2(div_shl_data[10]), .A3(n425), .A4(
        div_shl_data[9]), .Y(n479) );
  AO22X1_RVT U647 ( .A1(n22), .A2(div_shl_data[7]), .A3(n506), .A4(
        div_shl_data[8]), .Y(n478) );
  OR2X1_RVT U648 ( .A1(n479), .A2(n478), .Y(n634) );
  AO22X1_RVT U649 ( .A1(div_shl_cnta[2]), .A2(n633), .A3(n521), .A4(n634), .Y(
        n577) );
  AO222X1_RVT U650 ( .A1(n635), .A2(n715), .A3(n640), .A4(n21), .A5(n577), 
        .A6(div_shl_cnta[3]), .Y(n729) );
  AO22X1_RVT U651 ( .A1(n502), .A2(n783), .A3(n774), .A4(n729), .Y(n764) );
  AO22X1_RVT U652 ( .A1(n408), .A2(div_shl_data[30]), .A3(n425), .A4(
        div_shl_data[29]), .Y(n481) );
  AO22X1_RVT U653 ( .A1(n22), .A2(div_shl_data[27]), .A3(n506), .A4(
        div_shl_data[28]), .Y(n480) );
  NOR2X0_RVT U654 ( .A1(n481), .A2(n480), .Y(n630) );
  AO22X1_RVT U655 ( .A1(n408), .A2(div_shl_data[34]), .A3(n425), .A4(
        div_shl_data[33]), .Y(n483) );
  AO22X1_RVT U656 ( .A1(n22), .A2(div_shl_data[31]), .A3(n506), .A4(
        div_shl_data[32]), .Y(n482) );
  NOR2X0_RVT U657 ( .A1(n483), .A2(n482), .Y(n631) );
  OA22X1_RVT U658 ( .A1(n630), .A2(n604), .A3(n631), .A4(n710), .Y(n489) );
  AO22X1_RVT U659 ( .A1(n408), .A2(div_shl_data[22]), .A3(n425), .A4(
        div_shl_data[21]), .Y(n485) );
  AO22X1_RVT U660 ( .A1(n22), .A2(div_shl_data[19]), .A3(n506), .A4(
        div_shl_data[20]), .Y(n484) );
  NOR2X0_RVT U661 ( .A1(n485), .A2(n484), .Y(n636) );
  AO22X1_RVT U662 ( .A1(n408), .A2(div_shl_data[26]), .A3(n425), .A4(
        div_shl_data[25]), .Y(n487) );
  AO22X1_RVT U663 ( .A1(n22), .A2(div_shl_data[23]), .A3(n506), .A4(
        div_shl_data[24]), .Y(n486) );
  NOR2X0_RVT U664 ( .A1(n487), .A2(n486), .Y(n629) );
  OA22X1_RVT U665 ( .A1(n636), .A2(n537), .A3(n629), .A4(n34), .Y(n488) );
  NAND2X0_RVT U666 ( .A1(n489), .A2(n488), .Y(n728) );
  AO22X1_RVT U667 ( .A1(n408), .A2(div_shl_data[38]), .A3(n425), .A4(
        div_shl_data[37]), .Y(n491) );
  AO22X1_RVT U668 ( .A1(n22), .A2(div_shl_data[35]), .A3(n506), .A4(
        div_shl_data[36]), .Y(n490) );
  OR2X1_RVT U669 ( .A1(n491), .A2(n490), .Y(n569) );
  AO22X1_RVT U670 ( .A1(n408), .A2(div_shl_data[42]), .A3(n425), .A4(
        div_shl_data[41]), .Y(n493) );
  AO22X1_RVT U671 ( .A1(n22), .A2(div_shl_data[39]), .A3(n506), .A4(
        div_shl_data[40]), .Y(n492) );
  OR2X1_RVT U672 ( .A1(n493), .A2(n492), .Y(n570) );
  AO22X1_RVT U673 ( .A1(n408), .A2(div_shl_data[46]), .A3(n425), .A4(
        div_shl_data[45]), .Y(n495) );
  AO22X1_RVT U674 ( .A1(n22), .A2(div_shl_data[43]), .A3(n506), .A4(
        div_shl_data[44]), .Y(n494) );
  OR2X1_RVT U675 ( .A1(n495), .A2(n494), .Y(n534) );
  AO222X1_RVT U676 ( .A1(n569), .A2(n708), .A3(n570), .A4(n592), .A5(n534), 
        .A6(n715), .Y(n499) );
  AO22X1_RVT U677 ( .A1(n408), .A2(div_shl_data[50]), .A3(n425), .A4(
        div_shl_data[49]), .Y(n497) );
  AO22X1_RVT U678 ( .A1(n22), .A2(div_shl_data[47]), .A3(n506), .A4(
        div_shl_data[48]), .Y(n496) );
  OA21X1_RVT U679 ( .A1(n497), .A2(n496), .A3(n725), .Y(n498) );
  AO221X1_RVT U680 ( .A1(div_shl_cnta[4]), .A2(n728), .A3(n774), .A4(n499), 
        .A5(n498), .Y(n500) );
  AO22X1_RVT U681 ( .A1(div_shl_cnta[5]), .A2(n764), .A3(n775), .A4(n500), .Y(
        div_shl_tmp[103]) );
  NOR2X0_RVT U682 ( .A1(div_shl_tmp[103]), .A2(n761), .Y(
        div_frac_add_in2_in[50]) );
  AO22X1_RVT U683 ( .A1(div_shl_cnta[2]), .A2(n501), .A3(n521), .A4(n707), .Y(
        n591) );
  AO222X1_RVT U684 ( .A1(n709), .A2(n715), .A3(n716), .A4(n21), .A5(n591), 
        .A6(div_shl_cnta[3]), .Y(n731) );
  AO22X1_RVT U685 ( .A1(n502), .A2(n784), .A3(n774), .A4(n731), .Y(n765) );
  OA22X1_RVT U686 ( .A1(n649), .A2(n604), .A3(n704), .A4(n710), .Y(n504) );
  OA22X1_RVT U687 ( .A1(n711), .A2(n537), .A3(n647), .A4(n34), .Y(n503) );
  NAND2X0_RVT U688 ( .A1(n504), .A2(n503), .Y(n730) );
  AO222X1_RVT U689 ( .A1(n582), .A2(n708), .A3(n584), .A4(n592), .A5(n505), 
        .A6(n715), .Y(n510) );
  AO22X1_RVT U690 ( .A1(n408), .A2(div_shl_data[49]), .A3(n425), .A4(
        div_shl_data[48]), .Y(n508) );
  AO22X1_RVT U691 ( .A1(n22), .A2(div_shl_data[46]), .A3(n506), .A4(
        div_shl_data[47]), .Y(n507) );
  OA21X1_RVT U692 ( .A1(n508), .A2(n507), .A3(n725), .Y(n509) );
  AO221X1_RVT U693 ( .A1(div_shl_cnta[4]), .A2(n730), .A3(n774), .A4(n510), 
        .A5(n509), .Y(n511) );
  AO22X1_RVT U694 ( .A1(div_shl_cnta[5]), .A2(n765), .A3(n775), .A4(n511), .Y(
        div_shl_tmp[102]) );
  NOR2X0_RVT U695 ( .A1(div_shl_tmp[102]), .A2(n761), .Y(
        div_frac_add_in2_in[49]) );
  AOI22X1_RVT U697 ( .A1(n583), .A2(n544), .A3(n785), .A4(n512), .Y(n525) );
  INVX1_RVT U698 ( .A(n543), .Y(n598) );
  OA22X1_RVT U699 ( .A1(n598), .A2(n648), .A3(n597), .A4(n646), .Y(n524) );
  NAND2X0_RVT U700 ( .A1(n708), .A2(n601), .Y(n514) );
  OA22X1_RVT U701 ( .A1(n602), .A2(n34), .A3(n600), .A4(n710), .Y(n513) );
  AND2X1_RVT U702 ( .A1(n514), .A2(n513), .Y(n517) );
  NAND2X0_RVT U703 ( .A1(n515), .A2(n715), .Y(n516) );
  AND2X1_RVT U704 ( .A1(n517), .A2(n516), .Y(n734) );
  NAND4X0_RVT U705 ( .A1(n408), .A2(div_shl_data[0]), .A3(n779), .A4(n521), 
        .Y(n735) );
  AO22X1_RVT U706 ( .A1(div_shl_cnta[2]), .A2(n519), .A3(n521), .A4(n518), .Y(
        n606) );
  OAI22X1_RVT U707 ( .A1(n521), .A2(n520), .A3(div_shl_cnta[2]), .A4(n547), 
        .Y(n605) );
  AO22X1_RVT U708 ( .A1(div_shl_cnta[3]), .A2(n522), .A3(n779), .A4(n605), .Y(
        n733) );
  AO22X1_RVT U709 ( .A1(div_shl_cnta[4]), .A2(n735), .A3(n774), .A4(n733), .Y(
        n766) );
  OA22X1_RVT U710 ( .A1(n734), .A2(n758), .A3(n775), .A4(n766), .Y(n523) );
  NAND3X0_RVT U711 ( .A1(n525), .A2(n524), .A3(n523), .Y(div_shl_tmp[101]) );
  INVX1_RVT U712 ( .A(d4stg_fdiv), .Y(n761) );
  NOR2X0_RVT U713 ( .A1(n761), .A2(div_shl_tmp[101]), .Y(
        div_frac_add_in2_in[48]) );
  INVX1_RVT U714 ( .A(n556), .Y(n615) );
  OA22X1_RVT U715 ( .A1(n615), .A2(n648), .A3(n614), .A4(n646), .Y(n533) );
  AOI22X1_RVT U716 ( .A1(n583), .A2(n557), .A3(n785), .A4(n526), .Y(n532) );
  AO22X1_RVT U717 ( .A1(n715), .A2(n617), .A3(n21), .A4(n618), .Y(n528) );
  AO22X1_RVT U718 ( .A1(n708), .A2(n782), .A3(n592), .A4(n616), .Y(n527) );
  OR2X1_RVT U719 ( .A1(n528), .A2(n527), .Y(n767) );
  INVX1_RVT U720 ( .A(n767), .Y(n738) );
  OA22X1_RVT U721 ( .A1(n612), .A2(n604), .A3(n613), .A4(n710), .Y(n530) );
  OA22X1_RVT U722 ( .A1(n558), .A2(n537), .A3(n619), .A4(n34), .Y(n529) );
  AND2X1_RVT U723 ( .A1(n530), .A2(n529), .Y(n737) );
  OA22X1_RVT U724 ( .A1(n738), .A2(n736), .A3(n737), .A4(n758), .Y(n531) );
  NAND3X0_RVT U725 ( .A1(n533), .A2(n532), .A3(n531), .Y(div_shl_tmp[100]) );
  NOR2X0_RVT U726 ( .A1(n761), .A2(div_shl_tmp[100]), .Y(
        div_frac_add_in2_in[47]) );
  INVX1_RVT U727 ( .A(n569), .Y(n632) );
  OA22X1_RVT U728 ( .A1(n632), .A2(n648), .A3(n631), .A4(n646), .Y(n542) );
  AOI22X1_RVT U729 ( .A1(n583), .A2(n570), .A3(n785), .A4(n534), .Y(n541) );
  AO22X1_RVT U730 ( .A1(n715), .A2(n634), .A3(n21), .A4(n635), .Y(n536) );
  AO22X1_RVT U731 ( .A1(n708), .A2(n783), .A3(n592), .A4(n633), .Y(n535) );
  OR2X1_RVT U732 ( .A1(n536), .A2(n535), .Y(n768) );
  INVX1_RVT U733 ( .A(n768), .Y(n740) );
  OA22X1_RVT U734 ( .A1(n629), .A2(n604), .A3(n630), .A4(n710), .Y(n539) );
  OA22X1_RVT U735 ( .A1(n571), .A2(n537), .A3(n636), .A4(n34), .Y(n538) );
  AND2X1_RVT U736 ( .A1(n539), .A2(n538), .Y(n739) );
  OA22X1_RVT U737 ( .A1(n740), .A2(n736), .A3(n739), .A4(n758), .Y(n540) );
  NAND3X0_RVT U738 ( .A1(n542), .A2(n541), .A3(n540), .Y(div_shl_tmp[99]) );
  NOR2X0_RVT U739 ( .A1(n761), .A2(div_shl_tmp[99]), .Y(
        div_frac_add_in2_in[46]) );
  NOR2X0_RVT U740 ( .A1(n761), .A2(div_shl_tmp[98]), .Y(
        div_frac_add_in2_in[45]) );
  AOI22X1_RVT U741 ( .A1(n785), .A2(n544), .A3(n583), .A4(n543), .Y(n555) );
  OA22X1_RVT U742 ( .A1(n597), .A2(n648), .A3(n600), .A4(n646), .Y(n554) );
  NAND2X0_RVT U743 ( .A1(n592), .A2(n601), .Y(n546) );
  OA22X1_RVT U744 ( .A1(n602), .A2(n604), .A3(n599), .A4(n710), .Y(n545) );
  AND2X1_RVT U745 ( .A1(n546), .A2(n545), .Y(n549) );
  NAND2X0_RVT U746 ( .A1(n547), .A2(n708), .Y(n548) );
  AND2X1_RVT U747 ( .A1(n549), .A2(n548), .Y(n742) );
  AO22X1_RVT U748 ( .A1(div_shl_cnta[3]), .A2(n551), .A3(n779), .A4(n550), .Y(
        n770) );
  NAND2X0_RVT U749 ( .A1(n770), .A2(n774), .Y(n552) );
  OA22X1_RVT U750 ( .A1(n742), .A2(n758), .A3(n775), .A4(n552), .Y(n553) );
  NAND3X0_RVT U751 ( .A1(n555), .A2(n554), .A3(n553), .Y(div_shl_tmp[97]) );
  NOR2X0_RVT U752 ( .A1(n761), .A2(div_shl_tmp[97]), .Y(
        div_frac_add_in2_in[44]) );
  OA22X1_RVT U753 ( .A1(n614), .A2(n648), .A3(n613), .A4(n646), .Y(n568) );
  AOI22X1_RVT U754 ( .A1(n785), .A2(n557), .A3(n583), .A4(n556), .Y(n567) );
  NAND2X0_RVT U755 ( .A1(n708), .A2(n618), .Y(n560) );
  OA22X1_RVT U756 ( .A1(n558), .A2(n34), .A3(n612), .A4(n710), .Y(n559) );
  AND2X1_RVT U757 ( .A1(n560), .A2(n559), .Y(n563) );
  NAND2X0_RVT U758 ( .A1(n561), .A2(n715), .Y(n562) );
  AND2X1_RVT U759 ( .A1(n563), .A2(n562), .Y(n744) );
  AO22X1_RVT U760 ( .A1(n592), .A2(n782), .A3(n564), .A4(n779), .Y(n771) );
  NAND2X0_RVT U761 ( .A1(n774), .A2(n771), .Y(n565) );
  OA22X1_RVT U762 ( .A1(n744), .A2(n758), .A3(n775), .A4(n565), .Y(n566) );
  NAND3X0_RVT U763 ( .A1(n568), .A2(n567), .A3(n566), .Y(div_shl_tmp[96]) );
  NOR2X0_RVT U764 ( .A1(n761), .A2(div_shl_tmp[96]), .Y(
        div_frac_add_in2_in[43]) );
  OA22X1_RVT U765 ( .A1(n631), .A2(n648), .A3(n630), .A4(n646), .Y(n581) );
  AOI22X1_RVT U766 ( .A1(n785), .A2(n570), .A3(n583), .A4(n569), .Y(n580) );
  NAND2X0_RVT U767 ( .A1(n708), .A2(n635), .Y(n573) );
  OA22X1_RVT U768 ( .A1(n571), .A2(n34), .A3(n629), .A4(n710), .Y(n572) );
  AND2X1_RVT U769 ( .A1(n573), .A2(n572), .Y(n576) );
  NAND2X0_RVT U770 ( .A1(n574), .A2(n715), .Y(n575) );
  AND2X1_RVT U771 ( .A1(n576), .A2(n575), .Y(n746) );
  AO22X1_RVT U772 ( .A1(n592), .A2(n783), .A3(n577), .A4(n779), .Y(n772) );
  NAND2X0_RVT U773 ( .A1(n774), .A2(n772), .Y(n578) );
  OA22X1_RVT U774 ( .A1(n746), .A2(n758), .A3(n775), .A4(n578), .Y(n579) );
  NAND3X0_RVT U775 ( .A1(n581), .A2(n580), .A3(n579), .Y(div_shl_tmp[95]) );
  NOR2X0_RVT U776 ( .A1(n761), .A2(div_shl_tmp[95]), .Y(
        div_frac_add_in2_in[42]) );
  OA22X1_RVT U777 ( .A1(n704), .A2(n648), .A3(n649), .A4(n646), .Y(n596) );
  AOI22X1_RVT U778 ( .A1(n785), .A2(n584), .A3(n583), .A4(n582), .Y(n595) );
  NAND2X0_RVT U779 ( .A1(n708), .A2(n709), .Y(n587) );
  OA22X1_RVT U780 ( .A1(n585), .A2(n34), .A3(n647), .A4(n710), .Y(n586) );
  AND2X1_RVT U781 ( .A1(n587), .A2(n586), .Y(n590) );
  NAND2X0_RVT U782 ( .A1(n588), .A2(n715), .Y(n589) );
  AND2X1_RVT U783 ( .A1(n590), .A2(n589), .Y(n748) );
  AO22X1_RVT U784 ( .A1(n592), .A2(n784), .A3(n591), .A4(n779), .Y(n773) );
  NAND2X0_RVT U785 ( .A1(n774), .A2(n773), .Y(n593) );
  OA22X1_RVT U786 ( .A1(n748), .A2(n758), .A3(n775), .A4(n593), .Y(n594) );
  NAND3X0_RVT U787 ( .A1(n596), .A2(n595), .A3(n594), .Y(div_shl_tmp[94]) );
  NOR2X0_RVT U788 ( .A1(n761), .A2(div_shl_tmp[94]), .Y(
        div_frac_add_in2_in[41]) );
  OA22X1_RVT U789 ( .A1(n598), .A2(n705), .A3(n597), .A4(n650), .Y(n611) );
  OA22X1_RVT U790 ( .A1(n600), .A2(n648), .A3(n599), .A4(n646), .Y(n610) );
  OA222X1_RVT U791 ( .A1(n779), .A2(n605), .A3(n604), .A4(n603), .A5(n710), 
        .A6(n602), .Y(n750) );
  AO22X1_RVT U792 ( .A1(div_shl_cnta[3]), .A2(n607), .A3(n779), .A4(n606), .Y(
        n776) );
  NAND2X0_RVT U793 ( .A1(n776), .A2(n774), .Y(n608) );
  OA22X1_RVT U794 ( .A1(n750), .A2(n758), .A3(n775), .A4(n608), .Y(n609) );
  NAND3X0_RVT U795 ( .A1(n611), .A2(n610), .A3(n609), .Y(div_shl_tmp[93]) );
  NOR2X0_RVT U796 ( .A1(n761), .A2(div_shl_tmp[93]), .Y(
        div_frac_add_in2_in[40]) );
  OA22X1_RVT U797 ( .A1(n613), .A2(n648), .A3(n612), .A4(n646), .Y(n628) );
  OA22X1_RVT U798 ( .A1(n615), .A2(n705), .A3(n614), .A4(n650), .Y(n627) );
  AO22X1_RVT U799 ( .A1(n715), .A2(n782), .A3(n21), .A4(n616), .Y(n777) );
  INVX1_RVT U800 ( .A(n777), .Y(n754) );
  NAND2X0_RVT U801 ( .A1(n708), .A2(n617), .Y(n622) );
  OA22X1_RVT U802 ( .A1(n620), .A2(n34), .A3(n619), .A4(n710), .Y(n621) );
  AND2X1_RVT U803 ( .A1(n622), .A2(n621), .Y(n625) );
  NAND2X0_RVT U804 ( .A1(n623), .A2(n715), .Y(n624) );
  AND2X1_RVT U805 ( .A1(n625), .A2(n624), .Y(n753) );
  OA22X1_RVT U806 ( .A1(n754), .A2(n736), .A3(n753), .A4(n758), .Y(n626) );
  NAND3X0_RVT U807 ( .A1(n628), .A2(n627), .A3(n626), .Y(div_shl_tmp[92]) );
  NOR2X0_RVT U808 ( .A1(n761), .A2(div_shl_tmp[92]), .Y(
        div_frac_add_in2_in[39]) );
  OA22X1_RVT U809 ( .A1(n630), .A2(n648), .A3(n629), .A4(n646), .Y(n645) );
  OA22X1_RVT U810 ( .A1(n632), .A2(n705), .A3(n631), .A4(n650), .Y(n644) );
  AO22X1_RVT U811 ( .A1(n715), .A2(n783), .A3(n21), .A4(n633), .Y(n778) );
  INVX1_RVT U812 ( .A(n778), .Y(n756) );
  NAND2X0_RVT U813 ( .A1(n708), .A2(n634), .Y(n639) );
  OA22X1_RVT U814 ( .A1(n637), .A2(n34), .A3(n636), .A4(n710), .Y(n638) );
  AND2X1_RVT U815 ( .A1(n639), .A2(n638), .Y(n642) );
  NAND2X0_RVT U816 ( .A1(n640), .A2(n715), .Y(n641) );
  AND2X1_RVT U817 ( .A1(n642), .A2(n641), .Y(n755) );
  OA22X1_RVT U818 ( .A1(n756), .A2(n736), .A3(n755), .A4(n758), .Y(n643) );
  NAND3X0_RVT U819 ( .A1(n645), .A2(n644), .A3(n643), .Y(div_shl_tmp[91]) );
  NOR2X0_RVT U820 ( .A1(n761), .A2(div_shl_tmp[91]), .Y(
        div_frac_add_in2_in[38]) );
  OA22X1_RVT U821 ( .A1(n649), .A2(n648), .A3(n647), .A4(n646), .Y(n721) );
  OA22X1_RVT U822 ( .A1(n706), .A2(n705), .A3(n704), .A4(n650), .Y(n720) );
  NAND2X0_RVT U823 ( .A1(n708), .A2(n707), .Y(n714) );
  OA22X1_RVT U824 ( .A1(n712), .A2(n34), .A3(n711), .A4(n710), .Y(n713) );
  AND2X1_RVT U825 ( .A1(n714), .A2(n713), .Y(n718) );
  NAND2X0_RVT U826 ( .A1(n716), .A2(n715), .Y(n717) );
  AND2X1_RVT U827 ( .A1(n718), .A2(n717), .Y(n760) );
  NAND2X0_RVT U828 ( .A1(n780), .A2(n779), .Y(n757) );
  OA22X1_RVT U829 ( .A1(n760), .A2(n758), .A3(n736), .A4(n757), .Y(n719) );
  NAND3X0_RVT U830 ( .A1(n721), .A2(n720), .A3(n719), .Y(div_shl_tmp[90]) );
  NOR2X0_RVT U831 ( .A1(n761), .A2(div_shl_tmp[90]), .Y(
        div_frac_add_in2_in[37]) );
  AO222X1_RVT U832 ( .A1(n724), .A2(n25), .A3(n723), .A4(n752), .A5(n722), 
        .A6(n781), .Y(div_shl_tmp[89]) );
  NOR2X0_RVT U833 ( .A1(n761), .A2(div_shl_tmp[89]), .Y(
        div_frac_add_in2_in[36]) );
  AND2X1_RVT U834 ( .A1(div_shl_cnta[5]), .A2(n725), .Y(n732) );
  AO222X1_RVT U835 ( .A1(n782), .A2(n732), .A3(n727), .A4(n752), .A5(n726), 
        .A6(n25), .Y(div_shl_tmp[88]) );
  NOR2X0_RVT U836 ( .A1(n761), .A2(div_shl_tmp[88]), .Y(
        div_frac_add_in2_in[35]) );
  AO222X1_RVT U837 ( .A1(n783), .A2(n732), .A3(n729), .A4(n752), .A5(n728), 
        .A6(n25), .Y(div_shl_tmp[87]) );
  NOR2X0_RVT U838 ( .A1(n761), .A2(div_shl_tmp[87]), .Y(
        div_frac_add_in2_in[34]) );
  AO222X1_RVT U839 ( .A1(n784), .A2(n732), .A3(n731), .A4(n752), .A5(n730), 
        .A6(n25), .Y(div_shl_tmp[86]) );
  NOR2X0_RVT U840 ( .A1(n761), .A2(div_shl_tmp[86]), .Y(
        div_frac_add_in2_in[33]) );
  OAI222X1_RVT U841 ( .A1(n736), .A2(n735), .A3(n759), .A4(n734), .A5(n758), 
        .A6(n733), .Y(div_shl_tmp[85]) );
  NOR2X0_RVT U842 ( .A1(n761), .A2(div_shl_tmp[85]), .Y(
        div_frac_add_in2_in[32]) );
  OAI22X1_RVT U843 ( .A1(n738), .A2(n758), .A3(n737), .A4(n759), .Y(
        div_shl_tmp[84]) );
  NOR2X0_RVT U844 ( .A1(n761), .A2(div_shl_tmp[84]), .Y(
        div_frac_add_in2_in[31]) );
  OAI22X1_RVT U845 ( .A1(n740), .A2(n758), .A3(n739), .A4(n759), .Y(
        div_shl_tmp[83]) );
  NOR2X0_RVT U846 ( .A1(n761), .A2(div_shl_tmp[83]), .Y(
        div_frac_add_in2_in[30]) );
  AO22X1_RVT U847 ( .A1(d4stg_fdiv), .A2(n741), .A3(d6stg_fdiv), .A4(
        d6stg_fdivs), .Y(div_frac_add_in2_in[29]) );
  INVX1_RVT U848 ( .A(n742), .Y(n743) );
  AO22X1_RVT U849 ( .A1(n752), .A2(n770), .A3(n25), .A4(n743), .Y(
        div_shl_tmp[81]) );
  NOR2X0_RVT U850 ( .A1(n761), .A2(div_shl_tmp[81]), .Y(
        div_frac_add_in2_in[28]) );
  INVX1_RVT U851 ( .A(n744), .Y(n745) );
  AO22X1_RVT U852 ( .A1(n752), .A2(n771), .A3(n25), .A4(n745), .Y(
        div_shl_tmp[80]) );
  NOR2X0_RVT U853 ( .A1(n761), .A2(div_shl_tmp[80]), .Y(
        div_frac_add_in2_in[27]) );
  INVX1_RVT U854 ( .A(n746), .Y(n747) );
  AO22X1_RVT U855 ( .A1(n752), .A2(n772), .A3(n25), .A4(n747), .Y(
        div_shl_tmp[79]) );
  NOR2X0_RVT U856 ( .A1(n761), .A2(div_shl_tmp[79]), .Y(
        div_frac_add_in2_in[26]) );
  INVX1_RVT U857 ( .A(n748), .Y(n749) );
  AO22X1_RVT U858 ( .A1(n752), .A2(n773), .A3(n25), .A4(n749), .Y(
        div_shl_tmp[78]) );
  NOR2X0_RVT U859 ( .A1(n761), .A2(div_shl_tmp[78]), .Y(
        div_frac_add_in2_in[25]) );
  INVX1_RVT U860 ( .A(n750), .Y(n751) );
  AO22X1_RVT U861 ( .A1(n752), .A2(n776), .A3(n25), .A4(n751), .Y(
        div_shl_tmp[77]) );
  NOR2X0_RVT U862 ( .A1(n761), .A2(div_shl_tmp[77]), .Y(
        div_frac_add_in2_in[24]) );
  OAI22X1_RVT U863 ( .A1(n754), .A2(n758), .A3(n753), .A4(n759), .Y(
        div_shl_tmp[76]) );
  NOR2X0_RVT U864 ( .A1(n761), .A2(div_shl_tmp[76]), .Y(
        div_frac_add_in2_in[23]) );
  OAI22X1_RVT U865 ( .A1(n756), .A2(n758), .A3(n755), .A4(n759), .Y(
        div_shl_tmp[75]) );
  NOR2X0_RVT U866 ( .A1(n761), .A2(div_shl_tmp[75]), .Y(
        div_frac_add_in2_in[22]) );
  OAI22X1_RVT U867 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .Y(
        div_shl_tmp[74]) );
  NOR2X0_RVT U868 ( .A1(n761), .A2(div_shl_tmp[74]), .Y(
        div_frac_add_in2_in[21]) );
  AND2X1_RVT U869 ( .A1(n762), .A2(n775), .Y(div_shl_tmp[73]) );
  NOR2X0_RVT U870 ( .A1(div_shl_tmp[73]), .A2(n761), .Y(
        div_frac_add_in2_in[20]) );
  AND2X1_RVT U871 ( .A1(n775), .A2(n763), .Y(div_shl_tmp[72]) );
  NOR2X0_RVT U872 ( .A1(div_shl_tmp[72]), .A2(n761), .Y(
        div_frac_add_in2_in[19]) );
  AND2X1_RVT U873 ( .A1(n775), .A2(n764), .Y(div_shl_tmp[71]) );
  NOR2X0_RVT U874 ( .A1(div_shl_tmp[71]), .A2(n761), .Y(
        div_frac_add_in2_in[18]) );
  AND2X1_RVT U875 ( .A1(n775), .A2(n765), .Y(div_shl_tmp[70]) );
  NOR2X0_RVT U876 ( .A1(div_shl_tmp[70]), .A2(n761), .Y(
        div_frac_add_in2_in[17]) );
  NOR2X0_RVT U877 ( .A1(div_shl_cnta[5]), .A2(n766), .Y(div_shl_tmp[69]) );
  NOR2X0_RVT U878 ( .A1(div_shl_tmp[69]), .A2(n761), .Y(
        div_frac_add_in2_in[16]) );
  AND2X1_RVT U879 ( .A1(n25), .A2(n767), .Y(div_shl_tmp[68]) );
  NOR2X0_RVT U880 ( .A1(div_shl_tmp[68]), .A2(n761), .Y(
        div_frac_add_in2_in[15]) );
  AND2X1_RVT U881 ( .A1(n25), .A2(n768), .Y(div_shl_tmp[67]) );
  NOR2X0_RVT U882 ( .A1(div_shl_tmp[67]), .A2(n761), .Y(
        div_frac_add_in2_in[14]) );
  AND2X1_RVT U883 ( .A1(n25), .A2(n769), .Y(div_shl_tmp[66]) );
  NOR2X0_RVT U884 ( .A1(div_shl_tmp[66]), .A2(n761), .Y(
        div_frac_add_in2_in[13]) );
  AND3X1_RVT U885 ( .A1(n770), .A2(n775), .A3(n774), .Y(div_shl_tmp[65]) );
  NOR2X0_RVT U886 ( .A1(div_shl_tmp[65]), .A2(n761), .Y(
        div_frac_add_in2_in[12]) );
  AND3X1_RVT U887 ( .A1(n775), .A2(n774), .A3(n771), .Y(div_shl_tmp[64]) );
  NOR2X0_RVT U888 ( .A1(div_shl_tmp[64]), .A2(n761), .Y(
        div_frac_add_in2_in[11]) );
  AND3X1_RVT U889 ( .A1(n775), .A2(n774), .A3(n772), .Y(div_shl_tmp[63]) );
  NOR2X0_RVT U890 ( .A1(div_shl_tmp[63]), .A2(n761), .Y(
        div_frac_add_in2_in[10]) );
  AND3X1_RVT U891 ( .A1(n775), .A2(n774), .A3(n773), .Y(div_shl_tmp[62]) );
  NOR2X0_RVT U892 ( .A1(div_shl_tmp[62]), .A2(n761), .Y(div_frac_add_in2_in[9]) );
  AND3X1_RVT U893 ( .A1(n776), .A2(n775), .A3(n774), .Y(div_shl_tmp[61]) );
  NOR2X0_RVT U894 ( .A1(div_shl_tmp[61]), .A2(n761), .Y(div_frac_add_in2_in[8]) );
  AND2X1_RVT U895 ( .A1(n25), .A2(n777), .Y(div_shl_tmp[60]) );
  NOR2X0_RVT U896 ( .A1(div_shl_tmp[60]), .A2(n761), .Y(div_frac_add_in2_in[7]) );
  AND2X1_RVT U897 ( .A1(n25), .A2(n778), .Y(div_shl_tmp[59]) );
  NOR2X0_RVT U898 ( .A1(div_shl_tmp[59]), .A2(n761), .Y(div_frac_add_in2_in[6]) );
  AND3X1_RVT U899 ( .A1(n25), .A2(n780), .A3(n779), .Y(div_shl_tmp[58]) );
  NOR2X0_RVT U900 ( .A1(div_shl_tmp[58]), .A2(n761), .Y(div_frac_add_in2_in[5]) );
  AND2X1_RVT U901 ( .A1(n781), .A2(n25), .Y(div_shl_tmp[57]) );
  NOR2X0_RVT U902 ( .A1(div_shl_tmp[57]), .A2(n761), .Y(div_frac_add_in2_in[4]) );
  AND2X1_RVT U903 ( .A1(n785), .A2(n782), .Y(div_shl_tmp[56]) );
  NOR2X0_RVT U904 ( .A1(div_shl_tmp[56]), .A2(n761), .Y(div_frac_add_in2_in[3]) );
  AND2X1_RVT U905 ( .A1(n785), .A2(n783), .Y(div_shl_tmp[55]) );
  NOR2X0_RVT U906 ( .A1(div_shl_tmp[55]), .A2(n761), .Y(div_frac_add_in2_in[2]) );
  AND2X1_RVT U907 ( .A1(n785), .A2(n784), .Y(div_shl_tmp[54]) );
  NOR2X0_RVT U908 ( .A1(div_shl_tmp[54]), .A2(n761), .Y(div_frac_add_in2_in[1]) );
  AO22X1_RVT U909 ( .A1(d4stg_fdiv), .A2(n786), .A3(d6stg_fdiv), .A4(
        d6stg_fdivd), .Y(div_frac_add_in2_in[0]) );
  AO22X1_RVT U910 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[1]), .A3(n799), 
        .A4(div_frac_outa[0]), .Y(d6stg_frac_1) );
  AND2X1_RVT U911 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[0]), .Y(
        d6stg_frac_0) );
  AO222X1_RVT U912 ( .A1(d4stg_fdiv), .A2(div_shl_save[52]), .A3(n795), .A4(
        n787), .A5(n796), .A6(div_frac_add_in1[51]), .Y(
        div_frac_add_in1_in[52]) );
  AO22X1_RVT U913 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[31]), .A3(n799), .A4(div_frac_outa[30]), .Y(d6stg_frac_31) );
  AO22X1_RVT U914 ( .A1(d4stg_fdiv), .A2(div_shl_save[29]), .A3(d6stg_fdiv), 
        .A4(d6stg_frac_31), .Y(n790) );
  AO22X1_RVT U915 ( .A1(div_frac_add_in1[28]), .A2(n796), .A3(n795), .A4(n788), 
        .Y(n789) );
  OR2X1_RVT U916 ( .A1(n790), .A2(n789), .Y(div_frac_add_in1_in[29]) );
  AO22X1_RVT U917 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[30]), .A3(n799), .A4(div_frac_outa[29]), .Y(d6stg_frac_30) );
  AO22X1_RVT U918 ( .A1(d4stg_fdiv), .A2(div_shl_save[28]), .A3(n795), .A4(
        n791), .Y(n793) );
  AND2X1_RVT U919 ( .A1(d6stg_fdiv), .A2(d6stg_fdivd), .Y(n800) );
  AO22X1_RVT U920 ( .A1(n800), .A2(d6stg_frac_30), .A3(div_frac_add_in1[27]), 
        .A4(n796), .Y(n792) );
  OR2X1_RVT U921 ( .A1(n793), .A2(n792), .Y(div_frac_add_in1_in[28]) );
  AO22X1_RVT U922 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[29]), .A3(n799), .A4(div_frac_outa[28]), .Y(d6stg_frac_29) );
  AO22X1_RVT U923 ( .A1(d4stg_fdiv), .A2(div_shl_save[27]), .A3(n795), .A4(
        n794), .Y(n798) );
  AO22X1_RVT U924 ( .A1(n800), .A2(d6stg_frac_29), .A3(div_frac_add_in1[26]), 
        .A4(n796), .Y(n797) );
  OR2X1_RVT U925 ( .A1(n798), .A2(n797), .Y(div_frac_add_in1_in[27]) );
  AO22X1_RVT U926 ( .A1(d6stg_frac_out_nosh), .A2(div_frac_outa[2]), .A3(n799), 
        .A4(div_frac_outa[1]), .Y(d6stg_frac_2) );
  AO22X1_RVT U927 ( .A1(d4stg_fdiv), .A2(div_shl_save[0]), .A3(n800), .A4(
        d6stg_frac_2), .Y(div_frac_add_in1_in[0]) );
  NOR4X1_RVT U928 ( .A1(div_frac_add_in1[49]), .A2(div_frac_add_in1[50]), .A3(
        div_frac_add_in1[52]), .A4(div_frac_add_in1[54]), .Y(n817) );
  NOR4X1_RVT U929 ( .A1(div_frac_add_in1[48]), .A2(div_frac_add_in1[46]), .A3(
        div_frac_add_in1[47]), .A4(div_frac_add_in1[51]), .Y(n816) );
  NOR4X1_RVT U930 ( .A1(div_frac_add_in1[13]), .A2(div_frac_add_in1[14]), .A3(
        div_frac_add_in1[15]), .A4(div_frac_add_in1[16]), .Y(n804) );
  NOR4X1_RVT U931 ( .A1(div_frac_add_in1[19]), .A2(div_frac_add_in1[17]), .A3(
        div_frac_add_in1[18]), .A4(div_frac_add_in1[20]), .Y(n803) );
  NOR4X1_RVT U932 ( .A1(div_frac_add_in1[21]), .A2(div_frac_add_in1[22]), .A3(
        div_frac_add_in1[23]), .A4(div_frac_add_in1[26]), .Y(n802) );
  NOR4X1_RVT U933 ( .A1(div_frac_add_in1[24]), .A2(div_frac_add_in1[25]), .A3(
        div_frac_add_in1[27]), .A4(div_frac_add_in1[28]), .Y(n801) );
  AND4X1_RVT U934 ( .A1(n804), .A2(n803), .A3(n802), .A4(n801), .Y(n815) );
  NOR4X1_RVT U935 ( .A1(div_frac_add_in1[1]), .A2(div_frac_add_in1[2]), .A3(
        div_frac_add_in1[5]), .A4(div_frac_add_in1[3]), .Y(n813) );
  NOR4X1_RVT U936 ( .A1(div_frac_add_in1[4]), .A2(div_frac_add_in1[6]), .A3(
        div_frac_add_in1[7]), .A4(div_frac_add_in1[8]), .Y(n812) );
  OR4X1_RVT U937 ( .A1(div_frac_add_in1[9]), .A2(div_frac_add_in1[12]), .A3(
        div_frac_add_in1[10]), .A4(div_frac_add_in1[11]), .Y(n805) );
  NOR4X1_RVT U938 ( .A1(div_frac_add_in1[29]), .A2(div_frac_add_in1[0]), .A3(
        div_frac_add_in1[53]), .A4(n805), .Y(n811) );
  NOR4X1_RVT U939 ( .A1(div_frac_add_in1[30]), .A2(div_frac_add_in1[31]), .A3(
        div_frac_add_in1[34]), .A4(div_frac_add_in1[32]), .Y(n809) );
  NOR4X1_RVT U940 ( .A1(div_frac_add_in1[33]), .A2(div_frac_add_in1[35]), .A3(
        div_frac_add_in1[36]), .A4(div_frac_add_in1[37]), .Y(n808) );
  NOR4X1_RVT U941 ( .A1(div_frac_add_in1[38]), .A2(div_frac_add_in1[41]), .A3(
        div_frac_add_in1[39]), .A4(div_frac_add_in1[40]), .Y(n807) );
  NOR4X1_RVT U942 ( .A1(div_frac_add_in1[42]), .A2(div_frac_add_in1[43]), .A3(
        div_frac_add_in1[44]), .A4(div_frac_add_in1[45]), .Y(n806) );
  AND4X1_RVT U943 ( .A1(n809), .A2(n808), .A3(n807), .A4(n806), .Y(n810) );
  AND4X1_RVT U944 ( .A1(n813), .A2(n812), .A3(n811), .A4(n810), .Y(n814) );
  NAND4X0_RVT U945 ( .A1(n817), .A2(n816), .A3(n815), .A4(n814), .Y(
        div_frac_add_in1_neq_0) );
  AO22X1_RVT U946 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[54]), 
        .A3(div_norm_frac_in1_sng_dnrm), .A4(div_frac_in1[54]), .Y(n821) );
  AO22X1_RVT U947 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[51]), 
        .A3(div_frac_in1[51]), .A4(div_norm_frac_in1_dbl_dnrm), .Y(n819) );
  OR4X1_RVT U948 ( .A1(div_norm_frac_in2_dbl_norm), .A2(
        div_norm_frac_in1_dbl_norm), .A3(div_norm_qnan), .A4(
        div_norm_frac_in1_sng_norm), .Y(n818) );
  OR2X1_RVT U949 ( .A1(n819), .A2(n818), .Y(n820) );
  NOR4X1_RVT U950 ( .A1(div_norm_frac_in2_sng_norm), .A2(div_norm_inf), .A3(
        n821), .A4(n820), .Y(n703) );
  AO22X1_RVT U951 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[53]), 
        .A3(div_norm_frac_in2_dbl_dnrm), .A4(div_frac_in2[50]), .Y(n828) );
  OR2X1_RVT U952 ( .A1(div_frac_in2[51]), .A2(d1stg_snan_dbl_in2), .Y(n822) );
  AO22X1_RVT U953 ( .A1(div_norm_frac_in2_dbl_norm), .A2(n822), .A3(
        div_norm_frac_in1_sng_dnrm), .A4(div_frac_in1[53]), .Y(n827) );
  OA21X1_RVT U954 ( .A1(div_frac_in1[51]), .A2(d1stg_snan_dbl_in1), .A3(
        div_norm_frac_in1_dbl_norm), .Y(n823) );
  AO221X1_RVT U955 ( .A1(div_norm_frac_in2_sng_norm), .A2(d1stg_snan_sng_in2), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[54]), .A5(n823), .Y(
        n826) );
  AO221X1_RVT U956 ( .A1(div_norm_frac_in1_sng_norm), .A2(d1stg_snan_sng_in1), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[54]), .A5(
        div_norm_qnan), .Y(n824) );
  AO21X1_RVT U957 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[50]), 
        .A3(n824), .Y(n825) );
  NOR4X1_RVT U958 ( .A1(n828), .A2(n827), .A3(n826), .A4(n825), .Y(n702) );
  AO22X1_RVT U959 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[52]), 
        .A3(div_frac_in2[53]), .A4(div_norm_frac_in2_sng_norm), .Y(n833) );
  AO22X1_RVT U960 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[49]), 
        .A3(div_frac_in1[53]), .A4(div_norm_frac_in1_sng_norm), .Y(n832) );
  AO22X1_RVT U961 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[52]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[49]), .Y(n830) );
  AO22X1_RVT U962 ( .A1(div_frac_in2[50]), .A2(div_norm_frac_in2_dbl_norm), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[50]), .Y(n829) );
  OR2X1_RVT U963 ( .A1(n830), .A2(n829), .Y(n831) );
  NOR4X1_RVT U964 ( .A1(div_norm_qnan), .A2(n833), .A3(n832), .A4(n831), .Y(
        n701) );
  AO22X1_RVT U965 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[51]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[52]), .Y(n838) );
  AO22X1_RVT U966 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[48]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[52]), .Y(n837) );
  AO22X1_RVT U967 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[51]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[48]), .Y(n835) );
  AO22X1_RVT U968 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[49]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[49]), .Y(n834) );
  OR2X1_RVT U969 ( .A1(n835), .A2(n834), .Y(n836) );
  NOR4X1_RVT U970 ( .A1(div_norm_qnan), .A2(n838), .A3(n837), .A4(n836), .Y(
        n700) );
  AO22X1_RVT U971 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[50]), 
        .A3(div_frac_in2[51]), .A4(div_norm_frac_in2_sng_norm), .Y(n843) );
  AO22X1_RVT U972 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[47]), 
        .A3(div_frac_in1[51]), .A4(div_norm_frac_in1_sng_norm), .Y(n842) );
  AO22X1_RVT U973 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[50]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[47]), .Y(n840) );
  AO22X1_RVT U974 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[48]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[48]), .Y(n839) );
  OR2X1_RVT U975 ( .A1(n840), .A2(n839), .Y(n841) );
  NOR4X1_RVT U976 ( .A1(div_norm_qnan), .A2(n843), .A3(n842), .A4(n841), .Y(
        n699) );
  AO22X1_RVT U977 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[49]), 
        .A3(div_frac_in2[50]), .A4(div_norm_frac_in2_sng_norm), .Y(n848) );
  AO22X1_RVT U978 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[46]), 
        .A3(div_frac_in1[50]), .A4(div_norm_frac_in1_sng_norm), .Y(n847) );
  AO22X1_RVT U979 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[49]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[46]), .Y(n845) );
  AO22X1_RVT U980 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[47]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[47]), .Y(n844) );
  OR2X1_RVT U981 ( .A1(n845), .A2(n844), .Y(n846) );
  NOR4X1_RVT U982 ( .A1(div_norm_qnan), .A2(n848), .A3(n847), .A4(n846), .Y(
        n698) );
  AO22X1_RVT U983 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[48]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[49]), .Y(n853) );
  AO22X1_RVT U984 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[45]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[49]), .Y(n852) );
  AO22X1_RVT U985 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[48]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[45]), .Y(n850) );
  AO22X1_RVT U986 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[46]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[46]), .Y(n849) );
  OR2X1_RVT U987 ( .A1(n850), .A2(n849), .Y(n851) );
  NOR4X1_RVT U988 ( .A1(div_norm_qnan), .A2(n853), .A3(n852), .A4(n851), .Y(
        n697) );
  AO22X1_RVT U989 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[47]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[48]), .Y(n858) );
  AO22X1_RVT U990 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[44]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[48]), .Y(n857) );
  AO22X1_RVT U991 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[47]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[44]), .Y(n855) );
  AO22X1_RVT U992 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[45]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[45]), .Y(n854) );
  OR2X1_RVT U993 ( .A1(n855), .A2(n854), .Y(n856) );
  NOR4X1_RVT U994 ( .A1(div_norm_qnan), .A2(n858), .A3(n857), .A4(n856), .Y(
        n696) );
  AO22X1_RVT U995 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[46]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[47]), .Y(n863) );
  AO22X1_RVT U996 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[43]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[47]), .Y(n862) );
  AO22X1_RVT U997 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[46]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[43]), .Y(n860) );
  AO22X1_RVT U998 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[44]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[44]), .Y(n859) );
  OR2X1_RVT U999 ( .A1(n860), .A2(n859), .Y(n861) );
  NOR4X1_RVT U1000 ( .A1(div_norm_qnan), .A2(n863), .A3(n862), .A4(n861), .Y(
        n695) );
  AO22X1_RVT U1001 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[45]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[46]), .Y(n868) );
  AO22X1_RVT U1002 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[42]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[46]), .Y(n867) );
  AO22X1_RVT U1003 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[45]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[42]), .Y(n865) );
  AO22X1_RVT U1004 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[43]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[43]), .Y(n864) );
  OR2X1_RVT U1005 ( .A1(n865), .A2(n864), .Y(n866) );
  NOR4X1_RVT U1006 ( .A1(div_norm_qnan), .A2(n868), .A3(n867), .A4(n866), .Y(
        n694) );
  AO22X1_RVT U1007 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[44]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[45]), .Y(n873) );
  AO22X1_RVT U1008 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[41]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[45]), .Y(n872) );
  AO22X1_RVT U1009 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[44]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[41]), .Y(n870) );
  AO22X1_RVT U1010 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[42]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[42]), .Y(n869) );
  OR2X1_RVT U1011 ( .A1(n870), .A2(n869), .Y(n871) );
  NOR4X1_RVT U1012 ( .A1(div_norm_qnan), .A2(n873), .A3(n872), .A4(n871), .Y(
        n693) );
  AO22X1_RVT U1013 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[43]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[44]), .Y(n878) );
  AO22X1_RVT U1014 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[40]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[44]), .Y(n877) );
  AO22X1_RVT U1015 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[43]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[40]), .Y(n875) );
  AO22X1_RVT U1016 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[41]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[41]), .Y(n874) );
  OR2X1_RVT U1017 ( .A1(n875), .A2(n874), .Y(n876) );
  NOR4X1_RVT U1018 ( .A1(div_norm_qnan), .A2(n878), .A3(n877), .A4(n876), .Y(
        n692) );
  AO22X1_RVT U1019 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[42]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[43]), .Y(n883) );
  AO22X1_RVT U1020 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[39]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[43]), .Y(n882) );
  AO22X1_RVT U1021 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[42]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[39]), .Y(n880) );
  AO22X1_RVT U1022 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[40]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[40]), .Y(n879) );
  OR2X1_RVT U1023 ( .A1(n880), .A2(n879), .Y(n881) );
  NOR4X1_RVT U1024 ( .A1(div_norm_qnan), .A2(n883), .A3(n882), .A4(n881), .Y(
        n691) );
  AO22X1_RVT U1025 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[41]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[42]), .Y(n888) );
  AO22X1_RVT U1026 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[38]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[42]), .Y(n887) );
  AO22X1_RVT U1027 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[41]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[38]), .Y(n885) );
  AO22X1_RVT U1028 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[39]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[39]), .Y(n884) );
  OR2X1_RVT U1029 ( .A1(n885), .A2(n884), .Y(n886) );
  NOR4X1_RVT U1030 ( .A1(div_norm_qnan), .A2(n888), .A3(n887), .A4(n886), .Y(
        n690) );
  AO22X1_RVT U1031 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[40]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[41]), .Y(n893) );
  AO22X1_RVT U1032 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[37]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[41]), .Y(n892) );
  AO22X1_RVT U1033 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[40]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[37]), .Y(n890) );
  AO22X1_RVT U1034 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[38]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[38]), .Y(n889) );
  OR2X1_RVT U1035 ( .A1(n890), .A2(n889), .Y(n891) );
  NOR4X1_RVT U1036 ( .A1(div_norm_qnan), .A2(n893), .A3(n892), .A4(n891), .Y(
        n689) );
  AO22X1_RVT U1037 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[39]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[40]), .Y(n898) );
  AO22X1_RVT U1038 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[36]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[40]), .Y(n897) );
  AO22X1_RVT U1039 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[39]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[36]), .Y(n895) );
  AO22X1_RVT U1040 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[37]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[37]), .Y(n894) );
  OR2X1_RVT U1041 ( .A1(n895), .A2(n894), .Y(n896) );
  NOR4X1_RVT U1042 ( .A1(div_norm_qnan), .A2(n898), .A3(n897), .A4(n896), .Y(
        n688) );
  AO22X1_RVT U1043 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[38]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[39]), .Y(n903) );
  AO22X1_RVT U1044 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[35]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[39]), .Y(n902) );
  AO22X1_RVT U1045 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[38]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[35]), .Y(n900) );
  AO22X1_RVT U1046 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[36]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[36]), .Y(n899) );
  OR2X1_RVT U1047 ( .A1(n900), .A2(n899), .Y(n901) );
  NOR4X1_RVT U1048 ( .A1(div_norm_qnan), .A2(n903), .A3(n902), .A4(n901), .Y(
        n687) );
  AO22X1_RVT U1049 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[37]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[38]), .Y(n908) );
  AO22X1_RVT U1050 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[34]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[38]), .Y(n907) );
  AO22X1_RVT U1051 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[37]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[34]), .Y(n905) );
  AO22X1_RVT U1052 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[35]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[35]), .Y(n904) );
  OR2X1_RVT U1053 ( .A1(n905), .A2(n904), .Y(n906) );
  NOR4X1_RVT U1054 ( .A1(div_norm_qnan), .A2(n908), .A3(n907), .A4(n906), .Y(
        n686) );
  AO22X1_RVT U1055 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[36]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[37]), .Y(n913) );
  AO22X1_RVT U1056 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[33]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[37]), .Y(n912) );
  AO22X1_RVT U1057 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[36]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[33]), .Y(n910) );
  AO22X1_RVT U1058 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[34]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[34]), .Y(n909) );
  OR2X1_RVT U1059 ( .A1(n910), .A2(n909), .Y(n911) );
  NOR4X1_RVT U1060 ( .A1(div_norm_qnan), .A2(n913), .A3(n912), .A4(n911), .Y(
        n685) );
  AO22X1_RVT U1061 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[35]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[36]), .Y(n918) );
  AO22X1_RVT U1062 ( .A1(div_norm_frac_in1_dbl_norm), .A2(div_frac_in1[33]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[36]), .Y(n917) );
  AO22X1_RVT U1063 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[35]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[32]), .Y(n915) );
  AO22X1_RVT U1064 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[32]), 
        .A3(div_norm_frac_in2_dbl_norm), .A4(div_frac_in2[33]), .Y(n914) );
  OR2X1_RVT U1065 ( .A1(n915), .A2(n914), .Y(n916) );
  NOR4X1_RVT U1066 ( .A1(div_norm_qnan), .A2(n918), .A3(n917), .A4(n916), .Y(
        n684) );
  AO22X1_RVT U1067 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[34]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[35]), .Y(n923) );
  AO22X1_RVT U1068 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[31]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[35]), .Y(n922) );
  AO22X1_RVT U1069 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[34]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[31]), .Y(n920) );
  AO22X1_RVT U1070 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[32]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[32]), .Y(n919) );
  OR2X1_RVT U1071 ( .A1(n920), .A2(n919), .Y(n921) );
  NOR4X1_RVT U1072 ( .A1(div_norm_qnan), .A2(n923), .A3(n922), .A4(n921), .Y(
        n683) );
  AO22X1_RVT U1073 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[33]), 
        .A3(div_norm_frac_in2_sng_norm), .A4(div_frac_in2[34]), .Y(n928) );
  AO22X1_RVT U1074 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[30]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[34]), .Y(n927) );
  AO22X1_RVT U1075 ( .A1(div_norm_frac_in1_sng_dnrm), .A2(div_frac_in1[33]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[30]), .Y(n925) );
  AO22X1_RVT U1076 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[31]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[31]), .Y(n924) );
  OR2X1_RVT U1077 ( .A1(n925), .A2(n924), .Y(n926) );
  NOR4X1_RVT U1078 ( .A1(div_norm_qnan), .A2(n928), .A3(n927), .A4(n926), .Y(
        n682) );
  AO22X1_RVT U1079 ( .A1(div_norm_frac_in2_sng_dnrm), .A2(div_frac_in2[32]), 
        .A3(div_norm_frac_in1_sng_dnrm), .A4(div_frac_in1[32]), .Y(n933) );
  AO22X1_RVT U1080 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[29]), 
        .A3(div_norm_frac_in1_sng_norm), .A4(div_frac_in1[33]), .Y(n932) );
  AO22X1_RVT U1081 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[29]), 
        .A3(div_norm_frac_in2_dbl_norm), .A4(div_frac_in2[30]), .Y(n930) );
  AO22X1_RVT U1082 ( .A1(div_norm_frac_in2_sng_norm), .A2(div_frac_in2[33]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[30]), .Y(n929) );
  OR2X1_RVT U1083 ( .A1(n930), .A2(n929), .Y(n931) );
  NOR4X1_RVT U1084 ( .A1(div_norm_qnan), .A2(n933), .A3(n932), .A4(n931), .Y(
        n681) );
  AOI22X1_RVT U1085 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[28]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[28]), .Y(n935) );
  AND2X1_RVT U1086 ( .A1(div_norm_qnan), .A2(d1stg_dblop), .Y(n1020) );
  NAND2X0_RVT U1087 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[27]), 
        .Y(n934) );
  NAND3X0_RVT U1088 ( .A1(n935), .A2(n950), .A3(n934), .Y(n936) );
  AOI21X1_RVT U1089 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[27]), 
        .A3(n936), .Y(n679) );
  AOI22X1_RVT U1090 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[27]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[27]), .Y(n938) );
  NAND2X0_RVT U1091 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[26]), 
        .Y(n937) );
  NAND3X0_RVT U1092 ( .A1(n938), .A2(n950), .A3(n937), .Y(n939) );
  AOI21X1_RVT U1093 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[26]), 
        .A3(n939), .Y(n678) );
  AOI22X1_RVT U1094 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[26]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[26]), .Y(n941) );
  NAND2X0_RVT U1095 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[25]), 
        .Y(n940) );
  NAND3X0_RVT U1096 ( .A1(n941), .A2(n950), .A3(n940), .Y(n942) );
  AOI21X1_RVT U1097 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[25]), 
        .A3(n942), .Y(n677) );
  AOI22X1_RVT U1098 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[25]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[25]), .Y(n944) );
  NAND2X0_RVT U1099 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[24]), 
        .Y(n943) );
  NAND3X0_RVT U1100 ( .A1(n944), .A2(n950), .A3(n943), .Y(n945) );
  AOI21X1_RVT U1101 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[24]), 
        .A3(n945), .Y(n676) );
  AOI22X1_RVT U1102 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[24]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[24]), .Y(n947) );
  NAND2X0_RVT U1103 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[23]), 
        .Y(n946) );
  NAND3X0_RVT U1104 ( .A1(n947), .A2(n950), .A3(n946), .Y(n948) );
  AOI21X1_RVT U1105 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[23]), 
        .A3(n948), .Y(n675) );
  AOI22X1_RVT U1106 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[23]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[23]), .Y(n951) );
  INVX1_RVT U1107 ( .A(n1020), .Y(n950) );
  NAND2X0_RVT U1108 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[22]), 
        .Y(n949) );
  NAND3X0_RVT U1109 ( .A1(n951), .A2(n950), .A3(n949), .Y(n952) );
  AOI21X1_RVT U1110 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[22]), 
        .A3(n952), .Y(n674) );
  AOI22X1_RVT U1111 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[22]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[22]), .Y(n954) );
  NAND2X0_RVT U1112 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[21]), 
        .Y(n953) );
  NAND3X0_RVT U1113 ( .A1(n954), .A2(n950), .A3(n953), .Y(n955) );
  AOI21X1_RVT U1114 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[21]), 
        .A3(n955), .Y(n673) );
  AOI22X1_RVT U1115 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[21]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[21]), .Y(n957) );
  NAND2X0_RVT U1116 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[20]), 
        .Y(n956) );
  NAND3X0_RVT U1117 ( .A1(n957), .A2(n950), .A3(n956), .Y(n958) );
  AOI21X1_RVT U1118 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[20]), 
        .A3(n958), .Y(n672) );
  AOI22X1_RVT U1119 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[20]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[20]), .Y(n960) );
  NAND2X0_RVT U1120 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[19]), 
        .Y(n959) );
  NAND3X0_RVT U1121 ( .A1(n960), .A2(n950), .A3(n959), .Y(n961) );
  AOI21X1_RVT U1122 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[19]), 
        .A3(n961), .Y(n671) );
  AOI22X1_RVT U1123 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[19]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[19]), .Y(n963) );
  NAND2X0_RVT U1124 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[18]), 
        .Y(n962) );
  NAND3X0_RVT U1125 ( .A1(n963), .A2(n950), .A3(n962), .Y(n964) );
  AOI21X1_RVT U1126 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[18]), 
        .A3(n964), .Y(n670) );
  AOI22X1_RVT U1127 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[18]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[18]), .Y(n966) );
  NAND2X0_RVT U1128 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[17]), 
        .Y(n965) );
  NAND3X0_RVT U1129 ( .A1(n966), .A2(n950), .A3(n965), .Y(n967) );
  AOI21X1_RVT U1130 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[17]), 
        .A3(n967), .Y(n669) );
  AOI22X1_RVT U1131 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[17]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[17]), .Y(n969) );
  NAND2X0_RVT U1132 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[16]), 
        .Y(n968) );
  NAND3X0_RVT U1133 ( .A1(n969), .A2(n950), .A3(n968), .Y(n970) );
  AOI21X1_RVT U1134 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[16]), 
        .A3(n970), .Y(n668) );
  AOI22X1_RVT U1135 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[16]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[16]), .Y(n972) );
  NAND2X0_RVT U1136 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[15]), 
        .Y(n971) );
  NAND3X0_RVT U1137 ( .A1(n972), .A2(n950), .A3(n971), .Y(n973) );
  AOI21X1_RVT U1138 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[15]), 
        .A3(n973), .Y(n667) );
  AOI22X1_RVT U1139 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[15]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[15]), .Y(n975) );
  NAND2X0_RVT U1140 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[14]), 
        .Y(n974) );
  NAND3X0_RVT U1141 ( .A1(n975), .A2(n950), .A3(n974), .Y(n976) );
  AOI21X1_RVT U1142 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[14]), 
        .A3(n976), .Y(n666) );
  AOI22X1_RVT U1143 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[14]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[14]), .Y(n978) );
  NAND2X0_RVT U1144 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[13]), 
        .Y(n977) );
  NAND3X0_RVT U1145 ( .A1(n978), .A2(n950), .A3(n977), .Y(n979) );
  AOI21X1_RVT U1146 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[13]), 
        .A3(n979), .Y(n665) );
  AOI22X1_RVT U1147 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[13]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[13]), .Y(n981) );
  NAND2X0_RVT U1148 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[12]), 
        .Y(n980) );
  NAND3X0_RVT U1149 ( .A1(n981), .A2(n950), .A3(n980), .Y(n982) );
  AOI21X1_RVT U1150 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[12]), 
        .A3(n982), .Y(n664) );
  AOI22X1_RVT U1151 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[12]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[12]), .Y(n984) );
  NAND2X0_RVT U1152 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[11]), 
        .Y(n983) );
  NAND3X0_RVT U1153 ( .A1(n984), .A2(n950), .A3(n983), .Y(n985) );
  AOI21X1_RVT U1154 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[11]), 
        .A3(n985), .Y(n663) );
  AOI22X1_RVT U1155 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[11]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[11]), .Y(n987) );
  NAND2X0_RVT U1156 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[10]), 
        .Y(n986) );
  NAND3X0_RVT U1157 ( .A1(n987), .A2(n950), .A3(n986), .Y(n988) );
  AOI21X1_RVT U1158 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[10]), 
        .A3(n988), .Y(n662) );
  AOI22X1_RVT U1159 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[10]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[10]), .Y(n990) );
  NAND2X0_RVT U1160 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[9]), 
        .Y(n989) );
  NAND3X0_RVT U1161 ( .A1(n990), .A2(n950), .A3(n989), .Y(n991) );
  AOI21X1_RVT U1162 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[9]), 
        .A3(n991), .Y(n661) );
  AOI22X1_RVT U1163 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[9]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[9]), .Y(n993) );
  NAND2X0_RVT U1164 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[8]), 
        .Y(n992) );
  NAND3X0_RVT U1165 ( .A1(n993), .A2(n950), .A3(n992), .Y(n994) );
  AOI21X1_RVT U1166 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[8]), 
        .A3(n994), .Y(n660) );
  AOI22X1_RVT U1167 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[8]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[8]), .Y(n996) );
  NAND2X0_RVT U1168 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[7]), 
        .Y(n995) );
  NAND3X0_RVT U1169 ( .A1(n996), .A2(n950), .A3(n995), .Y(n997) );
  AOI21X1_RVT U1170 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[7]), 
        .A3(n997), .Y(n659) );
  AOI22X1_RVT U1171 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[7]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[7]), .Y(n999) );
  NAND2X0_RVT U1172 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[6]), 
        .Y(n998) );
  NAND3X0_RVT U1173 ( .A1(n999), .A2(n950), .A3(n998), .Y(n1000) );
  AOI21X1_RVT U1174 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[6]), 
        .A3(n1000), .Y(n658) );
  AOI22X1_RVT U1175 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[6]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[6]), .Y(n1002) );
  NAND2X0_RVT U1176 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[5]), 
        .Y(n1001) );
  NAND3X0_RVT U1177 ( .A1(n1002), .A2(n950), .A3(n1001), .Y(n1003) );
  AOI21X1_RVT U1178 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[5]), 
        .A3(n1003), .Y(n657) );
  AOI22X1_RVT U1179 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[5]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[5]), .Y(n1005) );
  NAND2X0_RVT U1180 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[4]), 
        .Y(n1004) );
  NAND3X0_RVT U1181 ( .A1(n1005), .A2(n950), .A3(n1004), .Y(n1006) );
  AOI21X1_RVT U1182 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[4]), 
        .A3(n1006), .Y(n656) );
  AOI22X1_RVT U1183 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[4]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[4]), .Y(n1008) );
  NAND2X0_RVT U1184 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[3]), 
        .Y(n1007) );
  NAND3X0_RVT U1185 ( .A1(n1008), .A2(n950), .A3(n1007), .Y(n1009) );
  AOI21X1_RVT U1186 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[3]), 
        .A3(n1009), .Y(n655) );
  AOI22X1_RVT U1187 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[3]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[3]), .Y(n1011) );
  NAND2X0_RVT U1188 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[2]), 
        .Y(n1010) );
  NAND3X0_RVT U1189 ( .A1(n1011), .A2(n950), .A3(n1010), .Y(n1012) );
  AOI21X1_RVT U1190 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[2]), 
        .A3(n1012), .Y(n654) );
  AOI22X1_RVT U1191 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[2]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[2]), .Y(n1014) );
  NAND2X0_RVT U1192 ( .A1(div_norm_frac_in1_dbl_dnrm), .A2(div_frac_in1[1]), 
        .Y(n1013) );
  NAND3X0_RVT U1193 ( .A1(n1014), .A2(n950), .A3(n1013), .Y(n1015) );
  AOI21X1_RVT U1194 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[1]), 
        .A3(n1015), .Y(n653) );
  AOI22X1_RVT U1195 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[1]), 
        .A3(div_norm_frac_in1_dbl_dnrm), .A4(div_frac_in1[0]), .Y(n1017) );
  NAND2X0_RVT U1196 ( .A1(div_norm_frac_in1_dbl_norm), .A2(div_frac_in1[1]), 
        .Y(n1016) );
  NAND3X0_RVT U1197 ( .A1(n1017), .A2(n950), .A3(n1016), .Y(n1018) );
  AOI21X1_RVT U1198 ( .A1(div_norm_frac_in2_dbl_dnrm), .A2(div_frac_in2[0]), 
        .A3(n1018), .Y(n652) );
  AO22X1_RVT U1199 ( .A1(div_norm_frac_in2_dbl_norm), .A2(div_frac_in2[0]), 
        .A3(div_norm_frac_in1_dbl_norm), .A4(div_frac_in1[0]), .Y(n1019) );
  NOR2X0_RVT U1200 ( .A1(n1020), .A2(n1019), .Y(n651) );
endmodule


module fpu_div ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_div, 
        fdiv_clken_l, fdiv_clken_l_div_exp_buf1, arst_l, grst_l, rclk, 
        div_pipe_active, d1stg_step, d8stg_fdiv_in, div_id_out_in, div_exc_out, 
        d8stg_fdivd, d8stg_fdivs, div_sign_out, div_exp_outa, div_frac_outa, 
        se, si, so, div_dest_rdy_BAR );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] div_id_out_in;
  output [4:0] div_exc_out;
  output [10:0] div_exp_outa;
  output [51:0] div_frac_outa;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_div, fdiv_clken_l, fdiv_clken_l_div_exp_buf1,
         arst_l, grst_l, rclk, se, si, div_dest_rdy_BAR;
  output div_pipe_active, d1stg_step, d8stg_fdiv_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, so;
  wire   div_dest_rdy, div_frac_add_52_inva, div_frac_add_in1_neq_0,
         d6stg_frac_0, d6stg_frac_1, d6stg_frac_2, d6stg_frac_29,
         d6stg_frac_30, d6stg_frac_31, \div_expadd2[12] , d1stg_snan_sng_in1,
         d1stg_snan_dbl_in1, d1stg_snan_sng_in2, d1stg_snan_dbl_in2,
         d1stg_dblop, d234stg_fdiv, d3stg_fdiv, d4stg_fdiv, d5stg_fdiva,
         d5stg_fdivb, d5stg_fdivs, d5stg_fdivd, d6stg_fdiv, d6stg_fdivs,
         d6stg_fdivd, d7stg_fdivd, div_norm_frac_in1_dbl_norm,
         div_norm_frac_in1_dbl_dnrm, div_norm_frac_in1_sng_norm,
         div_norm_frac_in1_sng_dnrm, div_norm_frac_in2_dbl_norm,
         div_norm_frac_in2_dbl_dnrm, div_norm_frac_in2_sng_norm,
         div_norm_frac_in2_sng_dnrm, div_norm_inf, div_norm_qnan,
         div_frac_add_in2_load, d6stg_frac_out_nosh, div_frac_add_in1_add,
         div_frac_add_in1_load, d7stg_rndup_inv, d7stg_to_0, d7stg_to_0_inv,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, div_frac_out_load,
         div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl,
         div_expadd1_in2_exp_in2_sng, div_exp1_expadd1, div_exp1_0835,
         div_exp1_0118, div_exp1_load, div_expadd2_in1_exp_out,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd22_inv,
         div_exp_out_expadd2, div_exp_out_of, div_exp_out_exp_out,
         div_exp_out_load, div_frac_add_52_inv, net211148, net211149,
         net211150, net211151, net211152, net211153, net211154;
  wire   [12:0] div_exp1;
  wire   [12:0] div_exp_out;
  wire   [54:53] div_frac_out;
  wire   [5:0] div_shl_cnt;
  assign div_dest_rdy = div_dest_rdy_BAR;

  fpu_div_ctl fpu_div_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_51(inq_in2[51]), .inq_in2_54(
        inq_in2[54]), .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(inq_op), .div_exp1(
        div_exp1), .inq_rnd_mode(inq_rnd_mode), .inq_id(inq_id), .inq_in1_63(
        inq_in1[63]), .inq_in2_63(inq_in2[63]), .inq_div(inq_div), 
        .div_exp_out(div_exp_out), .div_frac_add_52_inva(div_frac_add_52_inva), 
        .div_frac_add_in1_neq_0(div_frac_add_in1_neq_0), .div_frac_out_54(
        div_frac_out[54]), .d6stg_frac_0(d6stg_frac_0), .d6stg_frac_1(
        d6stg_frac_1), .d6stg_frac_2(d6stg_frac_2), .d6stg_frac_29(
        d6stg_frac_29), .d6stg_frac_30(d6stg_frac_30), .d6stg_frac_31(
        d6stg_frac_31), .div_frac_out_53(div_frac_out[53]), .div_expadd2_12(
        \div_expadd2[12] ), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), 
        .div_pipe_active(div_pipe_active), .d1stg_snan_sng_in1(
        d1stg_snan_sng_in1), .d1stg_snan_dbl_in1(d1stg_snan_dbl_in1), 
        .d1stg_snan_sng_in2(d1stg_snan_sng_in2), .d1stg_snan_dbl_in2(
        d1stg_snan_dbl_in2), .d1stg_step(d1stg_step), .d1stg_dblop(d1stg_dblop), .d234stg_fdiv(d234stg_fdiv), .d3stg_fdiv(d3stg_fdiv), .d4stg_fdiv(d4stg_fdiv), .d5stg_fdiva(d5stg_fdiva), .d5stg_fdivb(d5stg_fdivb), .d5stg_fdivs(
        d5stg_fdivs), .d5stg_fdivd(d5stg_fdivd), .d6stg_fdiv(d6stg_fdiv), 
        .d6stg_fdivs(d6stg_fdivs), .d6stg_fdivd(d6stg_fdivd), .d7stg_fdivd(
        d7stg_fdivd), .d8stg_fdiv_in(d8stg_fdiv_in), .d8stg_fdivs(d8stg_fdivs), 
        .d8stg_fdivd(d8stg_fdivd), .div_id_out_in(div_id_out_in), 
        .div_sign_out(div_sign_out), .div_exc_out(div_exc_out), 
        .div_norm_frac_in1_dbl_norm(div_norm_frac_in1_dbl_norm), 
        .div_norm_frac_in1_dbl_dnrm(div_norm_frac_in1_dbl_dnrm), 
        .div_norm_frac_in1_sng_norm(div_norm_frac_in1_sng_norm), 
        .div_norm_frac_in1_sng_dnrm(div_norm_frac_in1_sng_dnrm), 
        .div_norm_frac_in2_dbl_norm(div_norm_frac_in2_dbl_norm), 
        .div_norm_frac_in2_dbl_dnrm(div_norm_frac_in2_dbl_dnrm), 
        .div_norm_frac_in2_sng_norm(div_norm_frac_in2_sng_norm), 
        .div_norm_frac_in2_sng_dnrm(div_norm_frac_in2_sng_dnrm), 
        .div_norm_inf(div_norm_inf), .div_norm_qnan(div_norm_qnan), 
        .div_frac_add_in2_load(div_frac_add_in2_load), .d6stg_frac_out_nosh(
        d6stg_frac_out_nosh), .div_frac_add_in1_add(div_frac_add_in1_add), 
        .div_frac_add_in1_load(div_frac_add_in1_load), .d7stg_rndup_inv(
        d7stg_rndup_inv), .d7stg_to_0(d7stg_to_0), .d7stg_to_0_inv(
        d7stg_to_0_inv), .div_frac_out_add_in1(div_frac_out_add_in1), 
        .div_frac_out_add(div_frac_out_add), .div_frac_out_shl1_dbl(
        div_frac_out_shl1_dbl), .div_frac_out_shl1_sng(div_frac_out_shl1_sng), 
        .div_frac_out_of(div_frac_out_of), .div_frac_out_load(
        div_frac_out_load), .div_expadd1_in1_dbl(div_expadd1_in1_dbl), 
        .div_expadd1_in1_sng(div_expadd1_in1_sng), 
        .div_expadd1_in2_exp_in2_dbl(div_expadd1_in2_exp_in2_dbl), 
        .div_expadd1_in2_exp_in2_sng(div_expadd1_in2_exp_in2_sng), 
        .div_exp1_expadd1(div_exp1_expadd1), .div_exp1_0835(div_exp1_0835), 
        .div_exp1_0118(div_exp1_0118), .div_exp1_load(div_exp1_load), 
        .div_expadd2_in1_exp_out(div_expadd2_in1_exp_out), 
        .div_expadd2_no_decr_inv(div_expadd2_no_decr_inv), .div_expadd2_cin(
        div_expadd2_cin), .div_exp_out_expadd22_inv(div_exp_out_expadd22_inv), 
        .div_exp_out_expadd2(div_exp_out_expadd2), .div_exp_out_of(
        div_exp_out_of), .div_exp_out_exp_out(div_exp_out_exp_out), 
        .div_exp_out_load(div_exp_out_load), .se(se), .si(net211154), 
        .div_dest_rdy_BAR(div_dest_rdy) );
  fpu_div_exp_dp fpu_div_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .d1stg_step(d1stg_step), .d234stg_fdiv(d234stg_fdiv), 
        .div_expadd1_in1_dbl(div_expadd1_in1_dbl), .div_expadd1_in1_sng(
        div_expadd1_in1_sng), .div_expadd1_in2_exp_in2_dbl(
        div_expadd1_in2_exp_in2_dbl), .div_expadd1_in2_exp_in2_sng(
        div_expadd1_in2_exp_in2_sng), .d3stg_fdiv(d3stg_fdiv), .d4stg_fdiv(
        d4stg_fdiv), .div_shl_cnt(div_shl_cnt), .div_exp1_expadd1(
        div_exp1_expadd1), .div_exp1_0835(div_exp1_0835), .div_exp1_0118(
        div_exp1_0118), .div_exp1_zero(net211151), .div_exp1_load(
        div_exp1_load), .div_expadd2_in1_exp_out(div_expadd2_in1_exp_out), 
        .d5stg_fdiva(d5stg_fdiva), .d5stg_fdivd(d5stg_fdivd), .d5stg_fdivs(
        d5stg_fdivs), .d6stg_fdiv(d6stg_fdiv), .d7stg_fdiv(net211152), 
        .div_expadd2_no_decr_inv(div_expadd2_no_decr_inv), .div_expadd2_cin(
        div_expadd2_cin), .div_exp_out_expadd2(div_exp_out_expadd2), 
        .div_exp_out_expadd22_inv(div_exp_out_expadd22_inv), .div_exp_out_of(
        div_exp_out_of), .d7stg_to_0_inv(d7stg_to_0_inv), .d7stg_fdivd(
        d7stg_fdivd), .div_exp_out_exp_out(div_exp_out_exp_out), 
        .d7stg_rndup_inv(d7stg_rndup_inv), .div_frac_add_52_inv(
        div_frac_add_52_inv), .div_exp_out_load(div_exp_out_load), 
        .fdiv_clken_l(fdiv_clken_l_div_exp_buf1), .rclk(rclk), .div_exp1(
        div_exp1), .div_expadd2_12(\div_expadd2[12] ), .div_exp_out(
        div_exp_out), .div_exp_outa(div_exp_outa), .se(se), .si(net211153) );
  fpu_div_frac_dp fpu_div_frac_dp ( .inq_in1(inq_in1[54:0]), .inq_in2(
        inq_in2[54:0]), .d1stg_step(d1stg_step), .div_norm_frac_in1_dbl_norm(
        div_norm_frac_in1_dbl_norm), .div_norm_frac_in1_dbl_dnrm(
        div_norm_frac_in1_dbl_dnrm), .div_norm_frac_in1_sng_norm(
        div_norm_frac_in1_sng_norm), .div_norm_frac_in1_sng_dnrm(
        div_norm_frac_in1_sng_dnrm), .div_norm_frac_in2_dbl_norm(
        div_norm_frac_in2_dbl_norm), .div_norm_frac_in2_dbl_dnrm(
        div_norm_frac_in2_dbl_dnrm), .div_norm_frac_in2_sng_norm(
        div_norm_frac_in2_sng_norm), .div_norm_frac_in2_sng_dnrm(
        div_norm_frac_in2_sng_dnrm), .div_norm_inf(div_norm_inf), 
        .div_norm_qnan(div_norm_qnan), .d1stg_dblop(d1stg_dblop), 
        .div_norm_zero(net211148), .d1stg_snan_dbl_in1(d1stg_snan_dbl_in1), 
        .d1stg_snan_sng_in1(d1stg_snan_sng_in1), .d1stg_snan_dbl_in2(
        d1stg_snan_dbl_in2), .d1stg_snan_sng_in2(d1stg_snan_sng_in2), 
        .d3stg_fdiv(d3stg_fdiv), .d6stg_fdiv(d6stg_fdiv), .d6stg_fdivd(
        d6stg_fdivd), .d6stg_fdivs(d6stg_fdivs), .div_frac_add_in2_load(
        div_frac_add_in2_load), .d6stg_frac_out_shl1(net211149), 
        .d6stg_frac_out_nosh(d6stg_frac_out_nosh), .d4stg_fdiv(d4stg_fdiv), 
        .div_frac_add_in1_add(div_frac_add_in1_add), .div_frac_add_in1_load(
        div_frac_add_in1_load), .d5stg_fdivb(d5stg_fdivb), 
        .div_frac_out_add_in1(div_frac_out_add_in1), .div_frac_out_add(
        div_frac_out_add), .div_frac_out_shl1_dbl(div_frac_out_shl1_dbl), 
        .div_frac_out_shl1_sng(div_frac_out_shl1_sng), .div_frac_out_of(
        div_frac_out_of), .d7stg_to_0(d7stg_to_0), .div_frac_out_load(
        div_frac_out_load), .fdiv_clken_l(fdiv_clken_l), .rclk(rclk), 
        .div_shl_cnt(div_shl_cnt), .d6stg_frac_0(d6stg_frac_0), .d6stg_frac_1(
        d6stg_frac_1), .d6stg_frac_2(d6stg_frac_2), .d6stg_frac_29(
        d6stg_frac_29), .d6stg_frac_30(d6stg_frac_30), .d6stg_frac_31(
        d6stg_frac_31), .div_frac_add_in1_neq_0(div_frac_add_in1_neq_0), 
        .div_frac_add_52_inv(div_frac_add_52_inv), .div_frac_add_52_inva(
        div_frac_add_52_inva), .div_frac_out_54_53(div_frac_out), 
        .div_frac_outa(div_frac_outa), .se(se), .si(net211150) );
endmodule


module dffrl_async_SIZE1_1 ( din, clk, rst_l, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  output \q[0]_BAR ;
  wire   N4, n1;

  DFFARX1_RVT \q_reg[0]  ( .D(N4), .CLK(clk), .RSTB(rst_l), .QN(\q[0]_BAR ) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N4) );
endmodule


module dffre_SIZE1_1 ( din, rst, en, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  output \q[0]_BAR ;
  wire   \q[0] , n1, n2, n5;

  DFFX1_RVT \q_reg[0]  ( .D(n5), .CLK(clk), .Q(\q[0] ), .QN(\q[0]_BAR ) );
  INVX1_RVT U2 ( .A(en), .Y(n1) );
  AO22X1_RVT U3 ( .A1(en), .A2(\q[0] ), .A3(n1), .A4(\q[0]_BAR ), .Y(n2) );
  NOR3X0_RVT U4 ( .A1(rst), .A2(se), .A3(n2), .Y(n5) );
endmodule


module dff_SIZE8_2 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, n1;

  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
endmodule


module dff_SIZE2_1 ( din, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input clk, se;
  wire   N3, N4, n1;

  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
endmodule


module dff_SIZE3_0 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N3, N4, N5, n1;

  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
endmodule


module dff_SIZE1_5 ( din, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0]_BAR ;


  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\q[0]_BAR ) );
endmodule


module dff_SIZE1_4 ( din, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0]_BAR ;
  wire   N3, n2;

  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .QN(\q[0]_BAR ) );
  INVX1_RVT U3 ( .A(se), .Y(n2) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n2), .Y(N3) );
endmodule


module dff_SIZE1_3 ( din, clk, se, si, so, \q[0]_BAR  );
  input [0:0] din;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  output \q[0]_BAR ;


  DFFSSRX1_RVT \q_reg[0]  ( .D(1'b0), .SETB(se), .RSTB(din[0]), .CLK(clk), 
        .QN(\q[0]_BAR ) );
endmodule


module fpu_out_ctl ( d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, 
        div_id_out_in, m6stg_id_in, add_id_out_in, arst_l, grst_l, rclk, 
        fp_cpx_req_cq, req_thread, dest_rdy, se, si, so, add_dest_rdy_BAR, 
        div_dest_rdy_BAR, mul_dest_rdy_BAR );
  input [9:0] div_id_out_in;
  input [9:0] m6stg_id_in;
  input [9:0] add_id_out_in;
  output [7:0] fp_cpx_req_cq;
  output [1:0] req_thread;
  output [2:0] dest_rdy;
  input d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, arst_l, grst_l, rclk, se,
         si;
  output so, add_dest_rdy_BAR, div_dest_rdy_BAR, mul_dest_rdy_BAR;
  wire   add_dest_rdy, mul_dest_rdy, div_dest_rdy, out_ctl_rst_l, add_req,
         add_req_step, \dest_rdy_in[0] , n1, n2, n3, n4, n5, n6;
  wire   [9:0] out_id;
  assign add_dest_rdy_BAR = add_dest_rdy;
  assign mul_dest_rdy_BAR = mul_dest_rdy;
  assign div_dest_rdy_BAR = div_dest_rdy;
  assign so = 1'b0;

  dffrl_async_SIZE1_1 dffrl_out_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .se(se), .si(1'b0), .\q[0]_BAR (out_ctl_rst_l) );
  dffre_SIZE1_1 i_add_req ( .din(1'b0), .rst(out_ctl_rst_l), .en(add_req_step), 
        .clk(rclk), .se(se), .si(1'b0), .\q[0]_BAR (add_req) );
  dff_SIZE8_2 i_fp_cpx_req_cq ( .din(out_id[9:2]), .clk(rclk), .q(
        fp_cpx_req_cq), .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  dff_SIZE2_1 i_req_thread ( .din(out_id[1:0]), .clk(rclk), .q(req_thread), 
        .se(se), .si({1'b0, 1'b0}) );
  dff_SIZE3_0 i_dest_rdy ( .din({d8stg_fdiv_in, n6, \dest_rdy_in[0] }), .clk(
        rclk), .q(dest_rdy), .se(se), .si({1'b0, 1'b0, 1'b0}) );
  dff_SIZE1_5 i_add_dest_rdy ( .din(\dest_rdy_in[0] ), .clk(rclk), .se(se), 
        .si(1'b0), .\q[0]_BAR (add_dest_rdy) );
  dff_SIZE1_4 i_mul_dest_rdy ( .din(n6), .clk(rclk), .se(se), .si(1'b0), 
        .\q[0]_BAR (mul_dest_rdy) );
  dff_SIZE1_3 i_div_dest_rdy ( .din(d8stg_fdiv_in), .clk(rclk), .se(se), .si(
        1'b0), .\q[0]_BAR (div_dest_rdy) );
  INVX0_RVT U1 ( .A(add_req), .Y(n3) );
  INVX1_RVT U2 ( .A(d8stg_fdiv_in), .Y(n2) );
  NAND2X0_RVT U3 ( .A1(add_req), .A2(m6stg_fmul_in), .Y(n1) );
  AND3X1_RVT U4 ( .A1(n2), .A2(a6stg_fadd_in), .A3(n1), .Y(\dest_rdy_in[0] )
         );
  AND2X1_RVT U5 ( .A1(n2), .A2(m6stg_fmul_in), .Y(n5) );
  NAND2X0_RVT U6 ( .A1(n3), .A2(a6stg_fadd_in), .Y(n4) );
  AND2X1_RVT U7 ( .A1(n5), .A2(n4), .Y(n6) );
  OR2X1_RVT U10 ( .A1(n6), .A2(\dest_rdy_in[0] ), .Y(add_req_step) );
  AO222X1_RVT U11 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[9]), .A3(n6), .A4(
        m6stg_id_in[9]), .A5(\dest_rdy_in[0] ), .A6(add_id_out_in[9]), .Y(
        out_id[9]) );
  AO222X1_RVT U12 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[8]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[8]), .A5(m6stg_id_in[8]), .A6(n6), 
        .Y(out_id[8]) );
  AO222X1_RVT U13 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[7]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[7]), .A5(m6stg_id_in[7]), .A6(n6), 
        .Y(out_id[7]) );
  AO222X1_RVT U14 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[6]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[6]), .A5(m6stg_id_in[6]), .A6(n6), 
        .Y(out_id[6]) );
  AO222X1_RVT U15 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[5]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[5]), .A5(m6stg_id_in[5]), .A6(n6), 
        .Y(out_id[5]) );
  AO222X1_RVT U16 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[4]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[4]), .A5(m6stg_id_in[4]), .A6(n6), 
        .Y(out_id[4]) );
  AO222X1_RVT U17 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[3]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[3]), .A5(m6stg_id_in[3]), .A6(n6), 
        .Y(out_id[3]) );
  AO222X1_RVT U18 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[2]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[2]), .A5(m6stg_id_in[2]), .A6(n6), 
        .Y(out_id[2]) );
  AO222X1_RVT U19 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[1]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[1]), .A5(m6stg_id_in[1]), .A6(n6), 
        .Y(out_id[1]) );
  AO222X1_RVT U20 ( .A1(d8stg_fdiv_in), .A2(div_id_out_in[0]), .A3(
        \dest_rdy_in[0] ), .A4(add_id_out_in[0]), .A5(m6stg_id_in[0]), .A6(n6), 
        .Y(out_id[0]) );
endmodule


module clken_buf_3 ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   rclk;
  assign clk = rclk;

endmodule


module dff_SIZE8_1 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N3, N4, N9, n1;
  assign q[7] = q[6];

  DFFX1_RVT \q_reg[7]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[6]), .A2(n1), .Y(N9) );
endmodule


module dff_SIZE77 ( din, clk, q, se, si, so );
  input [76:0] din;
  output [76:0] q;
  input [76:0] si;
  output [76:0] so;
  input clk, se;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N68, N69, N70, N71, N72, N75, N76,
         N77, N78, N79, n1, n2, n3, n4, n5;

  DFFX1_RVT \q_reg[76]  ( .D(N79), .CLK(clk), .Q(q[76]) );
  DFFX1_RVT \q_reg[75]  ( .D(N78), .CLK(clk), .Q(q[75]) );
  DFFX1_RVT \q_reg[74]  ( .D(N77), .CLK(clk), .Q(q[74]) );
  DFFX1_RVT \q_reg[73]  ( .D(N76), .CLK(clk), .Q(q[73]) );
  DFFX1_RVT \q_reg[72]  ( .D(N75), .CLK(clk), .Q(q[72]) );
  DFFX1_RVT \q_reg[69]  ( .D(N72), .CLK(clk), .Q(q[69]) );
  DFFX1_RVT \q_reg[68]  ( .D(N71), .CLK(clk), .Q(q[68]) );
  DFFX1_RVT \q_reg[67]  ( .D(N70), .CLK(clk), .Q(q[67]) );
  DFFX1_RVT \q_reg[66]  ( .D(N69), .CLK(clk), .Q(q[66]) );
  DFFX1_RVT \q_reg[65]  ( .D(N68), .CLK(clk), .Q(q[65]) );
  DFFX1_RVT \q_reg[63]  ( .D(N66), .CLK(clk), .Q(q[63]) );
  DFFX1_RVT \q_reg[62]  ( .D(N65), .CLK(clk), .Q(q[62]) );
  DFFX1_RVT \q_reg[61]  ( .D(N64), .CLK(clk), .Q(q[61]) );
  DFFX1_RVT \q_reg[60]  ( .D(N63), .CLK(clk), .Q(q[60]) );
  DFFX1_RVT \q_reg[59]  ( .D(N62), .CLK(clk), .Q(q[59]) );
  DFFX1_RVT \q_reg[58]  ( .D(N61), .CLK(clk), .Q(q[58]) );
  DFFX1_RVT \q_reg[57]  ( .D(N60), .CLK(clk), .Q(q[57]) );
  DFFX1_RVT \q_reg[56]  ( .D(N59), .CLK(clk), .Q(q[56]) );
  DFFX1_RVT \q_reg[55]  ( .D(N58), .CLK(clk), .Q(q[55]) );
  DFFX1_RVT \q_reg[54]  ( .D(N57), .CLK(clk), .Q(q[54]) );
  DFFX1_RVT \q_reg[53]  ( .D(N56), .CLK(clk), .Q(q[53]) );
  DFFX1_RVT \q_reg[52]  ( .D(N55), .CLK(clk), .Q(q[52]) );
  DFFX1_RVT \q_reg[51]  ( .D(N54), .CLK(clk), .Q(q[51]) );
  DFFX1_RVT \q_reg[50]  ( .D(N53), .CLK(clk), .Q(q[50]) );
  DFFX1_RVT \q_reg[49]  ( .D(N52), .CLK(clk), .Q(q[49]) );
  DFFX1_RVT \q_reg[48]  ( .D(N51), .CLK(clk), .Q(q[48]) );
  DFFX1_RVT \q_reg[47]  ( .D(N50), .CLK(clk), .Q(q[47]) );
  DFFX1_RVT \q_reg[46]  ( .D(N49), .CLK(clk), .Q(q[46]) );
  DFFX1_RVT \q_reg[45]  ( .D(N48), .CLK(clk), .Q(q[45]) );
  DFFX1_RVT \q_reg[44]  ( .D(N47), .CLK(clk), .Q(q[44]) );
  DFFX1_RVT \q_reg[43]  ( .D(N46), .CLK(clk), .Q(q[43]) );
  DFFX1_RVT \q_reg[42]  ( .D(N45), .CLK(clk), .Q(q[42]) );
  DFFX1_RVT \q_reg[41]  ( .D(N44), .CLK(clk), .Q(q[41]) );
  DFFX1_RVT \q_reg[40]  ( .D(N43), .CLK(clk), .Q(q[40]) );
  DFFX1_RVT \q_reg[39]  ( .D(N42), .CLK(clk), .Q(q[39]) );
  DFFX1_RVT \q_reg[38]  ( .D(N41), .CLK(clk), .Q(q[38]) );
  DFFX1_RVT \q_reg[37]  ( .D(N40), .CLK(clk), .Q(q[37]) );
  DFFX1_RVT \q_reg[36]  ( .D(N39), .CLK(clk), .Q(q[36]) );
  DFFX1_RVT \q_reg[35]  ( .D(N38), .CLK(clk), .Q(q[35]) );
  DFFX1_RVT \q_reg[34]  ( .D(N37), .CLK(clk), .Q(q[34]) );
  DFFX1_RVT \q_reg[33]  ( .D(N36), .CLK(clk), .Q(q[33]) );
  DFFX1_RVT \q_reg[32]  ( .D(N35), .CLK(clk), .Q(q[32]) );
  DFFX1_RVT \q_reg[31]  ( .D(N34), .CLK(clk), .Q(q[31]) );
  DFFX1_RVT \q_reg[30]  ( .D(N33), .CLK(clk), .Q(q[30]) );
  DFFX1_RVT \q_reg[29]  ( .D(N32), .CLK(clk), .Q(q[29]) );
  DFFX1_RVT \q_reg[28]  ( .D(N31), .CLK(clk), .Q(q[28]) );
  DFFX1_RVT \q_reg[27]  ( .D(N30), .CLK(clk), .Q(q[27]) );
  DFFX1_RVT \q_reg[26]  ( .D(N29), .CLK(clk), .Q(q[26]) );
  DFFX1_RVT \q_reg[25]  ( .D(N28), .CLK(clk), .Q(q[25]) );
  DFFX1_RVT \q_reg[24]  ( .D(N27), .CLK(clk), .Q(q[24]) );
  DFFX1_RVT \q_reg[23]  ( .D(N26), .CLK(clk), .Q(q[23]) );
  DFFX1_RVT \q_reg[22]  ( .D(N25), .CLK(clk), .Q(q[22]) );
  DFFX1_RVT \q_reg[21]  ( .D(N24), .CLK(clk), .Q(q[21]) );
  DFFX1_RVT \q_reg[20]  ( .D(N23), .CLK(clk), .Q(q[20]) );
  DFFX1_RVT \q_reg[19]  ( .D(N22), .CLK(clk), .Q(q[19]) );
  DFFX1_RVT \q_reg[18]  ( .D(N21), .CLK(clk), .Q(q[18]) );
  DFFX1_RVT \q_reg[17]  ( .D(N20), .CLK(clk), .Q(q[17]) );
  DFFX1_RVT \q_reg[16]  ( .D(N19), .CLK(clk), .Q(q[16]) );
  DFFX1_RVT \q_reg[15]  ( .D(N18), .CLK(clk), .Q(q[15]) );
  DFFX1_RVT \q_reg[14]  ( .D(N17), .CLK(clk), .Q(q[14]) );
  DFFX1_RVT \q_reg[13]  ( .D(N16), .CLK(clk), .Q(q[13]) );
  DFFX1_RVT \q_reg[12]  ( .D(N15), .CLK(clk), .Q(q[12]) );
  DFFX1_RVT \q_reg[11]  ( .D(N14), .CLK(clk), .Q(q[11]) );
  DFFX1_RVT \q_reg[10]  ( .D(N13), .CLK(clk), .Q(q[10]) );
  DFFX1_RVT \q_reg[9]  ( .D(N12), .CLK(clk), .Q(q[9]) );
  DFFX1_RVT \q_reg[8]  ( .D(N11), .CLK(clk), .Q(q[8]) );
  DFFX1_RVT \q_reg[7]  ( .D(N10), .CLK(clk), .Q(q[7]) );
  DFFX1_RVT \q_reg[6]  ( .D(N9), .CLK(clk), .Q(q[6]) );
  DFFX1_RVT \q_reg[5]  ( .D(N8), .CLK(clk), .Q(q[5]) );
  DFFX1_RVT \q_reg[4]  ( .D(N7), .CLK(clk), .Q(q[4]) );
  DFFX1_RVT \q_reg[3]  ( .D(N6), .CLK(clk), .Q(q[3]) );
  DFFX1_RVT \q_reg[2]  ( .D(N5), .CLK(clk), .Q(q[2]) );
  DFFX1_RVT \q_reg[1]  ( .D(N4), .CLK(clk), .Q(q[1]) );
  DFFX1_RVT \q_reg[0]  ( .D(N3), .CLK(clk), .Q(q[0]) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND2X1_RVT U4 ( .A1(din[0]), .A2(n1), .Y(N3) );
  AND2X1_RVT U5 ( .A1(din[1]), .A2(n1), .Y(N4) );
  AND2X1_RVT U6 ( .A1(din[2]), .A2(n1), .Y(N5) );
  AND2X1_RVT U7 ( .A1(din[3]), .A2(n1), .Y(N6) );
  AND2X1_RVT U8 ( .A1(din[4]), .A2(n1), .Y(N7) );
  AND2X1_RVT U9 ( .A1(din[5]), .A2(n1), .Y(N8) );
  AND2X1_RVT U10 ( .A1(din[6]), .A2(n1), .Y(N9) );
  AND2X1_RVT U11 ( .A1(din[7]), .A2(n1), .Y(N10) );
  AND2X1_RVT U12 ( .A1(din[8]), .A2(n1), .Y(N11) );
  AND2X1_RVT U13 ( .A1(din[9]), .A2(n1), .Y(N12) );
  AND2X1_RVT U14 ( .A1(din[10]), .A2(n1), .Y(N13) );
  AND2X1_RVT U15 ( .A1(din[11]), .A2(n1), .Y(N14) );
  INVX1_RVT U16 ( .A(se), .Y(n2) );
  AND2X1_RVT U17 ( .A1(din[12]), .A2(n2), .Y(N15) );
  AND2X1_RVT U18 ( .A1(din[13]), .A2(n2), .Y(N16) );
  AND2X1_RVT U19 ( .A1(din[14]), .A2(n2), .Y(N17) );
  AND2X1_RVT U20 ( .A1(din[15]), .A2(n2), .Y(N18) );
  AND2X1_RVT U21 ( .A1(din[16]), .A2(n2), .Y(N19) );
  AND2X1_RVT U22 ( .A1(din[17]), .A2(n2), .Y(N20) );
  AND2X1_RVT U23 ( .A1(din[18]), .A2(n2), .Y(N21) );
  AND2X1_RVT U24 ( .A1(din[19]), .A2(n2), .Y(N22) );
  AND2X1_RVT U25 ( .A1(din[20]), .A2(n2), .Y(N23) );
  AND2X1_RVT U26 ( .A1(din[21]), .A2(n2), .Y(N24) );
  AND2X1_RVT U27 ( .A1(din[22]), .A2(n2), .Y(N25) );
  AND2X1_RVT U28 ( .A1(din[23]), .A2(n2), .Y(N26) );
  INVX1_RVT U29 ( .A(se), .Y(n3) );
  AND2X1_RVT U30 ( .A1(din[24]), .A2(n3), .Y(N27) );
  AND2X1_RVT U31 ( .A1(din[25]), .A2(n3), .Y(N28) );
  AND2X1_RVT U32 ( .A1(din[26]), .A2(n3), .Y(N29) );
  AND2X1_RVT U33 ( .A1(din[27]), .A2(n3), .Y(N30) );
  AND2X1_RVT U34 ( .A1(din[28]), .A2(n3), .Y(N31) );
  AND2X1_RVT U35 ( .A1(din[29]), .A2(n3), .Y(N32) );
  AND2X1_RVT U36 ( .A1(din[30]), .A2(n3), .Y(N33) );
  AND2X1_RVT U37 ( .A1(din[31]), .A2(n3), .Y(N34) );
  AND2X1_RVT U38 ( .A1(din[32]), .A2(n3), .Y(N35) );
  AND2X1_RVT U39 ( .A1(din[33]), .A2(n3), .Y(N36) );
  AND2X1_RVT U40 ( .A1(din[34]), .A2(n3), .Y(N37) );
  AND2X1_RVT U41 ( .A1(din[35]), .A2(n3), .Y(N38) );
  INVX1_RVT U42 ( .A(se), .Y(n4) );
  AND2X1_RVT U43 ( .A1(din[36]), .A2(n4), .Y(N39) );
  AND2X1_RVT U44 ( .A1(din[37]), .A2(n4), .Y(N40) );
  AND2X1_RVT U45 ( .A1(din[38]), .A2(n4), .Y(N41) );
  AND2X1_RVT U46 ( .A1(din[39]), .A2(n4), .Y(N42) );
  AND2X1_RVT U47 ( .A1(din[40]), .A2(n4), .Y(N43) );
  AND2X1_RVT U48 ( .A1(din[41]), .A2(n4), .Y(N44) );
  AND2X1_RVT U49 ( .A1(din[42]), .A2(n4), .Y(N45) );
  AND2X1_RVT U50 ( .A1(din[43]), .A2(n4), .Y(N46) );
  AND2X1_RVT U51 ( .A1(din[44]), .A2(n4), .Y(N47) );
  AND2X1_RVT U52 ( .A1(din[45]), .A2(n4), .Y(N48) );
  AND2X1_RVT U53 ( .A1(din[46]), .A2(n4), .Y(N49) );
  AND2X1_RVT U54 ( .A1(din[47]), .A2(n4), .Y(N50) );
  INVX1_RVT U55 ( .A(se), .Y(n5) );
  AND2X1_RVT U56 ( .A1(din[48]), .A2(n5), .Y(N51) );
  AND2X1_RVT U57 ( .A1(din[49]), .A2(n5), .Y(N52) );
  AND2X1_RVT U58 ( .A1(din[50]), .A2(n5), .Y(N53) );
  AND2X1_RVT U59 ( .A1(din[51]), .A2(n5), .Y(N54) );
  AND2X1_RVT U60 ( .A1(din[52]), .A2(n5), .Y(N55) );
  AND2X1_RVT U61 ( .A1(din[53]), .A2(n5), .Y(N56) );
  AND2X1_RVT U62 ( .A1(din[54]), .A2(n5), .Y(N57) );
  AND2X1_RVT U63 ( .A1(din[55]), .A2(n5), .Y(N58) );
  AND2X1_RVT U64 ( .A1(din[56]), .A2(n5), .Y(N59) );
  AND2X1_RVT U65 ( .A1(din[57]), .A2(n5), .Y(N60) );
  AND2X1_RVT U66 ( .A1(din[58]), .A2(n5), .Y(N61) );
  AND2X1_RVT U67 ( .A1(din[59]), .A2(n5), .Y(N62) );
  AND2X1_RVT U68 ( .A1(din[60]), .A2(n3), .Y(N63) );
  AND2X1_RVT U69 ( .A1(din[61]), .A2(n4), .Y(N64) );
  AND2X1_RVT U70 ( .A1(din[62]), .A2(n5), .Y(N65) );
  AND2X1_RVT U71 ( .A1(din[63]), .A2(n1), .Y(N66) );
  AND2X1_RVT U72 ( .A1(din[65]), .A2(n2), .Y(N68) );
  AND2X1_RVT U73 ( .A1(din[66]), .A2(n3), .Y(N69) );
  AND2X1_RVT U74 ( .A1(din[67]), .A2(n4), .Y(N70) );
  AND2X1_RVT U75 ( .A1(din[68]), .A2(n5), .Y(N71) );
  AND2X1_RVT U76 ( .A1(din[69]), .A2(n1), .Y(N72) );
  AND2X1_RVT U77 ( .A1(din[72]), .A2(n2), .Y(N75) );
  AND2X1_RVT U78 ( .A1(din[73]), .A2(n3), .Y(N76) );
  AND2X1_RVT U79 ( .A1(din[74]), .A2(n4), .Y(N77) );
  AND2X1_RVT U80 ( .A1(din[75]), .A2(n1), .Y(N78) );
  AND2X1_RVT U81 ( .A1(din[76]), .A2(n2), .Y(N79) );
endmodule


module fpu_out_dp ( dest_rdy, req_thread, div_exc_out, d8stg_fdivd, 
        d8stg_fdivs, div_sign_out, div_exp_out, div_frac_out, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, add_exc_out, a6stg_fcmpop, add_cc_out, add_fcc_out, 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        add_sign_out, add_exp_out, add_frac_out, rclk, fp_cpx_data_ca, se, si, 
        so );
  input [2:0] dest_rdy;
  input [1:0] req_thread;
  input [4:0] div_exc_out;
  input [10:0] div_exp_out;
  input [51:0] div_frac_out;
  input [4:0] mul_exc_out;
  input [10:0] mul_exp_out;
  input [51:0] mul_frac_out;
  input [4:0] add_exc_out;
  input [1:0] add_cc_out;
  input [1:0] add_fcc_out;
  input [10:0] add_exp_out;
  input [63:0] add_frac_out;
  output [144:0] fp_cpx_data_ca;
  input d8stg_fdivd, d8stg_fdivs, div_sign_out, m6stg_fmul_dbl_dst,
         m6stg_fmuls, mul_sign_out, a6stg_fcmpop, a6stg_dbl_dst, a6stg_sng_dst,
         a6stg_long_dst, a6stg_int_dst, add_sign_out, rclk, se, si;
  output so;
  wire   fp_cpx_data_ca_144, fp_cpx_data_ca_143, fp_cpx_data_ca_135,
         fp_cpx_data_ca_134, clk, \fp_cpx_data_ca_84_77_in[6] ,
         fp_cpx_data_ca_84_77_in_1, fp_cpx_data_ca_84_77_in_0,
         fp_cpx_data_ca_76_0_in_76, fp_cpx_data_ca_76_0_in_75,
         fp_cpx_data_ca_76_0_in_74, fp_cpx_data_ca_76_0_in_73,
         fp_cpx_data_ca_76_0_in_72, fp_cpx_data_ca_76_0_in_69,
         fp_cpx_data_ca_76_0_in_68, fp_cpx_data_ca_76_0_in_67,
         fp_cpx_data_ca_76_0_in_66, fp_cpx_data_ca_76_0_in_65, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232;
  wire   [63:0] fp_cpx_data_ca_76_0_in;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;
  assign fp_cpx_data_ca[144] = fp_cpx_data_ca_144;
  assign fp_cpx_data_ca[143] = fp_cpx_data_ca_143;
  assign fp_cpx_data_ca[135] = fp_cpx_data_ca_135;
  assign fp_cpx_data_ca[134] = fp_cpx_data_ca_134;
  assign fp_cpx_data_ca[139] = 1'b0;
  assign fp_cpx_data_ca[138] = 1'b0;
  assign fp_cpx_data_ca[137] = 1'b0;
  assign fp_cpx_data_ca[133] = 1'b0;
  assign fp_cpx_data_ca[132] = 1'b0;
  assign fp_cpx_data_ca[131] = 1'b0;
  assign fp_cpx_data_ca[130] = 1'b0;
  assign fp_cpx_data_ca[129] = 1'b0;
  assign fp_cpx_data_ca[128] = 1'b0;
  assign fp_cpx_data_ca[127] = 1'b0;
  assign fp_cpx_data_ca[126] = 1'b0;
  assign fp_cpx_data_ca[125] = 1'b0;
  assign fp_cpx_data_ca[124] = 1'b0;
  assign fp_cpx_data_ca[123] = 1'b0;
  assign fp_cpx_data_ca[122] = 1'b0;
  assign fp_cpx_data_ca[121] = 1'b0;
  assign fp_cpx_data_ca[120] = 1'b0;
  assign fp_cpx_data_ca[119] = 1'b0;
  assign fp_cpx_data_ca[118] = 1'b0;
  assign fp_cpx_data_ca[117] = 1'b0;
  assign fp_cpx_data_ca[116] = 1'b0;
  assign fp_cpx_data_ca[115] = 1'b0;
  assign fp_cpx_data_ca[114] = 1'b0;
  assign fp_cpx_data_ca[113] = 1'b0;
  assign fp_cpx_data_ca[112] = 1'b0;
  assign fp_cpx_data_ca[111] = 1'b0;
  assign fp_cpx_data_ca[110] = 1'b0;
  assign fp_cpx_data_ca[109] = 1'b0;
  assign fp_cpx_data_ca[108] = 1'b0;
  assign fp_cpx_data_ca[107] = 1'b0;
  assign fp_cpx_data_ca[106] = 1'b0;
  assign fp_cpx_data_ca[105] = 1'b0;
  assign fp_cpx_data_ca[104] = 1'b0;
  assign fp_cpx_data_ca[103] = 1'b0;
  assign fp_cpx_data_ca[102] = 1'b0;
  assign fp_cpx_data_ca[101] = 1'b0;
  assign fp_cpx_data_ca[100] = 1'b0;
  assign fp_cpx_data_ca[99] = 1'b0;
  assign fp_cpx_data_ca[98] = 1'b0;
  assign fp_cpx_data_ca[97] = 1'b0;
  assign fp_cpx_data_ca[96] = 1'b0;
  assign fp_cpx_data_ca[95] = 1'b0;
  assign fp_cpx_data_ca[94] = 1'b0;
  assign fp_cpx_data_ca[93] = 1'b0;
  assign fp_cpx_data_ca[92] = 1'b0;
  assign fp_cpx_data_ca[91] = 1'b0;
  assign fp_cpx_data_ca[90] = 1'b0;
  assign fp_cpx_data_ca[89] = 1'b0;
  assign fp_cpx_data_ca[88] = 1'b0;
  assign fp_cpx_data_ca[87] = 1'b0;
  assign fp_cpx_data_ca[86] = 1'b0;
  assign fp_cpx_data_ca[85] = 1'b0;
  assign fp_cpx_data_ca[84] = 1'b0;
  assign fp_cpx_data_ca[83] = 1'b0;
  assign fp_cpx_data_ca[82] = 1'b0;
  assign fp_cpx_data_ca[81] = 1'b0;
  assign fp_cpx_data_ca[80] = 1'b0;
  assign fp_cpx_data_ca[79] = 1'b0;
  assign fp_cpx_data_ca[78] = 1'b0;
  assign fp_cpx_data_ca[77] = 1'b0;
  assign so = 1'b0;

  clken_buf_3 ckbuf_out_dp ( .clk(clk), .rclk(rclk), .enb_l(1'b0), .tmb_l(1'b0) );
  dff_SIZE8_1 i_fp_cpx_data_ca_84_77 ( .din({1'b0, 
        \fp_cpx_data_ca_84_77_in[6] , 1'b0, 1'b0, 1'b0, 1'b0, 
        fp_cpx_data_ca_84_77_in_1, fp_cpx_data_ca_84_77_in_0}), .clk(clk), .q(
        {fp_cpx_data_ca_144, fp_cpx_data_ca_143, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, fp_cpx_data_ca_135, fp_cpx_data_ca_134}), 
        .se(se), .si({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  dff_SIZE77 i_fp_cpx_data_ca_76_0 ( .din({fp_cpx_data_ca_76_0_in_76, 
        fp_cpx_data_ca_76_0_in_75, fp_cpx_data_ca_76_0_in_74, 
        fp_cpx_data_ca_76_0_in_73, fp_cpx_data_ca_76_0_in_72, 1'b0, 1'b0, 
        fp_cpx_data_ca_76_0_in_69, fp_cpx_data_ca_76_0_in_68, 
        fp_cpx_data_ca_76_0_in_67, fp_cpx_data_ca_76_0_in_66, 
        fp_cpx_data_ca_76_0_in_65, 1'b0, fp_cpx_data_ca_76_0_in}), .clk(clk), 
        .q({fp_cpx_data_ca[76:72], SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, fp_cpx_data_ca[69:65], 
        SYNOPSYS_UNCONNECTED__6, fp_cpx_data_ca[63:0]}), .se(se), .si({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  OR3X1_RVT U2 ( .A1(dest_rdy[0]), .A2(dest_rdy[1]), .A3(dest_rdy[2]), .Y(
        \fp_cpx_data_ca_84_77_in[6] ) );
  AND2X1_RVT U5 ( .A1(dest_rdy[2]), .A2(div_exc_out[1]), .Y(
        fp_cpx_data_ca_76_0_in_73) );
  AND2X1_RVT U6 ( .A1(req_thread[1]), .A2(\fp_cpx_data_ca_84_77_in[6] ), .Y(
        fp_cpx_data_ca_84_77_in_1) );
  AND2X1_RVT U7 ( .A1(req_thread[0]), .A2(\fp_cpx_data_ca_84_77_in[6] ), .Y(
        fp_cpx_data_ca_84_77_in_0) );
  AO222X1_RVT U8 ( .A1(dest_rdy[0]), .A2(add_exc_out[4]), .A3(dest_rdy[2]), 
        .A4(div_exc_out[4]), .A5(dest_rdy[1]), .A6(mul_exc_out[4]), .Y(
        fp_cpx_data_ca_76_0_in_76) );
  AO222X1_RVT U9 ( .A1(dest_rdy[0]), .A2(add_exc_out[3]), .A3(dest_rdy[2]), 
        .A4(div_exc_out[3]), .A5(dest_rdy[1]), .A6(mul_exc_out[3]), .Y(
        fp_cpx_data_ca_76_0_in_75) );
  AO222X1_RVT U10 ( .A1(dest_rdy[0]), .A2(add_exc_out[2]), .A3(dest_rdy[2]), 
        .A4(div_exc_out[2]), .A5(dest_rdy[1]), .A6(mul_exc_out[2]), .Y(
        fp_cpx_data_ca_76_0_in_74) );
  AO222X1_RVT U11 ( .A1(dest_rdy[0]), .A2(add_exc_out[0]), .A3(dest_rdy[2]), 
        .A4(div_exc_out[0]), .A5(dest_rdy[1]), .A6(mul_exc_out[0]), .Y(
        fp_cpx_data_ca_76_0_in_72) );
  AND2X1_RVT U12 ( .A1(dest_rdy[0]), .A2(a6stg_fcmpop), .Y(
        fp_cpx_data_ca_76_0_in_69) );
  AND2X1_RVT U13 ( .A1(dest_rdy[0]), .A2(add_cc_out[1]), .Y(
        fp_cpx_data_ca_76_0_in_68) );
  AND2X1_RVT U14 ( .A1(dest_rdy[0]), .A2(add_cc_out[0]), .Y(
        fp_cpx_data_ca_76_0_in_67) );
  AND2X1_RVT U15 ( .A1(dest_rdy[0]), .A2(add_fcc_out[1]), .Y(
        fp_cpx_data_ca_76_0_in_66) );
  AND2X1_RVT U16 ( .A1(dest_rdy[0]), .A2(add_fcc_out[0]), .Y(
        fp_cpx_data_ca_76_0_in_65) );
  AND2X1_RVT U17 ( .A1(dest_rdy[0]), .A2(a6stg_dbl_dst), .Y(n228) );
  AND2X1_RVT U18 ( .A1(dest_rdy[0]), .A2(a6stg_sng_dst), .Y(n158) );
  AND2X1_RVT U19 ( .A1(dest_rdy[1]), .A2(m6stg_fmul_dbl_dst), .Y(n227) );
  AND2X1_RVT U20 ( .A1(dest_rdy[1]), .A2(m6stg_fmuls), .Y(n157) );
  OA21X1_RVT U21 ( .A1(a6stg_long_dst), .A2(a6stg_int_dst), .A3(dest_rdy[0]), 
        .Y(n159) );
  NAND2X0_RVT U22 ( .A1(dest_rdy[2]), .A2(d8stg_fdivd), .Y(n4) );
  NAND2X0_RVT U23 ( .A1(dest_rdy[2]), .A2(d8stg_fdivs), .Y(n5) );
  NAND2X0_RVT U24 ( .A1(n4), .A2(n5), .Y(n1) );
  AO22X1_RVT U25 ( .A1(add_frac_out[63]), .A2(n159), .A3(div_sign_out), .A4(n1), .Y(n2) );
  AO221X1_RVT U26 ( .A1(mul_sign_out), .A2(n227), .A3(mul_sign_out), .A4(n157), 
        .A5(n2), .Y(n3) );
  AO221X1_RVT U27 ( .A1(add_sign_out), .A2(n228), .A3(add_sign_out), .A4(n158), 
        .A5(n3), .Y(fp_cpx_data_ca_76_0_in[63]) );
  INVX1_RVT U28 ( .A(n4), .Y(n230) );
  INVX1_RVT U29 ( .A(n5), .Y(n156) );
  AO22X1_RVT U30 ( .A1(n230), .A2(div_exp_out[10]), .A3(n156), .A4(
        div_exp_out[7]), .Y(n10) );
  AOI22X1_RVT U31 ( .A1(n158), .A2(add_exp_out[7]), .A3(n157), .A4(
        mul_exp_out[7]), .Y(n8) );
  AOI22X1_RVT U32 ( .A1(n228), .A2(add_exp_out[10]), .A3(n227), .A4(
        mul_exp_out[10]), .Y(n7) );
  NAND2X0_RVT U33 ( .A1(add_frac_out[62]), .A2(n159), .Y(n6) );
  NAND3X0_RVT U34 ( .A1(n8), .A2(n7), .A3(n6), .Y(n9) );
  OR2X1_RVT U35 ( .A1(n10), .A2(n9), .Y(fp_cpx_data_ca_76_0_in[62]) );
  AO22X1_RVT U36 ( .A1(n230), .A2(div_exp_out[9]), .A3(n156), .A4(
        div_exp_out[6]), .Y(n15) );
  AOI22X1_RVT U37 ( .A1(n158), .A2(add_exp_out[6]), .A3(n157), .A4(
        mul_exp_out[6]), .Y(n13) );
  AOI22X1_RVT U38 ( .A1(n228), .A2(add_exp_out[9]), .A3(n227), .A4(
        mul_exp_out[9]), .Y(n12) );
  NAND2X0_RVT U39 ( .A1(add_frac_out[61]), .A2(n159), .Y(n11) );
  NAND3X0_RVT U40 ( .A1(n13), .A2(n12), .A3(n11), .Y(n14) );
  OR2X1_RVT U41 ( .A1(n15), .A2(n14), .Y(fp_cpx_data_ca_76_0_in[61]) );
  AO22X1_RVT U42 ( .A1(n230), .A2(div_exp_out[8]), .A3(n156), .A4(
        div_exp_out[5]), .Y(n20) );
  AOI22X1_RVT U43 ( .A1(n158), .A2(add_exp_out[5]), .A3(n157), .A4(
        mul_exp_out[5]), .Y(n18) );
  AOI22X1_RVT U44 ( .A1(n228), .A2(add_exp_out[8]), .A3(n227), .A4(
        mul_exp_out[8]), .Y(n17) );
  NAND2X0_RVT U45 ( .A1(add_frac_out[60]), .A2(n159), .Y(n16) );
  NAND3X0_RVT U46 ( .A1(n18), .A2(n17), .A3(n16), .Y(n19) );
  OR2X1_RVT U47 ( .A1(n20), .A2(n19), .Y(fp_cpx_data_ca_76_0_in[60]) );
  AO22X1_RVT U48 ( .A1(n230), .A2(div_exp_out[7]), .A3(n156), .A4(
        div_exp_out[4]), .Y(n25) );
  AOI22X1_RVT U49 ( .A1(n158), .A2(add_exp_out[4]), .A3(n157), .A4(
        mul_exp_out[4]), .Y(n23) );
  AOI22X1_RVT U50 ( .A1(n228), .A2(add_exp_out[7]), .A3(n227), .A4(
        mul_exp_out[7]), .Y(n22) );
  NAND2X0_RVT U51 ( .A1(add_frac_out[59]), .A2(n159), .Y(n21) );
  NAND3X0_RVT U52 ( .A1(n23), .A2(n22), .A3(n21), .Y(n24) );
  OR2X1_RVT U53 ( .A1(n25), .A2(n24), .Y(fp_cpx_data_ca_76_0_in[59]) );
  AO22X1_RVT U54 ( .A1(n230), .A2(div_exp_out[6]), .A3(n156), .A4(
        div_exp_out[3]), .Y(n30) );
  AOI22X1_RVT U55 ( .A1(n158), .A2(add_exp_out[3]), .A3(n157), .A4(
        mul_exp_out[3]), .Y(n28) );
  AOI22X1_RVT U56 ( .A1(n228), .A2(add_exp_out[6]), .A3(n227), .A4(
        mul_exp_out[6]), .Y(n27) );
  NAND2X0_RVT U57 ( .A1(add_frac_out[58]), .A2(n159), .Y(n26) );
  NAND3X0_RVT U58 ( .A1(n28), .A2(n27), .A3(n26), .Y(n29) );
  OR2X1_RVT U59 ( .A1(n30), .A2(n29), .Y(fp_cpx_data_ca_76_0_in[58]) );
  AO22X1_RVT U60 ( .A1(n230), .A2(div_exp_out[5]), .A3(n156), .A4(
        div_exp_out[2]), .Y(n35) );
  AOI22X1_RVT U61 ( .A1(n158), .A2(add_exp_out[2]), .A3(n157), .A4(
        mul_exp_out[2]), .Y(n33) );
  AOI22X1_RVT U62 ( .A1(n228), .A2(add_exp_out[5]), .A3(n227), .A4(
        mul_exp_out[5]), .Y(n32) );
  NAND2X0_RVT U63 ( .A1(add_frac_out[57]), .A2(n159), .Y(n31) );
  NAND3X0_RVT U64 ( .A1(n33), .A2(n32), .A3(n31), .Y(n34) );
  OR2X1_RVT U65 ( .A1(n35), .A2(n34), .Y(fp_cpx_data_ca_76_0_in[57]) );
  AO22X1_RVT U66 ( .A1(n230), .A2(div_exp_out[4]), .A3(n156), .A4(
        div_exp_out[1]), .Y(n40) );
  AOI22X1_RVT U67 ( .A1(n158), .A2(add_exp_out[1]), .A3(n157), .A4(
        mul_exp_out[1]), .Y(n38) );
  AOI22X1_RVT U68 ( .A1(n228), .A2(add_exp_out[4]), .A3(n227), .A4(
        mul_exp_out[4]), .Y(n37) );
  NAND2X0_RVT U69 ( .A1(add_frac_out[56]), .A2(n159), .Y(n36) );
  NAND3X0_RVT U70 ( .A1(n38), .A2(n37), .A3(n36), .Y(n39) );
  OR2X1_RVT U71 ( .A1(n40), .A2(n39), .Y(fp_cpx_data_ca_76_0_in[56]) );
  AO22X1_RVT U72 ( .A1(n230), .A2(div_exp_out[3]), .A3(n156), .A4(
        div_exp_out[0]), .Y(n45) );
  AOI22X1_RVT U73 ( .A1(n158), .A2(add_exp_out[0]), .A3(n157), .A4(
        mul_exp_out[0]), .Y(n43) );
  AOI22X1_RVT U74 ( .A1(n228), .A2(add_exp_out[3]), .A3(n227), .A4(
        mul_exp_out[3]), .Y(n42) );
  NAND2X0_RVT U75 ( .A1(add_frac_out[55]), .A2(n159), .Y(n41) );
  NAND3X0_RVT U76 ( .A1(n43), .A2(n42), .A3(n41), .Y(n44) );
  OR2X1_RVT U77 ( .A1(n45), .A2(n44), .Y(fp_cpx_data_ca_76_0_in[55]) );
  AO22X1_RVT U78 ( .A1(n230), .A2(div_exp_out[2]), .A3(n156), .A4(
        div_frac_out[51]), .Y(n50) );
  AOI22X1_RVT U79 ( .A1(n158), .A2(add_frac_out[62]), .A3(n157), .A4(
        mul_frac_out[51]), .Y(n48) );
  AOI22X1_RVT U80 ( .A1(n228), .A2(add_exp_out[2]), .A3(n227), .A4(
        mul_exp_out[2]), .Y(n47) );
  NAND2X0_RVT U81 ( .A1(add_frac_out[54]), .A2(n159), .Y(n46) );
  NAND3X0_RVT U82 ( .A1(n48), .A2(n47), .A3(n46), .Y(n49) );
  OR2X1_RVT U83 ( .A1(n50), .A2(n49), .Y(fp_cpx_data_ca_76_0_in[54]) );
  AO22X1_RVT U84 ( .A1(n230), .A2(div_exp_out[1]), .A3(n156), .A4(
        div_frac_out[50]), .Y(n55) );
  AOI22X1_RVT U85 ( .A1(n158), .A2(add_frac_out[61]), .A3(n157), .A4(
        mul_frac_out[50]), .Y(n53) );
  AOI22X1_RVT U86 ( .A1(n228), .A2(add_exp_out[1]), .A3(n227), .A4(
        mul_exp_out[1]), .Y(n52) );
  NAND2X0_RVT U87 ( .A1(add_frac_out[53]), .A2(n159), .Y(n51) );
  NAND3X0_RVT U88 ( .A1(n53), .A2(n52), .A3(n51), .Y(n54) );
  OR2X1_RVT U89 ( .A1(n55), .A2(n54), .Y(fp_cpx_data_ca_76_0_in[53]) );
  AO22X1_RVT U90 ( .A1(n230), .A2(div_exp_out[0]), .A3(n156), .A4(
        div_frac_out[49]), .Y(n60) );
  AOI22X1_RVT U91 ( .A1(n158), .A2(add_frac_out[60]), .A3(n157), .A4(
        mul_frac_out[49]), .Y(n58) );
  AOI22X1_RVT U92 ( .A1(n228), .A2(add_exp_out[0]), .A3(n227), .A4(
        mul_exp_out[0]), .Y(n57) );
  NAND2X0_RVT U93 ( .A1(add_frac_out[52]), .A2(n159), .Y(n56) );
  NAND3X0_RVT U94 ( .A1(n58), .A2(n57), .A3(n56), .Y(n59) );
  OR2X1_RVT U95 ( .A1(n60), .A2(n59), .Y(fp_cpx_data_ca_76_0_in[52]) );
  AO22X1_RVT U96 ( .A1(n230), .A2(div_frac_out[51]), .A3(n156), .A4(
        div_frac_out[48]), .Y(n65) );
  AOI22X1_RVT U97 ( .A1(n158), .A2(add_frac_out[59]), .A3(n157), .A4(
        mul_frac_out[48]), .Y(n63) );
  AOI22X1_RVT U98 ( .A1(n228), .A2(add_frac_out[62]), .A3(n227), .A4(
        mul_frac_out[51]), .Y(n62) );
  NAND2X0_RVT U99 ( .A1(add_frac_out[51]), .A2(n159), .Y(n61) );
  NAND3X0_RVT U100 ( .A1(n63), .A2(n62), .A3(n61), .Y(n64) );
  OR2X1_RVT U101 ( .A1(n65), .A2(n64), .Y(fp_cpx_data_ca_76_0_in[51]) );
  AO22X1_RVT U102 ( .A1(n230), .A2(div_frac_out[50]), .A3(n156), .A4(
        div_frac_out[47]), .Y(n70) );
  AOI22X1_RVT U103 ( .A1(n158), .A2(add_frac_out[58]), .A3(n157), .A4(
        mul_frac_out[47]), .Y(n68) );
  AOI22X1_RVT U104 ( .A1(n228), .A2(add_frac_out[61]), .A3(n227), .A4(
        mul_frac_out[50]), .Y(n67) );
  NAND2X0_RVT U105 ( .A1(add_frac_out[50]), .A2(n159), .Y(n66) );
  NAND3X0_RVT U106 ( .A1(n68), .A2(n67), .A3(n66), .Y(n69) );
  OR2X1_RVT U107 ( .A1(n70), .A2(n69), .Y(fp_cpx_data_ca_76_0_in[50]) );
  AO22X1_RVT U108 ( .A1(n230), .A2(div_frac_out[49]), .A3(n156), .A4(
        div_frac_out[46]), .Y(n75) );
  AOI22X1_RVT U109 ( .A1(n158), .A2(add_frac_out[57]), .A3(n157), .A4(
        mul_frac_out[46]), .Y(n73) );
  AOI22X1_RVT U110 ( .A1(n228), .A2(add_frac_out[60]), .A3(n227), .A4(
        mul_frac_out[49]), .Y(n72) );
  NAND2X0_RVT U111 ( .A1(add_frac_out[49]), .A2(n159), .Y(n71) );
  NAND3X0_RVT U112 ( .A1(n73), .A2(n72), .A3(n71), .Y(n74) );
  OR2X1_RVT U113 ( .A1(n75), .A2(n74), .Y(fp_cpx_data_ca_76_0_in[49]) );
  AO22X1_RVT U114 ( .A1(n230), .A2(div_frac_out[48]), .A3(n156), .A4(
        div_frac_out[45]), .Y(n80) );
  AOI22X1_RVT U115 ( .A1(n158), .A2(add_frac_out[56]), .A3(n157), .A4(
        mul_frac_out[45]), .Y(n78) );
  AOI22X1_RVT U116 ( .A1(n228), .A2(add_frac_out[59]), .A3(n227), .A4(
        mul_frac_out[48]), .Y(n77) );
  NAND2X0_RVT U117 ( .A1(add_frac_out[48]), .A2(n159), .Y(n76) );
  NAND3X0_RVT U118 ( .A1(n78), .A2(n77), .A3(n76), .Y(n79) );
  OR2X1_RVT U119 ( .A1(n80), .A2(n79), .Y(fp_cpx_data_ca_76_0_in[48]) );
  AO22X1_RVT U120 ( .A1(n230), .A2(div_frac_out[47]), .A3(n156), .A4(
        div_frac_out[44]), .Y(n85) );
  AOI22X1_RVT U121 ( .A1(n158), .A2(add_frac_out[55]), .A3(n157), .A4(
        mul_frac_out[44]), .Y(n83) );
  AOI22X1_RVT U122 ( .A1(n228), .A2(add_frac_out[58]), .A3(n227), .A4(
        mul_frac_out[47]), .Y(n82) );
  NAND2X0_RVT U123 ( .A1(add_frac_out[47]), .A2(n159), .Y(n81) );
  NAND3X0_RVT U124 ( .A1(n83), .A2(n82), .A3(n81), .Y(n84) );
  OR2X1_RVT U125 ( .A1(n85), .A2(n84), .Y(fp_cpx_data_ca_76_0_in[47]) );
  AO22X1_RVT U126 ( .A1(n230), .A2(div_frac_out[46]), .A3(n156), .A4(
        div_frac_out[43]), .Y(n90) );
  AOI22X1_RVT U127 ( .A1(n158), .A2(add_frac_out[54]), .A3(n157), .A4(
        mul_frac_out[43]), .Y(n88) );
  AOI22X1_RVT U128 ( .A1(n228), .A2(add_frac_out[57]), .A3(n227), .A4(
        mul_frac_out[46]), .Y(n87) );
  NAND2X0_RVT U129 ( .A1(add_frac_out[46]), .A2(n159), .Y(n86) );
  NAND3X0_RVT U130 ( .A1(n88), .A2(n87), .A3(n86), .Y(n89) );
  OR2X1_RVT U131 ( .A1(n90), .A2(n89), .Y(fp_cpx_data_ca_76_0_in[46]) );
  AO22X1_RVT U132 ( .A1(n230), .A2(div_frac_out[45]), .A3(n156), .A4(
        div_frac_out[42]), .Y(n95) );
  AOI22X1_RVT U133 ( .A1(n158), .A2(add_frac_out[53]), .A3(n157), .A4(
        mul_frac_out[42]), .Y(n93) );
  AOI22X1_RVT U134 ( .A1(n228), .A2(add_frac_out[56]), .A3(n227), .A4(
        mul_frac_out[45]), .Y(n92) );
  NAND2X0_RVT U135 ( .A1(add_frac_out[45]), .A2(n159), .Y(n91) );
  NAND3X0_RVT U136 ( .A1(n93), .A2(n92), .A3(n91), .Y(n94) );
  OR2X1_RVT U137 ( .A1(n95), .A2(n94), .Y(fp_cpx_data_ca_76_0_in[45]) );
  AO22X1_RVT U138 ( .A1(n230), .A2(div_frac_out[44]), .A3(n156), .A4(
        div_frac_out[41]), .Y(n100) );
  AOI22X1_RVT U139 ( .A1(n158), .A2(add_frac_out[52]), .A3(n157), .A4(
        mul_frac_out[41]), .Y(n98) );
  AOI22X1_RVT U140 ( .A1(n228), .A2(add_frac_out[55]), .A3(n227), .A4(
        mul_frac_out[44]), .Y(n97) );
  NAND2X0_RVT U141 ( .A1(add_frac_out[44]), .A2(n159), .Y(n96) );
  NAND3X0_RVT U142 ( .A1(n98), .A2(n97), .A3(n96), .Y(n99) );
  OR2X1_RVT U143 ( .A1(n100), .A2(n99), .Y(fp_cpx_data_ca_76_0_in[44]) );
  AO22X1_RVT U144 ( .A1(n230), .A2(div_frac_out[43]), .A3(n156), .A4(
        div_frac_out[40]), .Y(n105) );
  AOI22X1_RVT U145 ( .A1(n158), .A2(add_frac_out[51]), .A3(n157), .A4(
        mul_frac_out[40]), .Y(n103) );
  AOI22X1_RVT U146 ( .A1(n228), .A2(add_frac_out[54]), .A3(n227), .A4(
        mul_frac_out[43]), .Y(n102) );
  NAND2X0_RVT U147 ( .A1(add_frac_out[43]), .A2(n159), .Y(n101) );
  NAND3X0_RVT U148 ( .A1(n103), .A2(n102), .A3(n101), .Y(n104) );
  OR2X1_RVT U149 ( .A1(n105), .A2(n104), .Y(fp_cpx_data_ca_76_0_in[43]) );
  AO22X1_RVT U150 ( .A1(n230), .A2(div_frac_out[42]), .A3(n156), .A4(
        div_frac_out[39]), .Y(n110) );
  AOI22X1_RVT U151 ( .A1(n158), .A2(add_frac_out[50]), .A3(n157), .A4(
        mul_frac_out[39]), .Y(n108) );
  AOI22X1_RVT U152 ( .A1(n228), .A2(add_frac_out[53]), .A3(n227), .A4(
        mul_frac_out[42]), .Y(n107) );
  NAND2X0_RVT U153 ( .A1(add_frac_out[42]), .A2(n159), .Y(n106) );
  NAND3X0_RVT U154 ( .A1(n108), .A2(n107), .A3(n106), .Y(n109) );
  OR2X1_RVT U155 ( .A1(n110), .A2(n109), .Y(fp_cpx_data_ca_76_0_in[42]) );
  AO22X1_RVT U156 ( .A1(n230), .A2(div_frac_out[41]), .A3(n156), .A4(
        div_frac_out[38]), .Y(n115) );
  AOI22X1_RVT U157 ( .A1(n158), .A2(add_frac_out[49]), .A3(n157), .A4(
        mul_frac_out[38]), .Y(n113) );
  AOI22X1_RVT U158 ( .A1(n228), .A2(add_frac_out[52]), .A3(n227), .A4(
        mul_frac_out[41]), .Y(n112) );
  NAND2X0_RVT U159 ( .A1(add_frac_out[41]), .A2(n159), .Y(n111) );
  NAND3X0_RVT U160 ( .A1(n113), .A2(n112), .A3(n111), .Y(n114) );
  OR2X1_RVT U161 ( .A1(n115), .A2(n114), .Y(fp_cpx_data_ca_76_0_in[41]) );
  AO22X1_RVT U162 ( .A1(n230), .A2(div_frac_out[40]), .A3(n156), .A4(
        div_frac_out[37]), .Y(n120) );
  AOI22X1_RVT U163 ( .A1(n158), .A2(add_frac_out[48]), .A3(n157), .A4(
        mul_frac_out[37]), .Y(n118) );
  AOI22X1_RVT U164 ( .A1(n228), .A2(add_frac_out[51]), .A3(n227), .A4(
        mul_frac_out[40]), .Y(n117) );
  NAND2X0_RVT U165 ( .A1(add_frac_out[40]), .A2(n159), .Y(n116) );
  NAND3X0_RVT U166 ( .A1(n118), .A2(n117), .A3(n116), .Y(n119) );
  OR2X1_RVT U167 ( .A1(n120), .A2(n119), .Y(fp_cpx_data_ca_76_0_in[40]) );
  AO22X1_RVT U168 ( .A1(n230), .A2(div_frac_out[39]), .A3(n156), .A4(
        div_frac_out[36]), .Y(n125) );
  AOI22X1_RVT U169 ( .A1(n158), .A2(add_frac_out[47]), .A3(n157), .A4(
        mul_frac_out[36]), .Y(n123) );
  AOI22X1_RVT U170 ( .A1(n228), .A2(add_frac_out[50]), .A3(n227), .A4(
        mul_frac_out[39]), .Y(n122) );
  NAND2X0_RVT U171 ( .A1(add_frac_out[39]), .A2(n159), .Y(n121) );
  NAND3X0_RVT U172 ( .A1(n123), .A2(n122), .A3(n121), .Y(n124) );
  OR2X1_RVT U173 ( .A1(n125), .A2(n124), .Y(fp_cpx_data_ca_76_0_in[39]) );
  AO22X1_RVT U174 ( .A1(n230), .A2(div_frac_out[38]), .A3(n156), .A4(
        div_frac_out[35]), .Y(n130) );
  AOI22X1_RVT U175 ( .A1(n158), .A2(add_frac_out[46]), .A3(n157), .A4(
        mul_frac_out[35]), .Y(n128) );
  AOI22X1_RVT U176 ( .A1(n228), .A2(add_frac_out[49]), .A3(n227), .A4(
        mul_frac_out[38]), .Y(n127) );
  NAND2X0_RVT U177 ( .A1(add_frac_out[38]), .A2(n159), .Y(n126) );
  NAND3X0_RVT U178 ( .A1(n128), .A2(n127), .A3(n126), .Y(n129) );
  OR2X1_RVT U179 ( .A1(n130), .A2(n129), .Y(fp_cpx_data_ca_76_0_in[38]) );
  AO22X1_RVT U180 ( .A1(n230), .A2(div_frac_out[37]), .A3(n156), .A4(
        div_frac_out[34]), .Y(n135) );
  AOI22X1_RVT U181 ( .A1(n158), .A2(add_frac_out[45]), .A3(n157), .A4(
        mul_frac_out[34]), .Y(n133) );
  AOI22X1_RVT U182 ( .A1(n228), .A2(add_frac_out[48]), .A3(n227), .A4(
        mul_frac_out[37]), .Y(n132) );
  NAND2X0_RVT U183 ( .A1(add_frac_out[37]), .A2(n159), .Y(n131) );
  NAND3X0_RVT U184 ( .A1(n133), .A2(n132), .A3(n131), .Y(n134) );
  OR2X1_RVT U185 ( .A1(n135), .A2(n134), .Y(fp_cpx_data_ca_76_0_in[37]) );
  AO22X1_RVT U186 ( .A1(n230), .A2(div_frac_out[36]), .A3(n156), .A4(
        div_frac_out[33]), .Y(n140) );
  AOI22X1_RVT U187 ( .A1(n158), .A2(add_frac_out[44]), .A3(n157), .A4(
        mul_frac_out[33]), .Y(n138) );
  AOI22X1_RVT U188 ( .A1(n228), .A2(add_frac_out[47]), .A3(n227), .A4(
        mul_frac_out[36]), .Y(n137) );
  NAND2X0_RVT U189 ( .A1(add_frac_out[36]), .A2(n159), .Y(n136) );
  NAND3X0_RVT U190 ( .A1(n138), .A2(n137), .A3(n136), .Y(n139) );
  OR2X1_RVT U191 ( .A1(n140), .A2(n139), .Y(fp_cpx_data_ca_76_0_in[36]) );
  AO22X1_RVT U192 ( .A1(n230), .A2(div_frac_out[35]), .A3(n156), .A4(
        div_frac_out[32]), .Y(n145) );
  AOI22X1_RVT U193 ( .A1(n158), .A2(add_frac_out[43]), .A3(n157), .A4(
        mul_frac_out[32]), .Y(n143) );
  AOI22X1_RVT U194 ( .A1(n228), .A2(add_frac_out[46]), .A3(n227), .A4(
        mul_frac_out[35]), .Y(n142) );
  NAND2X0_RVT U195 ( .A1(add_frac_out[35]), .A2(n159), .Y(n141) );
  NAND3X0_RVT U196 ( .A1(n143), .A2(n142), .A3(n141), .Y(n144) );
  OR2X1_RVT U197 ( .A1(n145), .A2(n144), .Y(fp_cpx_data_ca_76_0_in[35]) );
  AO22X1_RVT U198 ( .A1(n230), .A2(div_frac_out[34]), .A3(n156), .A4(
        div_frac_out[31]), .Y(n150) );
  AOI22X1_RVT U199 ( .A1(n158), .A2(add_frac_out[42]), .A3(n157), .A4(
        mul_frac_out[31]), .Y(n148) );
  AOI22X1_RVT U200 ( .A1(n228), .A2(add_frac_out[45]), .A3(n227), .A4(
        mul_frac_out[34]), .Y(n147) );
  NAND2X0_RVT U201 ( .A1(add_frac_out[34]), .A2(n159), .Y(n146) );
  NAND3X0_RVT U202 ( .A1(n148), .A2(n147), .A3(n146), .Y(n149) );
  OR2X1_RVT U203 ( .A1(n150), .A2(n149), .Y(fp_cpx_data_ca_76_0_in[34]) );
  AO22X1_RVT U204 ( .A1(n230), .A2(div_frac_out[33]), .A3(n156), .A4(
        div_frac_out[30]), .Y(n155) );
  AOI22X1_RVT U205 ( .A1(n158), .A2(add_frac_out[41]), .A3(n157), .A4(
        mul_frac_out[30]), .Y(n153) );
  AOI22X1_RVT U206 ( .A1(n228), .A2(add_frac_out[44]), .A3(n227), .A4(
        mul_frac_out[33]), .Y(n152) );
  NAND2X0_RVT U207 ( .A1(add_frac_out[33]), .A2(n159), .Y(n151) );
  NAND3X0_RVT U208 ( .A1(n153), .A2(n152), .A3(n151), .Y(n154) );
  OR2X1_RVT U209 ( .A1(n155), .A2(n154), .Y(fp_cpx_data_ca_76_0_in[33]) );
  AO22X1_RVT U210 ( .A1(n230), .A2(div_frac_out[32]), .A3(n156), .A4(
        div_frac_out[29]), .Y(n164) );
  AOI22X1_RVT U211 ( .A1(n158), .A2(add_frac_out[40]), .A3(n157), .A4(
        mul_frac_out[29]), .Y(n162) );
  AOI22X1_RVT U212 ( .A1(n228), .A2(add_frac_out[43]), .A3(n227), .A4(
        mul_frac_out[32]), .Y(n161) );
  NAND2X0_RVT U213 ( .A1(add_frac_out[32]), .A2(n159), .Y(n160) );
  NAND3X0_RVT U214 ( .A1(n162), .A2(n161), .A3(n160), .Y(n163) );
  OR2X1_RVT U215 ( .A1(n164), .A2(n163), .Y(fp_cpx_data_ca_76_0_in[32]) );
  AO22X1_RVT U216 ( .A1(n228), .A2(add_frac_out[42]), .A3(n227), .A4(
        mul_frac_out[31]), .Y(n166) );
  AND2X1_RVT U217 ( .A1(dest_rdy[0]), .A2(a6stg_long_dst), .Y(n229) );
  AO22X1_RVT U218 ( .A1(n230), .A2(div_frac_out[31]), .A3(n229), .A4(
        add_frac_out[31]), .Y(n165) );
  OR2X1_RVT U219 ( .A1(n166), .A2(n165), .Y(fp_cpx_data_ca_76_0_in[31]) );
  AO22X1_RVT U220 ( .A1(n228), .A2(add_frac_out[41]), .A3(n227), .A4(
        mul_frac_out[30]), .Y(n168) );
  AO22X1_RVT U221 ( .A1(n230), .A2(div_frac_out[30]), .A3(n229), .A4(
        add_frac_out[30]), .Y(n167) );
  OR2X1_RVT U222 ( .A1(n168), .A2(n167), .Y(fp_cpx_data_ca_76_0_in[30]) );
  AO22X1_RVT U223 ( .A1(n228), .A2(add_frac_out[40]), .A3(n227), .A4(
        mul_frac_out[29]), .Y(n170) );
  AO22X1_RVT U224 ( .A1(n230), .A2(div_frac_out[29]), .A3(n229), .A4(
        add_frac_out[29]), .Y(n169) );
  OR2X1_RVT U225 ( .A1(n170), .A2(n169), .Y(fp_cpx_data_ca_76_0_in[29]) );
  AO22X1_RVT U226 ( .A1(n228), .A2(add_frac_out[39]), .A3(n227), .A4(
        mul_frac_out[28]), .Y(n172) );
  AO22X1_RVT U227 ( .A1(n230), .A2(div_frac_out[28]), .A3(n229), .A4(
        add_frac_out[28]), .Y(n171) );
  OR2X1_RVT U228 ( .A1(n172), .A2(n171), .Y(fp_cpx_data_ca_76_0_in[28]) );
  AO22X1_RVT U229 ( .A1(n228), .A2(add_frac_out[38]), .A3(n227), .A4(
        mul_frac_out[27]), .Y(n174) );
  AO22X1_RVT U230 ( .A1(n230), .A2(div_frac_out[27]), .A3(n229), .A4(
        add_frac_out[27]), .Y(n173) );
  OR2X1_RVT U231 ( .A1(n174), .A2(n173), .Y(fp_cpx_data_ca_76_0_in[27]) );
  AO22X1_RVT U232 ( .A1(n228), .A2(add_frac_out[37]), .A3(n227), .A4(
        mul_frac_out[26]), .Y(n176) );
  AO22X1_RVT U233 ( .A1(n230), .A2(div_frac_out[26]), .A3(n229), .A4(
        add_frac_out[26]), .Y(n175) );
  OR2X1_RVT U234 ( .A1(n176), .A2(n175), .Y(fp_cpx_data_ca_76_0_in[26]) );
  AO22X1_RVT U235 ( .A1(n228), .A2(add_frac_out[36]), .A3(n227), .A4(
        mul_frac_out[25]), .Y(n178) );
  AO22X1_RVT U236 ( .A1(n230), .A2(div_frac_out[25]), .A3(n229), .A4(
        add_frac_out[25]), .Y(n177) );
  OR2X1_RVT U237 ( .A1(n178), .A2(n177), .Y(fp_cpx_data_ca_76_0_in[25]) );
  AO22X1_RVT U238 ( .A1(n228), .A2(add_frac_out[35]), .A3(n227), .A4(
        mul_frac_out[24]), .Y(n180) );
  AO22X1_RVT U239 ( .A1(n230), .A2(div_frac_out[24]), .A3(n229), .A4(
        add_frac_out[24]), .Y(n179) );
  OR2X1_RVT U240 ( .A1(n180), .A2(n179), .Y(fp_cpx_data_ca_76_0_in[24]) );
  AO22X1_RVT U241 ( .A1(n228), .A2(add_frac_out[34]), .A3(n227), .A4(
        mul_frac_out[23]), .Y(n182) );
  AO22X1_RVT U242 ( .A1(n230), .A2(div_frac_out[23]), .A3(n229), .A4(
        add_frac_out[23]), .Y(n181) );
  OR2X1_RVT U243 ( .A1(n182), .A2(n181), .Y(fp_cpx_data_ca_76_0_in[23]) );
  AO22X1_RVT U244 ( .A1(n228), .A2(add_frac_out[33]), .A3(n227), .A4(
        mul_frac_out[22]), .Y(n184) );
  AO22X1_RVT U245 ( .A1(n230), .A2(div_frac_out[22]), .A3(n229), .A4(
        add_frac_out[22]), .Y(n183) );
  OR2X1_RVT U246 ( .A1(n184), .A2(n183), .Y(fp_cpx_data_ca_76_0_in[22]) );
  AO22X1_RVT U247 ( .A1(n228), .A2(add_frac_out[32]), .A3(n227), .A4(
        mul_frac_out[21]), .Y(n186) );
  AO22X1_RVT U248 ( .A1(n230), .A2(div_frac_out[21]), .A3(n229), .A4(
        add_frac_out[21]), .Y(n185) );
  OR2X1_RVT U249 ( .A1(n186), .A2(n185), .Y(fp_cpx_data_ca_76_0_in[21]) );
  AO22X1_RVT U250 ( .A1(n228), .A2(add_frac_out[31]), .A3(n227), .A4(
        mul_frac_out[20]), .Y(n188) );
  AO22X1_RVT U251 ( .A1(n230), .A2(div_frac_out[20]), .A3(n229), .A4(
        add_frac_out[20]), .Y(n187) );
  OR2X1_RVT U252 ( .A1(n188), .A2(n187), .Y(fp_cpx_data_ca_76_0_in[20]) );
  AO22X1_RVT U253 ( .A1(n228), .A2(add_frac_out[30]), .A3(n227), .A4(
        mul_frac_out[19]), .Y(n190) );
  AO22X1_RVT U254 ( .A1(n230), .A2(div_frac_out[19]), .A3(n229), .A4(
        add_frac_out[19]), .Y(n189) );
  OR2X1_RVT U255 ( .A1(n190), .A2(n189), .Y(fp_cpx_data_ca_76_0_in[19]) );
  AO22X1_RVT U256 ( .A1(n228), .A2(add_frac_out[29]), .A3(n227), .A4(
        mul_frac_out[18]), .Y(n192) );
  AO22X1_RVT U257 ( .A1(n230), .A2(div_frac_out[18]), .A3(n229), .A4(
        add_frac_out[18]), .Y(n191) );
  OR2X1_RVT U258 ( .A1(n192), .A2(n191), .Y(fp_cpx_data_ca_76_0_in[18]) );
  AO22X1_RVT U259 ( .A1(n228), .A2(add_frac_out[28]), .A3(n227), .A4(
        mul_frac_out[17]), .Y(n194) );
  AO22X1_RVT U260 ( .A1(n230), .A2(div_frac_out[17]), .A3(n229), .A4(
        add_frac_out[17]), .Y(n193) );
  OR2X1_RVT U261 ( .A1(n194), .A2(n193), .Y(fp_cpx_data_ca_76_0_in[17]) );
  AO22X1_RVT U262 ( .A1(n228), .A2(add_frac_out[27]), .A3(n227), .A4(
        mul_frac_out[16]), .Y(n196) );
  AO22X1_RVT U263 ( .A1(n230), .A2(div_frac_out[16]), .A3(n229), .A4(
        add_frac_out[16]), .Y(n195) );
  OR2X1_RVT U264 ( .A1(n196), .A2(n195), .Y(fp_cpx_data_ca_76_0_in[16]) );
  AO22X1_RVT U265 ( .A1(n228), .A2(add_frac_out[26]), .A3(n227), .A4(
        mul_frac_out[15]), .Y(n198) );
  AO22X1_RVT U266 ( .A1(n230), .A2(div_frac_out[15]), .A3(n229), .A4(
        add_frac_out[15]), .Y(n197) );
  OR2X1_RVT U267 ( .A1(n198), .A2(n197), .Y(fp_cpx_data_ca_76_0_in[15]) );
  AO22X1_RVT U268 ( .A1(n228), .A2(add_frac_out[25]), .A3(n227), .A4(
        mul_frac_out[14]), .Y(n200) );
  AO22X1_RVT U269 ( .A1(n230), .A2(div_frac_out[14]), .A3(n229), .A4(
        add_frac_out[14]), .Y(n199) );
  OR2X1_RVT U270 ( .A1(n200), .A2(n199), .Y(fp_cpx_data_ca_76_0_in[14]) );
  AO22X1_RVT U271 ( .A1(n228), .A2(add_frac_out[24]), .A3(n227), .A4(
        mul_frac_out[13]), .Y(n202) );
  AO22X1_RVT U272 ( .A1(n230), .A2(div_frac_out[13]), .A3(n229), .A4(
        add_frac_out[13]), .Y(n201) );
  OR2X1_RVT U273 ( .A1(n202), .A2(n201), .Y(fp_cpx_data_ca_76_0_in[13]) );
  AO22X1_RVT U274 ( .A1(n228), .A2(add_frac_out[23]), .A3(n227), .A4(
        mul_frac_out[12]), .Y(n204) );
  AO22X1_RVT U275 ( .A1(n230), .A2(div_frac_out[12]), .A3(n229), .A4(
        add_frac_out[12]), .Y(n203) );
  OR2X1_RVT U276 ( .A1(n204), .A2(n203), .Y(fp_cpx_data_ca_76_0_in[12]) );
  AO22X1_RVT U277 ( .A1(n228), .A2(add_frac_out[22]), .A3(n227), .A4(
        mul_frac_out[11]), .Y(n206) );
  AO22X1_RVT U278 ( .A1(n230), .A2(div_frac_out[11]), .A3(n229), .A4(
        add_frac_out[11]), .Y(n205) );
  OR2X1_RVT U279 ( .A1(n206), .A2(n205), .Y(fp_cpx_data_ca_76_0_in[11]) );
  AO22X1_RVT U280 ( .A1(n228), .A2(add_frac_out[21]), .A3(n227), .A4(
        mul_frac_out[10]), .Y(n208) );
  AO22X1_RVT U281 ( .A1(n230), .A2(div_frac_out[10]), .A3(n229), .A4(
        add_frac_out[10]), .Y(n207) );
  OR2X1_RVT U282 ( .A1(n208), .A2(n207), .Y(fp_cpx_data_ca_76_0_in[10]) );
  AO22X1_RVT U283 ( .A1(n228), .A2(add_frac_out[20]), .A3(n227), .A4(
        mul_frac_out[9]), .Y(n210) );
  AO22X1_RVT U284 ( .A1(n230), .A2(div_frac_out[9]), .A3(n229), .A4(
        add_frac_out[9]), .Y(n209) );
  OR2X1_RVT U285 ( .A1(n210), .A2(n209), .Y(fp_cpx_data_ca_76_0_in[9]) );
  AO22X1_RVT U286 ( .A1(n228), .A2(add_frac_out[19]), .A3(n227), .A4(
        mul_frac_out[8]), .Y(n212) );
  AO22X1_RVT U287 ( .A1(n230), .A2(div_frac_out[8]), .A3(n229), .A4(
        add_frac_out[8]), .Y(n211) );
  OR2X1_RVT U288 ( .A1(n212), .A2(n211), .Y(fp_cpx_data_ca_76_0_in[8]) );
  AO22X1_RVT U289 ( .A1(n228), .A2(add_frac_out[18]), .A3(n227), .A4(
        mul_frac_out[7]), .Y(n214) );
  AO22X1_RVT U290 ( .A1(n230), .A2(div_frac_out[7]), .A3(n229), .A4(
        add_frac_out[7]), .Y(n213) );
  OR2X1_RVT U291 ( .A1(n214), .A2(n213), .Y(fp_cpx_data_ca_76_0_in[7]) );
  AO22X1_RVT U292 ( .A1(n228), .A2(add_frac_out[17]), .A3(n227), .A4(
        mul_frac_out[6]), .Y(n216) );
  AO22X1_RVT U293 ( .A1(n230), .A2(div_frac_out[6]), .A3(n229), .A4(
        add_frac_out[6]), .Y(n215) );
  OR2X1_RVT U294 ( .A1(n216), .A2(n215), .Y(fp_cpx_data_ca_76_0_in[6]) );
  AO22X1_RVT U295 ( .A1(n228), .A2(add_frac_out[16]), .A3(n227), .A4(
        mul_frac_out[5]), .Y(n218) );
  AO22X1_RVT U296 ( .A1(n230), .A2(div_frac_out[5]), .A3(n229), .A4(
        add_frac_out[5]), .Y(n217) );
  OR2X1_RVT U297 ( .A1(n218), .A2(n217), .Y(fp_cpx_data_ca_76_0_in[5]) );
  AO22X1_RVT U298 ( .A1(n228), .A2(add_frac_out[15]), .A3(n227), .A4(
        mul_frac_out[4]), .Y(n220) );
  AO22X1_RVT U299 ( .A1(n230), .A2(div_frac_out[4]), .A3(n229), .A4(
        add_frac_out[4]), .Y(n219) );
  OR2X1_RVT U300 ( .A1(n220), .A2(n219), .Y(fp_cpx_data_ca_76_0_in[4]) );
  AO22X1_RVT U301 ( .A1(n228), .A2(add_frac_out[14]), .A3(n227), .A4(
        mul_frac_out[3]), .Y(n222) );
  AO22X1_RVT U302 ( .A1(n230), .A2(div_frac_out[3]), .A3(n229), .A4(
        add_frac_out[3]), .Y(n221) );
  OR2X1_RVT U303 ( .A1(n222), .A2(n221), .Y(fp_cpx_data_ca_76_0_in[3]) );
  AO22X1_RVT U304 ( .A1(n228), .A2(add_frac_out[13]), .A3(n227), .A4(
        mul_frac_out[2]), .Y(n224) );
  AO22X1_RVT U305 ( .A1(n230), .A2(div_frac_out[2]), .A3(n229), .A4(
        add_frac_out[2]), .Y(n223) );
  OR2X1_RVT U306 ( .A1(n224), .A2(n223), .Y(fp_cpx_data_ca_76_0_in[2]) );
  AO22X1_RVT U307 ( .A1(n228), .A2(add_frac_out[12]), .A3(n227), .A4(
        mul_frac_out[1]), .Y(n226) );
  AO22X1_RVT U308 ( .A1(n230), .A2(div_frac_out[1]), .A3(n229), .A4(
        add_frac_out[1]), .Y(n225) );
  OR2X1_RVT U309 ( .A1(n226), .A2(n225), .Y(fp_cpx_data_ca_76_0_in[1]) );
  AO22X1_RVT U310 ( .A1(n228), .A2(add_frac_out[11]), .A3(n227), .A4(
        mul_frac_out[0]), .Y(n232) );
  AO22X1_RVT U311 ( .A1(n230), .A2(div_frac_out[0]), .A3(n229), .A4(
        add_frac_out[0]), .Y(n231) );
  OR2X1_RVT U312 ( .A1(n232), .A2(n231), .Y(fp_cpx_data_ca_76_0_in[0]) );
endmodule


module fpu_out ( d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, div_id_out_in, 
        m6stg_id_in, add_id_out_in, div_exc_out, d8stg_fdivd, d8stg_fdivs, 
        div_sign_out, div_exp_out, div_frac_out, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, add_exc_out, a6stg_fcmpop, add_cc_out, add_fcc_out, 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        add_sign_out, add_exp_out, add_frac_out, arst_l, grst_l, rclk, 
        fp_cpx_req_cq, fp_cpx_data_ca, se, si, so, add_dest_rdy_BAR, 
        div_dest_rdy_BAR, mul_dest_rdy_BAR );
  input [9:0] div_id_out_in;
  input [9:0] m6stg_id_in;
  input [9:0] add_id_out_in;
  input [4:0] div_exc_out;
  input [10:0] div_exp_out;
  input [51:0] div_frac_out;
  input [4:0] mul_exc_out;
  input [10:0] mul_exp_out;
  input [51:0] mul_frac_out;
  input [4:0] add_exc_out;
  input [1:0] add_cc_out;
  input [1:0] add_fcc_out;
  input [10:0] add_exp_out;
  input [63:0] add_frac_out;
  output [7:0] fp_cpx_req_cq;
  output [144:0] fp_cpx_data_ca;
  input d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out,
         a6stg_fcmpop, a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst,
         a6stg_int_dst, add_sign_out, arst_l, grst_l, rclk, se, si;
  output so, add_dest_rdy_BAR, div_dest_rdy_BAR, mul_dest_rdy_BAR;
  wire   add_dest_rdy, mul_dest_rdy, div_dest_rdy, net211144, net211145,
         net211146, net211147;
  wire   [1:0] req_thread;
  wire   [2:0] dest_rdy;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66;
  assign add_dest_rdy_BAR = add_dest_rdy;
  assign mul_dest_rdy_BAR = mul_dest_rdy;
  assign div_dest_rdy_BAR = div_dest_rdy;

  fpu_out_ctl fpu_out_ctl ( .d8stg_fdiv_in(d8stg_fdiv_in), .m6stg_fmul_in(
        m6stg_fmul_in), .a6stg_fadd_in(a6stg_fadd_in), .div_id_out_in(
        div_id_out_in), .m6stg_id_in(m6stg_id_in), .add_id_out_in(
        add_id_out_in), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), 
        .fp_cpx_req_cq(fp_cpx_req_cq), .req_thread(req_thread), .dest_rdy(
        dest_rdy), .se(se), .si(net211147), .add_dest_rdy_BAR(add_dest_rdy), 
        .div_dest_rdy_BAR(div_dest_rdy), .mul_dest_rdy_BAR(mul_dest_rdy) );
  fpu_out_dp fpu_out_dp ( .dest_rdy(dest_rdy), .req_thread(req_thread), 
        .div_exc_out(div_exc_out), .d8stg_fdivd(d8stg_fdivd), .d8stg_fdivs(
        d8stg_fdivs), .div_sign_out(div_sign_out), .div_exp_out(div_exp_out), 
        .div_frac_out(div_frac_out), .mul_exc_out({mul_exc_out[4:2], net211144, 
        mul_exc_out[0]}), .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), 
        .m6stg_fmuls(m6stg_fmuls), .mul_sign_out(mul_sign_out), .mul_exp_out(
        mul_exp_out), .mul_frac_out(mul_frac_out), .add_exc_out({
        add_exc_out[4:2], net211145, add_exc_out[0]}), .a6stg_fcmpop(
        a6stg_fcmpop), .add_cc_out(add_cc_out), .add_fcc_out(add_fcc_out), 
        .a6stg_dbl_dst(a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), 
        .a6stg_long_dst(a6stg_long_dst), .a6stg_int_dst(a6stg_int_dst), 
        .add_sign_out(add_sign_out), .add_exp_out(add_exp_out), .add_frac_out(
        add_frac_out), .rclk(rclk), .fp_cpx_data_ca({fp_cpx_data_ca[144:143], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, fp_cpx_data_ca[135:134], 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, fp_cpx_data_ca[76:72], 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        fp_cpx_data_ca[69:65], SYNOPSYS_UNCONNECTED__66, fp_cpx_data_ca[63:0]}), .se(se), .si(net211146) );
endmodule


module test_stub_scan ( mux_drive_disable, mem_write_disable, sehold, se, 
        testmode_l, mem_bypass, so_0, so_1, so_2, ctu_tst_pre_grst_l, arst_l, 
        global_shift_enable, ctu_tst_scan_disable, ctu_tst_scanmode, 
        ctu_tst_macrotest, ctu_tst_short_chain, long_chain_so_0, 
        short_chain_so_0, long_chain_so_1, short_chain_so_1, long_chain_so_2, 
        short_chain_so_2 );
  input ctu_tst_pre_grst_l, arst_l, global_shift_enable, ctu_tst_scan_disable,
         ctu_tst_scanmode, ctu_tst_macrotest, ctu_tst_short_chain,
         long_chain_so_0, short_chain_so_0, long_chain_so_1, short_chain_so_1,
         long_chain_so_2, short_chain_so_2;
  output mux_drive_disable, mem_write_disable, sehold, se, testmode_l,
         mem_bypass, so_0, so_1, so_2;
  wire   global_shift_enable, n1, n2;
  assign se = global_shift_enable;

  NAND2X0_RVT U1 ( .A1(ctu_tst_scanmode), .A2(ctu_tst_short_chain), .Y(n1) );
  OA221X1_RVT U2 ( .A1(n1), .A2(ctu_tst_scan_disable), .A3(n1), .A4(
        global_shift_enable), .A5(long_chain_so_0), .Y(so_0) );
  INVX1_RVT U3 ( .A(global_shift_enable), .Y(n2) );
  NAND2X0_RVT U4 ( .A1(ctu_tst_pre_grst_l), .A2(n2), .Y(mem_write_disable) );
  AND2X1_RVT U5 ( .A1(ctu_tst_macrotest), .A2(n2), .Y(sehold) );
endmodule


module bw_u1_scanl_2x_0 ( so, ck, sd_BAR );
  input ck, sd_BAR;
  output so;
  wire   sd, n3;
  assign sd = sd_BAR;

  LATCHX1_RVT so_l_reg ( .CLK(n3), .D(sd), .QN(so) );
  INVX0_RVT U4 ( .A(ck), .Y(n3) );
endmodule


module zsoffasr_prim_0 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   N10, n1;

  DFFASRX1_RVT q_reg ( .D(N10), .CLK(ck), .RSTB(r_l), .SETB(1'b1), .Q(q) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  AND3X1_RVT U4 ( .A1(r_l), .A2(d), .A3(n1), .Y(N10) );
  OR2X1_RVT U6 ( .A1(q), .A2(n1), .Y(so) );
endmodule


module bw_u1_soffasr_2x_0 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   net210538, net210539;

  zsoffasr_prim_0 i0 ( .q(q), .so(so), .ck(ck), .d(d), .r_l(r_l), .s_l(
        net210538), .se(se), .sd(net210539) );
endmodule


module bw_u1_scanl_2x_2 ( so, sd, ck );
  input sd, ck;
  output so;
  wire   n4, n5;

  LATCHX1_RVT so_l_reg ( .CLK(n4), .D(n5), .QN(so) );
  INVX0_RVT U4 ( .A(ck), .Y(n4) );
  INVX1_RVT U3 ( .A(sd), .Y(n5) );
endmodule


module zsoffasr_prim_3 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   N10, n1;

  DFFARX1_RVT q_reg ( .D(N10), .CLK(ck), .RSTB(r_l), .Q(q) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OA221X1_RVT U4 ( .A1(se), .A2(d), .A3(n1), .A4(sd), .A5(r_l), .Y(N10) );
  OR2X1_RVT U5 ( .A1(q), .A2(n1), .Y(so) );
endmodule


module bw_u1_soffasr_2x_3 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   net210264;

  zsoffasr_prim_3 i0 ( .q(q), .so(so), .ck(ck), .d(d), .r_l(r_l), .s_l(
        net210264), .se(se), .sd(sd) );
endmodule


module synchronizer_asr_0 ( sync_out, so, async_in, gclk, rclk, arst_l, si, se
 );
  input async_in, gclk, rclk, arst_l, si, se;
  output sync_out, so;
  wire   pre_sync_out, so_rptr, so_lockup, net210785;

  bw_u1_soffasr_2x_0 repeater ( .q(pre_sync_out), .so(so_rptr), .ck(gclk), .d(
        async_in), .r_l(arst_l), .s_l(1'b1), .se(se), .sd(net210785) );
  bw_u1_scanl_2x_2 lockup ( .so(so_lockup), .sd(so_rptr), .ck(gclk) );
  bw_u1_soffasr_2x_3 syncff ( .q(sync_out), .so(so), .ck(rclk), .d(
        pre_sync_out), .r_l(arst_l), .s_l(1'b1), .se(se), .sd(so_lockup) );
endmodule


module bw_u1_scanl_2x_1 ( so, sd, ck );
  input sd, ck;
  output so;
  wire   n4, n5;

  LATCHX1_RVT so_l_reg ( .CLK(n4), .D(n5), .QN(so) );
  INVX0_RVT U4 ( .A(ck), .Y(n4) );
  INVX1_RVT U3 ( .A(sd), .Y(n5) );
endmodule


module zsoffasr_prim_1 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   N10, n1;

  DFFASRX1_RVT q_reg ( .D(N10), .CLK(ck), .RSTB(1'b1), .SETB(1'b1), .Q(q) );
  INVX1_RVT U4 ( .A(se), .Y(n1) );
  OR2X1_RVT U5 ( .A1(q), .A2(n1), .Y(so) );
  AO22X1_RVT U6 ( .A1(se), .A2(sd), .A3(n1), .A4(d), .Y(N10) );
endmodule


module bw_u1_soffasr_2x_1 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   net210268, net210269;

  zsoffasr_prim_1 i0 ( .so(so), .ck(ck), .d(d), .r_l(net210268), .s_l(
        net210269), .se(se), .sd(sd) );
endmodule


module zsoffasr_prim_2 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   N10, n1;

  DFFX1_RVT q_reg ( .D(N10), .CLK(ck), .Q(q) );
  INVX1_RVT U3 ( .A(se), .Y(n1) );
  OR2X1_RVT U4 ( .A1(sd), .A2(n1), .Y(N10) );
  OR2X1_RVT U5 ( .A1(q), .A2(n1), .Y(so) );
endmodule


module bw_u1_soffasr_2x_2 ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   net210265, net210266, net210267;

  zsoffasr_prim_2 i0 ( .q(q), .so(so), .ck(ck), .d(net210265), .r_l(net210266), 
        .s_l(net210267), .se(se), .sd(sd) );
endmodule


module synchronizer_asr_1 ( sync_out, so, async_in, gclk, rclk, arst_l, si, se
 );
  input async_in, gclk, rclk, arst_l, si, se;
  output sync_out, so;
  wire   pre_sync_out, so_rptr, so_lockup, net210270, net210271, net210272;

  bw_u1_soffasr_2x_2 repeater ( .q(pre_sync_out), .so(so_rptr), .ck(gclk), .d(
        net210271), .r_l(net210272), .s_l(1'b1), .se(se), .sd(si) );
  bw_u1_scanl_2x_1 lockup ( .so(so_lockup), .sd(so_rptr), .ck(gclk) );
  bw_u1_soffasr_2x_1 syncff ( .so(so), .ck(rclk), .d(pre_sync_out), .r_l(
        net210270), .s_l(1'b1), .se(se), .sd(so_lockup) );
endmodule


module bw_u1_syncff_4x ( so, ck, d, se, sd, q_BAR );
  input ck, d, se, sd;
  output so, q_BAR;
  wire   N3;
  assign N3 = d;

  DFFX1_RVT q_r_reg ( .D(N3), .CLK(ck), .QN(q_BAR) );
endmodule


module cluster_header ( dbginit_l, cluster_grst_l, rclk, so, gclk, 
        cluster_cken, arst_l, grst_l, adbginit_l, gdbginit_l, si, se );
  input gclk, cluster_cken, arst_l, grst_l, adbginit_l, gdbginit_l, si, se;
  output dbginit_l, cluster_grst_l, rclk, so;
  wire   pre_sync_enable, sync_enable, rst_sync_so, net210932, net210933,
         net210934;

  bw_u1_syncff_4x sync_cluster_master ( .ck(gclk), .d(cluster_cken), .se(1'b0), 
        .sd(1'b0), .q_BAR(pre_sync_enable) );
  bw_u1_scanl_2x_0 sync_cluster_slave ( .so(sync_enable), .ck(gclk), .sd_BAR(
        pre_sync_enable) );
  synchronizer_asr_0 rst_repeater ( .sync_out(cluster_grst_l), .so(rst_sync_so), .async_in(grst_l), .gclk(gclk), .rclk(rclk), .arst_l(arst_l), .si(net210934), 
        .se(se) );
  synchronizer_asr_1 dbginit_repeater ( .so(so), .async_in(net210932), .gclk(
        gclk), .rclk(rclk), .arst_l(net210933), .si(rst_sync_so), .se(se) );
  AND2X1_RVT U3 ( .A1(sync_enable), .A2(gclk), .Y(rclk) );
endmodule


module bw_clk_cl_fpu_cmp ( so, dbginit_l, cluster_grst_l, rclk, si, se, 
        adbginit_l, gdbginit_l, arst_l, grst_l, cluster_cken, gclk );
  input si, se, adbginit_l, gdbginit_l, arst_l, grst_l, cluster_cken, gclk;
  output so, dbginit_l, cluster_grst_l, rclk;
  wire   net211141, net211142, net211143;

  cluster_header I0 ( .cluster_grst_l(cluster_grst_l), .rclk(rclk), .so(so), 
        .gclk(gclk), .cluster_cken(cluster_cken), .arst_l(arst_l), .grst_l(
        grst_l), .adbginit_l(net211141), .gdbginit_l(net211142), .si(net211143), .se(se) );
endmodule


module fpu_bufrpt_grp32_0 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp64_0 ( in, out );
  input [63:0] in;
  output [63:0] out;

  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[55];
  assign out[54] = in[54];
  assign out[53] = in[53];
  assign out[52] = in[52];
  assign out[51] = in[51];
  assign out[50] = in[50];
  assign out[49] = in[49];
  assign out[48] = in[48];
  assign out[47] = in[47];
  assign out[46] = in[46];
  assign out[45] = in[45];
  assign out[44] = in[44];
  assign out[43] = in[43];
  assign out[42] = in[42];
  assign out[41] = in[41];
  assign out[40] = in[40];
  assign out[39] = in[39];
  assign out[38] = in[38];
  assign out[37] = in[37];
  assign out[36] = in[36];
  assign out[35] = in[35];
  assign out[34] = in[34];
  assign out[33] = in[33];
  assign out[32] = in[32];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp4_0 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_0 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_0 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[11] = in[11];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_inq ( in, out );
  input [155:0] in;
  output [155:0] out;

  assign out[155] = in[155];
  assign out[154] = in[154];
  assign out[153] = in[153];
  assign out[152] = in[152];
  assign out[151] = in[151];
  assign out[150] = in[150];
  assign out[149] = in[149];
  assign out[148] = in[148];
  assign out[147] = in[147];
  assign out[146] = in[146];
  assign out[145] = in[145];
  assign out[144] = in[144];
  assign out[143] = in[143];
  assign out[142] = in[142];
  assign out[141] = in[141];
  assign out[140] = in[140];
  assign out[139] = in[139];
  assign out[138] = in[138];
  assign out[137] = in[137];
  assign out[136] = in[136];
  assign out[135] = in[135];
  assign out[134] = in[134];
  assign out[133] = in[133];
  assign out[132] = in[132];
  assign out[131] = in[131];
  assign out[130] = in[130];
  assign out[129] = in[129];
  assign out[128] = in[128];
  assign out[127] = in[127];
  assign out[126] = in[126];
  assign out[125] = in[125];
  assign out[124] = in[124];
  assign out[123] = in[123];
  assign out[122] = in[122];
  assign out[121] = in[121];
  assign out[120] = in[120];
  assign out[119] = in[119];
  assign out[118] = in[118];
  assign out[117] = in[117];
  assign out[116] = in[116];
  assign out[115] = in[115];
  assign out[114] = in[114];
  assign out[113] = in[113];
  assign out[112] = in[112];
  assign out[111] = in[111];
  assign out[110] = in[110];
  assign out[109] = in[109];
  assign out[108] = in[108];
  assign out[107] = in[107];
  assign out[106] = in[106];
  assign out[105] = in[105];
  assign out[104] = in[104];
  assign out[103] = in[103];
  assign out[102] = in[102];
  assign out[101] = in[101];
  assign out[100] = in[100];
  assign out[99] = in[99];
  assign out[98] = in[98];
  assign out[97] = in[97];
  assign out[96] = in[96];
  assign out[95] = in[95];
  assign out[94] = in[94];
  assign out[93] = in[93];
  assign out[92] = in[92];
  assign out[91] = in[91];
  assign out[90] = in[90];
  assign out[89] = in[89];
  assign out[88] = in[88];
  assign out[87] = in[87];
  assign out[86] = in[86];
  assign out[85] = in[85];
  assign out[84] = in[84];
  assign out[83] = in[83];
  assign out[82] = in[82];
  assign out[81] = in[81];
  assign out[80] = in[80];
  assign out[79] = in[79];
  assign out[78] = in[78];
  assign out[77] = in[77];
  assign out[76] = in[76];
  assign out[75] = in[75];
  assign out[74] = in[74];
  assign out[73] = in[73];
  assign out[72] = in[72];
  assign out[71] = in[71];
  assign out[70] = in[70];
  assign out[69] = in[69];
  assign out[68] = in[68];
  assign out[67] = in[67];
  assign out[66] = in[66];
  assign out[65] = in[65];
  assign out[64] = in[64];
  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[55];
  assign out[54] = in[54];
  assign out[53] = in[53];
  assign out[52] = in[52];
  assign out[51] = in[51];
  assign out[50] = in[50];
  assign out[49] = in[49];
  assign out[48] = in[48];
  assign out[47] = in[47];
  assign out[46] = in[46];
  assign out[45] = in[45];
  assign out[44] = in[44];
  assign out[43] = in[43];
  assign out[42] = in[42];
  assign out[41] = in[41];
  assign out[40] = in[40];
  assign out[39] = in[39];
  assign out[38] = in[38];
  assign out[37] = in[37];
  assign out[36] = in[36];
  assign out[35] = in[35];
  assign out[34] = in[34];
  assign out[33] = in[33];
  assign out[32] = in[32];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];

endmodule


module fpu_bufrpt_grp64_1 ( in, out );
  input [63:0] in;
  output [63:0] out;

  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[55];
  assign out[54] = in[54];
  assign out[53] = in[53];
  assign out[52] = in[52];
  assign out[51] = in[51];
  assign out[50] = in[50];
  assign out[49] = in[49];
  assign out[48] = in[48];
  assign out[47] = in[47];
  assign out[46] = in[46];
  assign out[45] = in[45];
  assign out[44] = in[44];
  assign out[43] = in[43];
  assign out[42] = in[42];
  assign out[41] = in[41];
  assign out[40] = in[40];
  assign out[39] = in[39];
  assign out[38] = in[38];
  assign out[37] = in[37];
  assign out[36] = in[36];
  assign out[35] = in[35];
  assign out[34] = in[34];
  assign out[33] = in[33];
  assign out[32] = in[32];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_1 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[9] = in[9];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];

endmodule


module fpu_rptr_fp_cpx_grp16_3 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[3] = in[3];

endmodule


module fpu_rptr_fp_cpx_grp16_5 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[5] = in[5];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_6 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_7 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_8 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16_9 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_1 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_2 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_3 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_4 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_5 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16_6 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];

endmodule


module fpu_bufrpt_grp32_1 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_2 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_3 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_4 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_5 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_6 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_7 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_8 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_9 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp32_10 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp4_2 ( in, out );
  input [3:0] in;
  output [3:0] out;
  wire   \in[3] ;
  assign out[3] = \in[3] ;
  assign \in[3]  = in[3];

endmodule


module fpu_bufrpt_grp4_3 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];

endmodule


module fpu_bufrpt_grp4_4 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp4_5 ( in, out );
  input [3:0] in;
  output [3:0] out;
  wire   \in[3] ;
  assign out[3] = \in[3] ;
  assign \in[3]  = in[3];

endmodule


module fpu_bufrpt_grp4_6 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];

endmodule


module fpu_bufrpt_grp4_7 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];

endmodule


module fpu_bufrpt_grp4_8 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];

endmodule


module fpu_bufrpt_grp4_9 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];

endmodule


module fpu_bufrpt_grp4_10 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];

endmodule


module fpu_rptr_groups ( inq_in1, inq_in2, inq_id, inq_op, inq_rnd_mode, 
        inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0, 
        inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, 
        inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l, 
        ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain, 
        global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l, 
        fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf, 
        pcx_fpio_data_px2, pcx_fpio_data_rdy_px2, fp_cpx_req_cq, 
        fp_cpx_data_ca, inq_sram_din_unbuf, inq_in1_add_buf1, inq_in1_mul_buf1, 
        inq_in1_div_buf1, inq_in2_add_buf1, inq_in2_mul_buf1, inq_in2_div_buf1, 
        inq_id_add_buf1, inq_id_mul_buf1, inq_id_div_buf1, inq_op_add_buf1, 
        inq_op_div_buf1, inq_op_mul_buf1, inq_rnd_mode_add_buf1, 
        inq_rnd_mode_div_buf1, inq_rnd_mode_mul_buf1, 
        inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1, 
        inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1, 
        inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1, 
        inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1, 
        inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1, 
        inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1, 
        inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1, 
        inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1, 
        inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1, 
        inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1, 
        inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1, 
        inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1, 
        inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1, 
        inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1, 
        inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1, 
        ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1, 
        ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1, 
        ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1, 
        cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2, 
        se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4, 
        se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2, 
        arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3, 
        arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2, 
        fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1, 
        fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so, 
        pcx_fpio_data_px2_buf1, pcx_fpio_data_rdy_px2_buf1, fp_cpx_req_cq_buf1, 
        fp_cpx_data_ca_buf1, inq_sram_din_buf1 );
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  input [4:0] inq_id;
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [123:0] pcx_fpio_data_px2;
  input [7:0] fp_cpx_req_cq;
  input [144:0] fp_cpx_data_ca;
  input [155:0] inq_sram_din_unbuf;
  output [63:0] inq_in1_add_buf1;
  output [63:0] inq_in1_mul_buf1;
  output [63:0] inq_in1_div_buf1;
  output [63:0] inq_in2_add_buf1;
  output [63:0] inq_in2_mul_buf1;
  output [63:0] inq_in2_div_buf1;
  output [4:0] inq_id_add_buf1;
  output [4:0] inq_id_mul_buf1;
  output [4:0] inq_id_div_buf1;
  output [7:0] inq_op_add_buf1;
  output [7:0] inq_op_div_buf1;
  output [7:0] inq_op_mul_buf1;
  output [1:0] inq_rnd_mode_add_buf1;
  output [1:0] inq_rnd_mode_div_buf1;
  output [1:0] inq_rnd_mode_mul_buf1;
  output [123:0] pcx_fpio_data_px2_buf1;
  output [7:0] fp_cpx_req_cq_buf1;
  output [144:0] fp_cpx_data_ca_buf1;
  output [155:0] inq_sram_din_buf1;
  input inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0,
         inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l,
         ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain,
         global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l,
         fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf,
         pcx_fpio_data_rdy_px2;
  output inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1,
         inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1,
         inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1,
         inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1,
         inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1,
         inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1,
         inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1,
         inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1,
         inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1,
         inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1,
         inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1,
         inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1,
         inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1,
         inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1,
         inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1,
         ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1,
         ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1,
         ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1,
         cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2,
         se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4,
         se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2,
         arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3,
         arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2,
         fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1,
         fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so,
         pcx_fpio_data_rdy_px2_buf1;
  wire   se_add_buf1, se_mul64_buf1, so_buf1, arst_l_buf1, net211105,
         net211106, net211107, net211108, net211109, net211110, net211111,
         net211112, net211113, net211114, net211115, net211116, net211117,
         net211118, net211119, net211120, net211121, net211122, net211123,
         net211124, net211125, net211126, net211127, net211128, net211129,
         net211130, net211131, net211132, net211133, net211134, net211135,
         net211136, net211137, net211138, net211139, net211140;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97;

  fpu_bufrpt_grp32_0 i_inq_in1_add_buf1_hi ( .in(inq_in1[63:32]), .out(
        inq_in1_add_buf1[63:32]) );
  fpu_bufrpt_grp32_10 i_inq_in1_add_buf1_lo ( .in(inq_in1[31:0]), .out(
        inq_in1_add_buf1[31:0]) );
  fpu_bufrpt_grp32_9 i_inq_in1_mul_buf1_hi ( .in(inq_in1[63:32]), .out(
        inq_in1_mul_buf1[63:32]) );
  fpu_bufrpt_grp32_8 i_inq_in1_mul_buf1_lo ( .in(inq_in1[31:0]), .out(
        inq_in1_mul_buf1[31:0]) );
  fpu_bufrpt_grp64_0 i_inq_in1_div_buf1 ( .in(inq_in1), .out(inq_in1_div_buf1)
         );
  fpu_bufrpt_grp32_7 i_inq_in2_add_buf1_hi ( .in(inq_in2[63:32]), .out(
        inq_in2_add_buf1[63:32]) );
  fpu_bufrpt_grp32_6 i_inq_in2_add_buf1_lo ( .in(inq_in2[31:0]), .out(
        inq_in2_add_buf1[31:0]) );
  fpu_bufrpt_grp32_5 i_inq_in2_mul_buf1_hi ( .in(inq_in2[63:32]), .out(
        inq_in2_mul_buf1[63:32]) );
  fpu_bufrpt_grp32_4 i_inq_in2_mul_buf1_lo ( .in(inq_in2[31:0]), .out(
        inq_in2_mul_buf1[31:0]) );
  fpu_bufrpt_grp64_1 i_inq_in2_div_buf1 ( .in(inq_in2), .out(inq_in2_div_buf1)
         );
  fpu_bufrpt_grp32_3 i_inq_id_add_buf1 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 
        se_out_buf2, arst_l_out_buf3, fpu_grst_l_in_buf2, inq_id, inq_op, 
        inq_rnd_mode, inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, 
        inq_in2_50_0_neq_0, inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs}), .out({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, se_in_buf3, arst_l_add_buf4, 
        fpu_grst_l_add_buf3, inq_id_add_buf1, inq_op_add_buf1, 
        inq_rnd_mode_add_buf1, inq_in1_50_0_neq_0_add_buf1, 
        SYNOPSYS_UNCONNECTED__4, inq_in1_53_32_neq_0_add_buf1, 
        inq_in1_exp_eq_0_add_buf1, inq_in1_exp_neq_ffs_add_buf1, 
        inq_in2_50_0_neq_0_add_buf1, SYNOPSYS_UNCONNECTED__5, 
        inq_in2_53_32_neq_0_add_buf1, inq_in2_exp_eq_0_add_buf1, 
        inq_in2_exp_neq_ffs_add_buf1}) );
  fpu_bufrpt_grp32_2 i_inq_id_mul_buf1 ( .in({1'b0, 1'b0, 1'b0, se_in_buf3, 
        arst_l_mul_buf2, fpu_grst_l_mul_buf1, fmul_clken_l, inq_id, inq_op, 
        inq_rnd_mode, inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, 
        inq_in2_50_0_neq_0, inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs}), .out({SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, se_mul_buf4, 
        arst_l_out_buf3, fpu_grst_l_in_buf2, fmul_clken_l_buf1, 
        inq_id_mul_buf1, inq_op_mul_buf1, inq_rnd_mode_mul_buf1, 
        inq_in1_50_0_neq_0_mul_buf1, SYNOPSYS_UNCONNECTED__9, 
        inq_in1_53_32_neq_0_mul_buf1, inq_in1_exp_eq_0_mul_buf1, 
        inq_in1_exp_neq_ffs_mul_buf1, inq_in2_50_0_neq_0_mul_buf1, 
        SYNOPSYS_UNCONNECTED__10, inq_in2_53_32_neq_0_mul_buf1, 
        inq_in2_exp_eq_0_mul_buf1, inq_in2_exp_neq_ffs_mul_buf1}) );
  fpu_bufrpt_grp32_1 i_inq_id_div_buf1 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        se_mul_buf4, arst_l_mul_buf2, inq_id, inq_op, inq_rnd_mode, 
        inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0, 
        inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, 
        inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs}), .out({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, se_div_buf5, 
        arst_l_in_buf3, inq_id_div_buf1, inq_op_div_buf1, 
        inq_rnd_mode_div_buf1, inq_in1_50_0_neq_0_div_buf1, 
        inq_in1_53_0_neq_0_div_buf1, inq_in1_53_32_neq_0_div_buf1, 
        inq_in1_exp_eq_0_div_buf1, inq_in1_exp_neq_ffs_div_buf1, 
        inq_in2_50_0_neq_0_div_buf1, inq_in2_53_0_neq_0_div_buf1, 
        inq_in2_53_32_neq_0_div_buf1, inq_in2_exp_eq_0_div_buf1, 
        inq_in2_exp_neq_ffs_div_buf1}) );
  fpu_bufrpt_grp4_0 i_ctu_tst_buf1_hi ( .in({ctu_tst_short_chain, 
        ctu_tst_macrotest, ctu_tst_scan_disable, ctu_tst_pre_grst_l}), .out({
        ctu_tst_short_chain_buf1, ctu_tst_macrotest_buf1, 
        ctu_tst_scan_disable_buf1, ctu_tst_pre_grst_l_buf1}) );
  fpu_bufrpt_grp4_10 i_ctu_tst_buf1_lo ( .in({ctu_tst_scanmode, 
        global_shift_enable, 1'b0, 1'b0}), .out({ctu_tst_scanmode_buf1, 
        global_shift_enable_buf1, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17}) );
  fpu_bufrpt_grp4_9 i_cluster_cken_buf1 ( .in({cluster_cken, grst_l, 1'b0, 
        1'b0}), .out({cluster_cken_buf1, grst_l_buf1, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19}) );
  fpu_bufrpt_grp4_8 i_se_buf1 ( .in({se, se, so_unbuf, 1'b0}), .out({
        se_add_buf1, se_mul64_buf1, so_buf1, SYNOPSYS_UNCONNECTED__20}) );
  fpu_bufrpt_grp4_7 i_se_add_buf2 ( .in({se_add_buf1, se_add_buf1, se_add_buf1, 
        1'b0}), .out({se_add_exp_buf2, se_add_frac_buf2, se_out_buf2, 
        SYNOPSYS_UNCONNECTED__21}) );
  fpu_bufrpt_grp4_6 i_se_mul64_buf2 ( .in({se_mul64_buf1, se_mul64_buf1, 1'b0, 
        1'b0}), .out({se_mul64_buf2, se_cluster_header_buf2, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  fpu_bufrpt_grp4_5 i_arst_l_buf1 ( .in({arst_l, 1'b0, 1'b0, 1'b0}), .out({
        arst_l_buf1, SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26}) );
  fpu_bufrpt_grp4_4 i_arst_l_buf2 ( .in({arst_l_buf1, arst_l_buf1, arst_l_buf1, 
        fpu_grst_l}), .out({arst_l_mul_buf2, arst_l_cluster_header_buf2, 
        arst_l_div_buf2, fpu_grst_l_mul_buf1}) );
  fpu_bufrpt_grp4_3 i_fdiv_clken_l_buf1 ( .in({fdiv_clken_l, fdiv_clken_l, 
        1'b0, 1'b0}), .out({fdiv_clken_l_div_exp_buf1, 
        fdiv_clken_l_div_frac_buf1, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28}) );
  fpu_bufrpt_grp4_2 i_so_cluster_header_buf1 ( .in({scan_manual_6, 1'b0, 1'b0, 
        1'b0}), .out({scan_manual_6_buf1, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31}) );
  fpu_rptr_pcx_fpio_grp16_0 i_pcx_fpio_buf1_0 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 
        pcx_fpio_data_px2[112], pcx_fpio_data_px2[113], pcx_fpio_data_px2[114], 
        pcx_fpio_data_px2[115], pcx_fpio_data_px2[116], 1'b0, 
        pcx_fpio_data_px2[118], pcx_fpio_data_px2[119], pcx_fpio_data_px2[120], 
        pcx_fpio_data_px2[121], pcx_fpio_data_px2[122], pcx_fpio_data_px2[123]}), .out({SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        pcx_fpio_data_px2_buf1[112], pcx_fpio_data_px2_buf1[113], 
        pcx_fpio_data_px2_buf1[114], pcx_fpio_data_px2_buf1[115], 
        pcx_fpio_data_px2_buf1[116], SYNOPSYS_UNCONNECTED__36, 
        pcx_fpio_data_px2_buf1[118], pcx_fpio_data_px2_buf1[119], 
        pcx_fpio_data_px2_buf1[120], pcx_fpio_data_px2_buf1[121], 
        pcx_fpio_data_px2_buf1[122], pcx_fpio_data_px2_buf1[123]}) );
  fpu_rptr_pcx_fpio_grp16_6 i_pcx_fpio_buf1_2 ( .in({pcx_fpio_data_px2[76], 
        pcx_fpio_data_px2[77], pcx_fpio_data_px2[78], pcx_fpio_data_px2[79], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .out({pcx_fpio_data_px2_buf1[76], pcx_fpio_data_px2_buf1[77], 
        pcx_fpio_data_px2_buf1[78], pcx_fpio_data_px2_buf1[79], 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48}) );
  fpu_rptr_pcx_fpio_grp16_5 i_pcx_fpio_buf1_3 ( .in({pcx_fpio_data_px2[3:0], 
        pcx_fpio_data_px2[64], pcx_fpio_data_px2[65], pcx_fpio_data_px2[66], 
        pcx_fpio_data_px2[67], 1'b0, 1'b0, 1'b0, 1'b0, pcx_fpio_data_px2[72], 
        pcx_fpio_data_px2[73], pcx_fpio_data_px2[74], pcx_fpio_data_px2[75]}), 
        .out({pcx_fpio_data_px2_buf1[3:0], pcx_fpio_data_px2_buf1[64], 
        pcx_fpio_data_px2_buf1[65], pcx_fpio_data_px2_buf1[66], 
        pcx_fpio_data_px2_buf1[67], SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, pcx_fpio_data_px2_buf1[72], 
        pcx_fpio_data_px2_buf1[73], pcx_fpio_data_px2_buf1[74], 
        pcx_fpio_data_px2_buf1[75]}) );
  fpu_rptr_pcx_fpio_grp16_4 i_pcx_fpio_buf1_4 ( .in(pcx_fpio_data_px2[19:4]), 
        .out(pcx_fpio_data_px2_buf1[19:4]) );
  fpu_rptr_pcx_fpio_grp16_3 i_pcx_fpio_buf1_5 ( .in(pcx_fpio_data_px2[35:20]), 
        .out(pcx_fpio_data_px2_buf1[35:20]) );
  fpu_rptr_pcx_fpio_grp16_2 i_pcx_fpio_buf1_6 ( .in({pcx_fpio_data_rdy_px2, 
        pcx_fpio_data_px2[50:36]}), .out({pcx_fpio_data_rdy_px2_buf1, 
        pcx_fpio_data_px2_buf1[50:36]}) );
  fpu_rptr_pcx_fpio_grp16_1 i_pcx_fpio_buf1_7 ( .in({1'b0, 1'b0, 1'b0, 
        pcx_fpio_data_px2[63:51]}), .out({SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        pcx_fpio_data_px2_buf1[63:51]}) );
  fpu_rptr_fp_cpx_grp16_0 i_fp_cpx_buf1_0 ( .in({net211134, net211135, 
        net211136, net211137, fp_cpx_data_ca[134], net211138, net211139, 
        net211140, fp_cpx_req_cq[6], fp_cpx_req_cq[7], fp_cpx_req_cq[3:2], 
        fp_cpx_req_cq[5], fp_cpx_req_cq[1:0], fp_cpx_req_cq[4]}), .out({
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        fp_cpx_data_ca_buf1[134], SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        fp_cpx_req_cq_buf1[6], fp_cpx_req_cq_buf1[7], fp_cpx_req_cq_buf1[3:2], 
        fp_cpx_req_cq_buf1[5], fp_cpx_req_cq_buf1[1:0], fp_cpx_req_cq_buf1[4]}) );
  fpu_rptr_fp_cpx_grp16_9 i_fp_cpx_buf1_1 ( .in({fp_cpx_data_ca[34], 
        fp_cpx_data_ca[36], fp_cpx_data_ca[38], fp_cpx_data_ca[40], 
        fp_cpx_data_ca[42], fp_cpx_data_ca[44], fp_cpx_data_ca[46], 
        fp_cpx_data_ca[48], fp_cpx_data_ca[50], fp_cpx_data_ca[52], 
        fp_cpx_data_ca[54], fp_cpx_data_ca[56], fp_cpx_data_ca[58], 
        fp_cpx_data_ca[60], fp_cpx_data_ca[62], fp_cpx_data_ca[144]}), .out({
        fp_cpx_data_ca_buf1[34], fp_cpx_data_ca_buf1[36], 
        fp_cpx_data_ca_buf1[38], fp_cpx_data_ca_buf1[40], 
        fp_cpx_data_ca_buf1[42], fp_cpx_data_ca_buf1[44], 
        fp_cpx_data_ca_buf1[46], fp_cpx_data_ca_buf1[48], 
        fp_cpx_data_ca_buf1[50], fp_cpx_data_ca_buf1[52], 
        fp_cpx_data_ca_buf1[54], fp_cpx_data_ca_buf1[56], 
        fp_cpx_data_ca_buf1[58], fp_cpx_data_ca_buf1[60], 
        fp_cpx_data_ca_buf1[62], fp_cpx_data_ca_buf1[144]}) );
  fpu_rptr_fp_cpx_grp16_8 i_fp_cpx_buf1_2 ( .in({fp_cpx_data_ca[2], 
        fp_cpx_data_ca[4], fp_cpx_data_ca[6], fp_cpx_data_ca[8], 
        fp_cpx_data_ca[10], fp_cpx_data_ca[12], fp_cpx_data_ca[14], 
        fp_cpx_data_ca[16], fp_cpx_data_ca[18], fp_cpx_data_ca[20], 
        fp_cpx_data_ca[22], fp_cpx_data_ca[24], fp_cpx_data_ca[26], 
        fp_cpx_data_ca[28], fp_cpx_data_ca[30], fp_cpx_data_ca[32]}), .out({
        fp_cpx_data_ca_buf1[2], fp_cpx_data_ca_buf1[4], fp_cpx_data_ca_buf1[6], 
        fp_cpx_data_ca_buf1[8], fp_cpx_data_ca_buf1[10], 
        fp_cpx_data_ca_buf1[12], fp_cpx_data_ca_buf1[14], 
        fp_cpx_data_ca_buf1[16], fp_cpx_data_ca_buf1[18], 
        fp_cpx_data_ca_buf1[20], fp_cpx_data_ca_buf1[22], 
        fp_cpx_data_ca_buf1[24], fp_cpx_data_ca_buf1[26], 
        fp_cpx_data_ca_buf1[28], fp_cpx_data_ca_buf1[30], 
        fp_cpx_data_ca_buf1[32]}) );
  fpu_rptr_fp_cpx_grp16_7 i_fp_cpx_buf1_3 ( .in({fp_cpx_data_ca[31], 
        fp_cpx_data_ca[27], fp_cpx_data_ca[23], fp_cpx_data_ca[25], 
        fp_cpx_data_ca[21], fp_cpx_data_ca[17], fp_cpx_data_ca[19], 
        fp_cpx_data_ca[15], fp_cpx_data_ca[11], fp_cpx_data_ca[13], 
        fp_cpx_data_ca[9], fp_cpx_data_ca[5], fp_cpx_data_ca[7], 
        fp_cpx_data_ca[3], fp_cpx_data_ca[0], fp_cpx_data_ca[1]}), .out({
        fp_cpx_data_ca_buf1[31], fp_cpx_data_ca_buf1[27], 
        fp_cpx_data_ca_buf1[23], fp_cpx_data_ca_buf1[25], 
        fp_cpx_data_ca_buf1[21], fp_cpx_data_ca_buf1[17], 
        fp_cpx_data_ca_buf1[19], fp_cpx_data_ca_buf1[15], 
        fp_cpx_data_ca_buf1[11], fp_cpx_data_ca_buf1[13], 
        fp_cpx_data_ca_buf1[9], fp_cpx_data_ca_buf1[5], fp_cpx_data_ca_buf1[7], 
        fp_cpx_data_ca_buf1[3], fp_cpx_data_ca_buf1[0], fp_cpx_data_ca_buf1[1]}) );
  fpu_rptr_fp_cpx_grp16_6 i_fp_cpx_buf1_4 ( .in({fp_cpx_data_ca[59], 
        fp_cpx_data_ca[61], fp_cpx_data_ca[57], fp_cpx_data_ca[53], 
        fp_cpx_data_ca[55], fp_cpx_data_ca[51], fp_cpx_data_ca[47], 
        fp_cpx_data_ca[49], fp_cpx_data_ca[45], fp_cpx_data_ca[41], 
        fp_cpx_data_ca[43], fp_cpx_data_ca[39], fp_cpx_data_ca[35], 
        fp_cpx_data_ca[37], fp_cpx_data_ca[33], fp_cpx_data_ca[29]}), .out({
        fp_cpx_data_ca_buf1[59], fp_cpx_data_ca_buf1[61], 
        fp_cpx_data_ca_buf1[57], fp_cpx_data_ca_buf1[53], 
        fp_cpx_data_ca_buf1[55], fp_cpx_data_ca_buf1[51], 
        fp_cpx_data_ca_buf1[47], fp_cpx_data_ca_buf1[49], 
        fp_cpx_data_ca_buf1[45], fp_cpx_data_ca_buf1[41], 
        fp_cpx_data_ca_buf1[43], fp_cpx_data_ca_buf1[39], 
        fp_cpx_data_ca_buf1[35], fp_cpx_data_ca_buf1[37], 
        fp_cpx_data_ca_buf1[33], fp_cpx_data_ca_buf1[29]}) );
  fpu_rptr_fp_cpx_grp16_5 i_fp_cpx_buf1_5 ( .in({net211121, net211122, 
        net211123, net211124, net211125, net211126, net211127, net211128, 
        net211129, net211130, fp_cpx_data_ca[135], net211131, net211132, 
        net211133, fp_cpx_data_ca[143], fp_cpx_data_ca[63]}), .out({
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        fp_cpx_data_ca_buf1[135], SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        fp_cpx_data_ca_buf1[143], fp_cpx_data_ca_buf1[63]}) );
  fpu_rptr_fp_cpx_grp16_3 i_fp_cpx_buf1_7 ( .in({net211110, net211111, 
        net211112, net211113, net211114, net211115, net211116, 
        fp_cpx_data_ca[65], fp_cpx_data_ca[67], fp_cpx_data_ca[69], 
        fp_cpx_data_ca[73], net211117, fp_cpx_data_ca[75], net211118, 
        net211119, net211120}), .out({SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        fp_cpx_data_ca_buf1[65], fp_cpx_data_ca_buf1[67], 
        fp_cpx_data_ca_buf1[69], fp_cpx_data_ca_buf1[73], 
        SYNOPSYS_UNCONNECTED__83, fp_cpx_data_ca_buf1[75], 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86}) );
  fpu_rptr_fp_cpx_grp16_1 i_fp_cpx_buf1_9 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, so_buf1, net211106, fp_cpx_data_ca[66], fp_cpx_data_ca[68], 
        net211107, fp_cpx_data_ca[72], fp_cpx_data_ca[74], fp_cpx_data_ca[76], 
        net211108, net211109}), .out({SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, so, SYNOPSYS_UNCONNECTED__93, 
        fp_cpx_data_ca_buf1[66], fp_cpx_data_ca_buf1[68], 
        SYNOPSYS_UNCONNECTED__94, fp_cpx_data_ca_buf1[72], 
        fp_cpx_data_ca_buf1[74], fp_cpx_data_ca_buf1[76], 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96}) );
  fpu_rptr_inq i_inq_sram_din_buf1 ( .in({inq_sram_din_unbuf[155:1], net211105}), .out({inq_sram_din_buf1[155:1], SYNOPSYS_UNCONNECTED__97}) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bw_r_rf16x160_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CGLPPRX2_RVT latch ( .CLK(CLK), .EN(EN), .SE(TE), .GCLK(ENCLK) );
endmodule


module bw_r_rf16x160 ( dout, so_w, so_r, din, rd_adr, wr_adr, read_en, wr_en, 
        rst_tri_en, word_wen, byte_wen, rd_clk, wr_clk, se, si_r, si_w, 
        reset_l, sehold );
  output [159:0] dout;
  input [159:0] din;
  input [3:0] rd_adr;
  input [3:0] wr_adr;
  input [3:0] word_wen;
  input [19:0] byte_wen;
  input read_en, wr_en, rst_tri_en, rd_clk, wr_clk, se, si_r, si_w, reset_l,
         sehold;
  output so_w, so_r;
  wire   wr_en_d1, \inq_ary[15][159] , \inq_ary[15][158] , \inq_ary[15][157] ,
         \inq_ary[15][156] , \inq_ary[15][155] , \inq_ary[15][154] ,
         \inq_ary[15][153] , \inq_ary[15][152] , \inq_ary[15][151] ,
         \inq_ary[15][150] , \inq_ary[15][149] , \inq_ary[15][148] ,
         \inq_ary[15][147] , \inq_ary[15][146] , \inq_ary[15][145] ,
         \inq_ary[15][144] , \inq_ary[15][143] , \inq_ary[15][142] ,
         \inq_ary[15][141] , \inq_ary[15][140] , \inq_ary[15][139] ,
         \inq_ary[15][138] , \inq_ary[15][137] , \inq_ary[15][136] ,
         \inq_ary[15][135] , \inq_ary[15][134] , \inq_ary[15][133] ,
         \inq_ary[15][132] , \inq_ary[15][131] , \inq_ary[15][130] ,
         \inq_ary[15][129] , \inq_ary[15][128] , \inq_ary[15][127] ,
         \inq_ary[15][126] , \inq_ary[15][125] , \inq_ary[15][124] ,
         \inq_ary[15][123] , \inq_ary[15][122] , \inq_ary[15][121] ,
         \inq_ary[15][120] , \inq_ary[15][119] , \inq_ary[15][118] ,
         \inq_ary[15][117] , \inq_ary[15][116] , \inq_ary[15][115] ,
         \inq_ary[15][114] , \inq_ary[15][113] , \inq_ary[15][112] ,
         \inq_ary[15][111] , \inq_ary[15][110] , \inq_ary[15][109] ,
         \inq_ary[15][108] , \inq_ary[15][107] , \inq_ary[15][106] ,
         \inq_ary[15][105] , \inq_ary[15][104] , \inq_ary[15][103] ,
         \inq_ary[15][102] , \inq_ary[15][101] , \inq_ary[15][100] ,
         \inq_ary[15][99] , \inq_ary[15][98] , \inq_ary[15][97] ,
         \inq_ary[15][96] , \inq_ary[15][95] , \inq_ary[15][94] ,
         \inq_ary[15][93] , \inq_ary[15][92] , \inq_ary[15][91] ,
         \inq_ary[15][90] , \inq_ary[15][89] , \inq_ary[15][88] ,
         \inq_ary[15][87] , \inq_ary[15][86] , \inq_ary[15][85] ,
         \inq_ary[15][84] , \inq_ary[15][83] , \inq_ary[15][82] ,
         \inq_ary[15][81] , \inq_ary[15][80] , \inq_ary[15][79] ,
         \inq_ary[15][78] , \inq_ary[15][77] , \inq_ary[15][76] ,
         \inq_ary[15][75] , \inq_ary[15][74] , \inq_ary[15][73] ,
         \inq_ary[15][72] , \inq_ary[15][71] , \inq_ary[15][70] ,
         \inq_ary[15][69] , \inq_ary[15][68] , \inq_ary[15][67] ,
         \inq_ary[15][66] , \inq_ary[15][65] , \inq_ary[15][64] ,
         \inq_ary[15][63] , \inq_ary[15][62] , \inq_ary[15][61] ,
         \inq_ary[15][60] , \inq_ary[15][59] , \inq_ary[15][58] ,
         \inq_ary[15][57] , \inq_ary[15][56] , \inq_ary[15][55] ,
         \inq_ary[15][54] , \inq_ary[15][53] , \inq_ary[15][52] ,
         \inq_ary[15][51] , \inq_ary[15][50] , \inq_ary[15][49] ,
         \inq_ary[15][48] , \inq_ary[15][47] , \inq_ary[15][46] ,
         \inq_ary[15][45] , \inq_ary[15][44] , \inq_ary[15][43] ,
         \inq_ary[15][42] , \inq_ary[15][41] , \inq_ary[15][40] ,
         \inq_ary[15][39] , \inq_ary[15][38] , \inq_ary[15][37] ,
         \inq_ary[15][36] , \inq_ary[15][35] , \inq_ary[15][34] ,
         \inq_ary[15][33] , \inq_ary[15][32] , \inq_ary[15][31] ,
         \inq_ary[15][30] , \inq_ary[15][29] , \inq_ary[15][28] ,
         \inq_ary[15][27] , \inq_ary[15][26] , \inq_ary[15][25] ,
         \inq_ary[15][24] , \inq_ary[15][23] , \inq_ary[15][22] ,
         \inq_ary[15][21] , \inq_ary[15][20] , \inq_ary[15][19] ,
         \inq_ary[15][18] , \inq_ary[15][17] , \inq_ary[15][16] ,
         \inq_ary[15][15] , \inq_ary[15][14] , \inq_ary[15][13] ,
         \inq_ary[15][12] , \inq_ary[15][11] , \inq_ary[15][10] ,
         \inq_ary[15][9] , \inq_ary[15][8] , \inq_ary[15][7] ,
         \inq_ary[15][6] , \inq_ary[15][5] , \inq_ary[14][159] ,
         \inq_ary[14][158] , \inq_ary[14][157] , \inq_ary[14][156] ,
         \inq_ary[14][155] , \inq_ary[14][154] , \inq_ary[14][153] ,
         \inq_ary[14][152] , \inq_ary[14][151] , \inq_ary[14][150] ,
         \inq_ary[14][149] , \inq_ary[14][148] , \inq_ary[14][147] ,
         \inq_ary[14][146] , \inq_ary[14][145] , \inq_ary[14][144] ,
         \inq_ary[14][143] , \inq_ary[14][142] , \inq_ary[14][141] ,
         \inq_ary[14][140] , \inq_ary[14][139] , \inq_ary[14][138] ,
         \inq_ary[14][137] , \inq_ary[14][136] , \inq_ary[14][135] ,
         \inq_ary[14][134] , \inq_ary[14][133] , \inq_ary[14][132] ,
         \inq_ary[14][131] , \inq_ary[14][130] , \inq_ary[14][129] ,
         \inq_ary[14][128] , \inq_ary[14][127] , \inq_ary[14][126] ,
         \inq_ary[14][125] , \inq_ary[14][124] , \inq_ary[14][123] ,
         \inq_ary[14][122] , \inq_ary[14][121] , \inq_ary[14][120] ,
         \inq_ary[14][119] , \inq_ary[14][118] , \inq_ary[14][117] ,
         \inq_ary[14][116] , \inq_ary[14][115] , \inq_ary[14][114] ,
         \inq_ary[14][113] , \inq_ary[14][112] , \inq_ary[14][111] ,
         \inq_ary[14][110] , \inq_ary[14][109] , \inq_ary[14][108] ,
         \inq_ary[14][107] , \inq_ary[14][106] , \inq_ary[14][105] ,
         \inq_ary[14][104] , \inq_ary[14][103] , \inq_ary[14][102] ,
         \inq_ary[14][101] , \inq_ary[14][100] , \inq_ary[14][99] ,
         \inq_ary[14][98] , \inq_ary[14][97] , \inq_ary[14][96] ,
         \inq_ary[14][95] , \inq_ary[14][94] , \inq_ary[14][93] ,
         \inq_ary[14][92] , \inq_ary[14][91] , \inq_ary[14][90] ,
         \inq_ary[14][89] , \inq_ary[14][88] , \inq_ary[14][87] ,
         \inq_ary[14][86] , \inq_ary[14][85] , \inq_ary[14][84] ,
         \inq_ary[14][83] , \inq_ary[14][82] , \inq_ary[14][81] ,
         \inq_ary[14][80] , \inq_ary[14][79] , \inq_ary[14][78] ,
         \inq_ary[14][77] , \inq_ary[14][76] , \inq_ary[14][75] ,
         \inq_ary[14][74] , \inq_ary[14][73] , \inq_ary[14][72] ,
         \inq_ary[14][71] , \inq_ary[14][70] , \inq_ary[14][69] ,
         \inq_ary[14][68] , \inq_ary[14][67] , \inq_ary[14][66] ,
         \inq_ary[14][65] , \inq_ary[14][64] , \inq_ary[14][63] ,
         \inq_ary[14][62] , \inq_ary[14][61] , \inq_ary[14][60] ,
         \inq_ary[14][59] , \inq_ary[14][58] , \inq_ary[14][57] ,
         \inq_ary[14][56] , \inq_ary[14][55] , \inq_ary[14][54] ,
         \inq_ary[14][53] , \inq_ary[14][52] , \inq_ary[14][51] ,
         \inq_ary[14][50] , \inq_ary[14][49] , \inq_ary[14][48] ,
         \inq_ary[14][47] , \inq_ary[14][46] , \inq_ary[14][45] ,
         \inq_ary[14][44] , \inq_ary[14][43] , \inq_ary[14][42] ,
         \inq_ary[14][41] , \inq_ary[14][40] , \inq_ary[14][39] ,
         \inq_ary[14][38] , \inq_ary[14][37] , \inq_ary[14][36] ,
         \inq_ary[14][35] , \inq_ary[14][34] , \inq_ary[14][33] ,
         \inq_ary[14][32] , \inq_ary[14][31] , \inq_ary[14][30] ,
         \inq_ary[14][29] , \inq_ary[14][28] , \inq_ary[14][27] ,
         \inq_ary[14][26] , \inq_ary[14][25] , \inq_ary[14][24] ,
         \inq_ary[14][23] , \inq_ary[14][22] , \inq_ary[14][21] ,
         \inq_ary[14][20] , \inq_ary[14][19] , \inq_ary[14][18] ,
         \inq_ary[14][17] , \inq_ary[14][16] , \inq_ary[14][15] ,
         \inq_ary[14][14] , \inq_ary[14][13] , \inq_ary[14][12] ,
         \inq_ary[14][11] , \inq_ary[14][10] , \inq_ary[14][9] ,
         \inq_ary[14][8] , \inq_ary[14][7] , \inq_ary[14][6] ,
         \inq_ary[14][5] , \inq_ary[13][159] , \inq_ary[13][158] ,
         \inq_ary[13][157] , \inq_ary[13][156] , \inq_ary[13][155] ,
         \inq_ary[13][154] , \inq_ary[13][153] , \inq_ary[13][152] ,
         \inq_ary[13][151] , \inq_ary[13][150] , \inq_ary[13][149] ,
         \inq_ary[13][148] , \inq_ary[13][147] , \inq_ary[13][146] ,
         \inq_ary[13][145] , \inq_ary[13][144] , \inq_ary[13][143] ,
         \inq_ary[13][142] , \inq_ary[13][141] , \inq_ary[13][140] ,
         \inq_ary[13][139] , \inq_ary[13][138] , \inq_ary[13][137] ,
         \inq_ary[13][136] , \inq_ary[13][135] , \inq_ary[13][134] ,
         \inq_ary[13][133] , \inq_ary[13][132] , \inq_ary[13][131] ,
         \inq_ary[13][130] , \inq_ary[13][129] , \inq_ary[13][128] ,
         \inq_ary[13][127] , \inq_ary[13][126] , \inq_ary[13][125] ,
         \inq_ary[13][124] , \inq_ary[13][123] , \inq_ary[13][122] ,
         \inq_ary[13][121] , \inq_ary[13][120] , \inq_ary[13][119] ,
         \inq_ary[13][118] , \inq_ary[13][117] , \inq_ary[13][116] ,
         \inq_ary[13][115] , \inq_ary[13][114] , \inq_ary[13][113] ,
         \inq_ary[13][112] , \inq_ary[13][111] , \inq_ary[13][110] ,
         \inq_ary[13][109] , \inq_ary[13][108] , \inq_ary[13][107] ,
         \inq_ary[13][106] , \inq_ary[13][105] , \inq_ary[13][104] ,
         \inq_ary[13][103] , \inq_ary[13][102] , \inq_ary[13][101] ,
         \inq_ary[13][100] , \inq_ary[13][99] , \inq_ary[13][98] ,
         \inq_ary[13][97] , \inq_ary[13][96] , \inq_ary[13][95] ,
         \inq_ary[13][94] , \inq_ary[13][93] , \inq_ary[13][92] ,
         \inq_ary[13][91] , \inq_ary[13][90] , \inq_ary[13][89] ,
         \inq_ary[13][88] , \inq_ary[13][87] , \inq_ary[13][86] ,
         \inq_ary[13][85] , \inq_ary[13][84] , \inq_ary[13][83] ,
         \inq_ary[13][82] , \inq_ary[13][81] , \inq_ary[13][80] ,
         \inq_ary[13][79] , \inq_ary[13][78] , \inq_ary[13][77] ,
         \inq_ary[13][76] , \inq_ary[13][75] , \inq_ary[13][74] ,
         \inq_ary[13][73] , \inq_ary[13][72] , \inq_ary[13][71] ,
         \inq_ary[13][70] , \inq_ary[13][69] , \inq_ary[13][68] ,
         \inq_ary[13][67] , \inq_ary[13][66] , \inq_ary[13][65] ,
         \inq_ary[13][64] , \inq_ary[13][63] , \inq_ary[13][62] ,
         \inq_ary[13][61] , \inq_ary[13][60] , \inq_ary[13][59] ,
         \inq_ary[13][58] , \inq_ary[13][57] , \inq_ary[13][56] ,
         \inq_ary[13][55] , \inq_ary[13][54] , \inq_ary[13][53] ,
         \inq_ary[13][52] , \inq_ary[13][51] , \inq_ary[13][50] ,
         \inq_ary[13][49] , \inq_ary[13][48] , \inq_ary[13][47] ,
         \inq_ary[13][46] , \inq_ary[13][45] , \inq_ary[13][44] ,
         \inq_ary[13][43] , \inq_ary[13][42] , \inq_ary[13][41] ,
         \inq_ary[13][40] , \inq_ary[13][39] , \inq_ary[13][38] ,
         \inq_ary[13][37] , \inq_ary[13][36] , \inq_ary[13][35] ,
         \inq_ary[13][34] , \inq_ary[13][33] , \inq_ary[13][32] ,
         \inq_ary[13][31] , \inq_ary[13][30] , \inq_ary[13][29] ,
         \inq_ary[13][28] , \inq_ary[13][27] , \inq_ary[13][26] ,
         \inq_ary[13][25] , \inq_ary[13][24] , \inq_ary[13][23] ,
         \inq_ary[13][22] , \inq_ary[13][21] , \inq_ary[13][20] ,
         \inq_ary[13][19] , \inq_ary[13][18] , \inq_ary[13][17] ,
         \inq_ary[13][16] , \inq_ary[13][15] , \inq_ary[13][14] ,
         \inq_ary[13][13] , \inq_ary[13][12] , \inq_ary[13][11] ,
         \inq_ary[13][10] , \inq_ary[13][9] , \inq_ary[13][8] ,
         \inq_ary[13][7] , \inq_ary[13][6] , \inq_ary[13][5] ,
         \inq_ary[12][159] , \inq_ary[12][158] , \inq_ary[12][157] ,
         \inq_ary[12][156] , \inq_ary[12][155] , \inq_ary[12][154] ,
         \inq_ary[12][153] , \inq_ary[12][152] , \inq_ary[12][151] ,
         \inq_ary[12][150] , \inq_ary[12][149] , \inq_ary[12][148] ,
         \inq_ary[12][147] , \inq_ary[12][146] , \inq_ary[12][145] ,
         \inq_ary[12][144] , \inq_ary[12][143] , \inq_ary[12][142] ,
         \inq_ary[12][141] , \inq_ary[12][140] , \inq_ary[12][139] ,
         \inq_ary[12][138] , \inq_ary[12][137] , \inq_ary[12][136] ,
         \inq_ary[12][135] , \inq_ary[12][134] , \inq_ary[12][133] ,
         \inq_ary[12][132] , \inq_ary[12][131] , \inq_ary[12][130] ,
         \inq_ary[12][129] , \inq_ary[12][128] , \inq_ary[12][127] ,
         \inq_ary[12][126] , \inq_ary[12][125] , \inq_ary[12][124] ,
         \inq_ary[12][123] , \inq_ary[12][122] , \inq_ary[12][121] ,
         \inq_ary[12][120] , \inq_ary[12][119] , \inq_ary[12][118] ,
         \inq_ary[12][117] , \inq_ary[12][116] , \inq_ary[12][115] ,
         \inq_ary[12][114] , \inq_ary[12][113] , \inq_ary[12][112] ,
         \inq_ary[12][111] , \inq_ary[12][110] , \inq_ary[12][109] ,
         \inq_ary[12][108] , \inq_ary[12][107] , \inq_ary[12][106] ,
         \inq_ary[12][105] , \inq_ary[12][104] , \inq_ary[12][103] ,
         \inq_ary[12][102] , \inq_ary[12][101] , \inq_ary[12][100] ,
         \inq_ary[12][99] , \inq_ary[12][98] , \inq_ary[12][97] ,
         \inq_ary[12][96] , \inq_ary[12][95] , \inq_ary[12][94] ,
         \inq_ary[12][93] , \inq_ary[12][92] , \inq_ary[12][91] ,
         \inq_ary[12][90] , \inq_ary[12][89] , \inq_ary[12][88] ,
         \inq_ary[12][87] , \inq_ary[12][86] , \inq_ary[12][85] ,
         \inq_ary[12][84] , \inq_ary[12][83] , \inq_ary[12][82] ,
         \inq_ary[12][81] , \inq_ary[12][80] , \inq_ary[12][79] ,
         \inq_ary[12][78] , \inq_ary[12][77] , \inq_ary[12][76] ,
         \inq_ary[12][75] , \inq_ary[12][74] , \inq_ary[12][73] ,
         \inq_ary[12][72] , \inq_ary[12][71] , \inq_ary[12][70] ,
         \inq_ary[12][69] , \inq_ary[12][68] , \inq_ary[12][67] ,
         \inq_ary[12][66] , \inq_ary[12][65] , \inq_ary[12][64] ,
         \inq_ary[12][63] , \inq_ary[12][62] , \inq_ary[12][61] ,
         \inq_ary[12][60] , \inq_ary[12][59] , \inq_ary[12][58] ,
         \inq_ary[12][57] , \inq_ary[12][56] , \inq_ary[12][55] ,
         \inq_ary[12][54] , \inq_ary[12][53] , \inq_ary[12][52] ,
         \inq_ary[12][51] , \inq_ary[12][50] , \inq_ary[12][49] ,
         \inq_ary[12][48] , \inq_ary[12][47] , \inq_ary[12][46] ,
         \inq_ary[12][45] , \inq_ary[12][44] , \inq_ary[12][43] ,
         \inq_ary[12][42] , \inq_ary[12][41] , \inq_ary[12][40] ,
         \inq_ary[12][39] , \inq_ary[12][38] , \inq_ary[12][37] ,
         \inq_ary[12][36] , \inq_ary[12][35] , \inq_ary[12][34] ,
         \inq_ary[12][33] , \inq_ary[12][32] , \inq_ary[12][31] ,
         \inq_ary[12][30] , \inq_ary[12][29] , \inq_ary[12][28] ,
         \inq_ary[12][27] , \inq_ary[12][26] , \inq_ary[12][25] ,
         \inq_ary[12][24] , \inq_ary[12][23] , \inq_ary[12][22] ,
         \inq_ary[12][21] , \inq_ary[12][20] , \inq_ary[12][19] ,
         \inq_ary[12][18] , \inq_ary[12][17] , \inq_ary[12][16] ,
         \inq_ary[12][15] , \inq_ary[12][14] , \inq_ary[12][13] ,
         \inq_ary[12][12] , \inq_ary[12][11] , \inq_ary[12][10] ,
         \inq_ary[12][9] , \inq_ary[12][8] , \inq_ary[12][7] ,
         \inq_ary[12][6] , \inq_ary[12][5] , \inq_ary[11][159] ,
         \inq_ary[11][158] , \inq_ary[11][157] , \inq_ary[11][156] ,
         \inq_ary[11][155] , \inq_ary[11][154] , \inq_ary[11][153] ,
         \inq_ary[11][152] , \inq_ary[11][151] , \inq_ary[11][150] ,
         \inq_ary[11][149] , \inq_ary[11][148] , \inq_ary[11][147] ,
         \inq_ary[11][146] , \inq_ary[11][145] , \inq_ary[11][144] ,
         \inq_ary[11][143] , \inq_ary[11][142] , \inq_ary[11][141] ,
         \inq_ary[11][140] , \inq_ary[11][139] , \inq_ary[11][138] ,
         \inq_ary[11][137] , \inq_ary[11][136] , \inq_ary[11][135] ,
         \inq_ary[11][134] , \inq_ary[11][133] , \inq_ary[11][132] ,
         \inq_ary[11][131] , \inq_ary[11][130] , \inq_ary[11][129] ,
         \inq_ary[11][128] , \inq_ary[11][127] , \inq_ary[11][126] ,
         \inq_ary[11][125] , \inq_ary[11][124] , \inq_ary[11][123] ,
         \inq_ary[11][122] , \inq_ary[11][121] , \inq_ary[11][120] ,
         \inq_ary[11][119] , \inq_ary[11][118] , \inq_ary[11][117] ,
         \inq_ary[11][116] , \inq_ary[11][115] , \inq_ary[11][114] ,
         \inq_ary[11][113] , \inq_ary[11][112] , \inq_ary[11][111] ,
         \inq_ary[11][110] , \inq_ary[11][109] , \inq_ary[11][108] ,
         \inq_ary[11][107] , \inq_ary[11][106] , \inq_ary[11][105] ,
         \inq_ary[11][104] , \inq_ary[11][103] , \inq_ary[11][102] ,
         \inq_ary[11][101] , \inq_ary[11][100] , \inq_ary[11][99] ,
         \inq_ary[11][98] , \inq_ary[11][97] , \inq_ary[11][96] ,
         \inq_ary[11][95] , \inq_ary[11][94] , \inq_ary[11][93] ,
         \inq_ary[11][92] , \inq_ary[11][91] , \inq_ary[11][90] ,
         \inq_ary[11][89] , \inq_ary[11][88] , \inq_ary[11][87] ,
         \inq_ary[11][86] , \inq_ary[11][85] , \inq_ary[11][84] ,
         \inq_ary[11][83] , \inq_ary[11][82] , \inq_ary[11][81] ,
         \inq_ary[11][80] , \inq_ary[11][79] , \inq_ary[11][78] ,
         \inq_ary[11][77] , \inq_ary[11][76] , \inq_ary[11][75] ,
         \inq_ary[11][74] , \inq_ary[11][73] , \inq_ary[11][72] ,
         \inq_ary[11][71] , \inq_ary[11][70] , \inq_ary[11][69] ,
         \inq_ary[11][68] , \inq_ary[11][67] , \inq_ary[11][66] ,
         \inq_ary[11][65] , \inq_ary[11][64] , \inq_ary[11][63] ,
         \inq_ary[11][62] , \inq_ary[11][61] , \inq_ary[11][60] ,
         \inq_ary[11][59] , \inq_ary[11][58] , \inq_ary[11][57] ,
         \inq_ary[11][56] , \inq_ary[11][55] , \inq_ary[11][54] ,
         \inq_ary[11][53] , \inq_ary[11][52] , \inq_ary[11][51] ,
         \inq_ary[11][50] , \inq_ary[11][49] , \inq_ary[11][48] ,
         \inq_ary[11][47] , \inq_ary[11][46] , \inq_ary[11][45] ,
         \inq_ary[11][44] , \inq_ary[11][43] , \inq_ary[11][42] ,
         \inq_ary[11][41] , \inq_ary[11][40] , \inq_ary[11][39] ,
         \inq_ary[11][38] , \inq_ary[11][37] , \inq_ary[11][36] ,
         \inq_ary[11][35] , \inq_ary[11][34] , \inq_ary[11][33] ,
         \inq_ary[11][32] , \inq_ary[11][31] , \inq_ary[11][30] ,
         \inq_ary[11][29] , \inq_ary[11][28] , \inq_ary[11][27] ,
         \inq_ary[11][26] , \inq_ary[11][25] , \inq_ary[11][24] ,
         \inq_ary[11][23] , \inq_ary[11][22] , \inq_ary[11][21] ,
         \inq_ary[11][20] , \inq_ary[11][19] , \inq_ary[11][18] ,
         \inq_ary[11][17] , \inq_ary[11][16] , \inq_ary[11][15] ,
         \inq_ary[11][14] , \inq_ary[11][13] , \inq_ary[11][12] ,
         \inq_ary[11][11] , \inq_ary[11][10] , \inq_ary[11][9] ,
         \inq_ary[11][8] , \inq_ary[11][7] , \inq_ary[11][6] ,
         \inq_ary[11][5] , \inq_ary[10][159] , \inq_ary[10][158] ,
         \inq_ary[10][157] , \inq_ary[10][156] , \inq_ary[10][155] ,
         \inq_ary[10][154] , \inq_ary[10][153] , \inq_ary[10][152] ,
         \inq_ary[10][151] , \inq_ary[10][150] , \inq_ary[10][149] ,
         \inq_ary[10][148] , \inq_ary[10][147] , \inq_ary[10][146] ,
         \inq_ary[10][145] , \inq_ary[10][144] , \inq_ary[10][143] ,
         \inq_ary[10][142] , \inq_ary[10][141] , \inq_ary[10][140] ,
         \inq_ary[10][139] , \inq_ary[10][138] , \inq_ary[10][137] ,
         \inq_ary[10][136] , \inq_ary[10][135] , \inq_ary[10][134] ,
         \inq_ary[10][133] , \inq_ary[10][132] , \inq_ary[10][131] ,
         \inq_ary[10][130] , \inq_ary[10][129] , \inq_ary[10][128] ,
         \inq_ary[10][127] , \inq_ary[10][126] , \inq_ary[10][125] ,
         \inq_ary[10][124] , \inq_ary[10][123] , \inq_ary[10][122] ,
         \inq_ary[10][121] , \inq_ary[10][120] , \inq_ary[10][119] ,
         \inq_ary[10][118] , \inq_ary[10][117] , \inq_ary[10][116] ,
         \inq_ary[10][115] , \inq_ary[10][114] , \inq_ary[10][113] ,
         \inq_ary[10][112] , \inq_ary[10][111] , \inq_ary[10][110] ,
         \inq_ary[10][109] , \inq_ary[10][108] , \inq_ary[10][107] ,
         \inq_ary[10][106] , \inq_ary[10][105] , \inq_ary[10][104] ,
         \inq_ary[10][103] , \inq_ary[10][102] , \inq_ary[10][101] ,
         \inq_ary[10][100] , \inq_ary[10][99] , \inq_ary[10][98] ,
         \inq_ary[10][97] , \inq_ary[10][96] , \inq_ary[10][95] ,
         \inq_ary[10][94] , \inq_ary[10][93] , \inq_ary[10][92] ,
         \inq_ary[10][91] , \inq_ary[10][90] , \inq_ary[10][89] ,
         \inq_ary[10][88] , \inq_ary[10][87] , \inq_ary[10][86] ,
         \inq_ary[10][85] , \inq_ary[10][84] , \inq_ary[10][83] ,
         \inq_ary[10][82] , \inq_ary[10][81] , \inq_ary[10][80] ,
         \inq_ary[10][79] , \inq_ary[10][78] , \inq_ary[10][77] ,
         \inq_ary[10][76] , \inq_ary[10][75] , \inq_ary[10][74] ,
         \inq_ary[10][73] , \inq_ary[10][72] , \inq_ary[10][71] ,
         \inq_ary[10][70] , \inq_ary[10][69] , \inq_ary[10][68] ,
         \inq_ary[10][67] , \inq_ary[10][66] , \inq_ary[10][65] ,
         \inq_ary[10][64] , \inq_ary[10][63] , \inq_ary[10][62] ,
         \inq_ary[10][61] , \inq_ary[10][60] , \inq_ary[10][59] ,
         \inq_ary[10][58] , \inq_ary[10][57] , \inq_ary[10][56] ,
         \inq_ary[10][55] , \inq_ary[10][54] , \inq_ary[10][53] ,
         \inq_ary[10][52] , \inq_ary[10][51] , \inq_ary[10][50] ,
         \inq_ary[10][49] , \inq_ary[10][48] , \inq_ary[10][47] ,
         \inq_ary[10][46] , \inq_ary[10][45] , \inq_ary[10][44] ,
         \inq_ary[10][43] , \inq_ary[10][42] , \inq_ary[10][41] ,
         \inq_ary[10][40] , \inq_ary[10][39] , \inq_ary[10][38] ,
         \inq_ary[10][37] , \inq_ary[10][36] , \inq_ary[10][35] ,
         \inq_ary[10][34] , \inq_ary[10][33] , \inq_ary[10][32] ,
         \inq_ary[10][31] , \inq_ary[10][30] , \inq_ary[10][29] ,
         \inq_ary[10][28] , \inq_ary[10][27] , \inq_ary[10][26] ,
         \inq_ary[10][25] , \inq_ary[10][24] , \inq_ary[10][23] ,
         \inq_ary[10][22] , \inq_ary[10][21] , \inq_ary[10][20] ,
         \inq_ary[10][19] , \inq_ary[10][18] , \inq_ary[10][17] ,
         \inq_ary[10][16] , \inq_ary[10][15] , \inq_ary[10][14] ,
         \inq_ary[10][13] , \inq_ary[10][12] , \inq_ary[10][11] ,
         \inq_ary[10][10] , \inq_ary[10][9] , \inq_ary[10][8] ,
         \inq_ary[10][7] , \inq_ary[10][6] , \inq_ary[10][5] ,
         \inq_ary[9][159] , \inq_ary[9][158] , \inq_ary[9][157] ,
         \inq_ary[9][156] , \inq_ary[9][155] , \inq_ary[9][154] ,
         \inq_ary[9][153] , \inq_ary[9][152] , \inq_ary[9][151] ,
         \inq_ary[9][150] , \inq_ary[9][149] , \inq_ary[9][148] ,
         \inq_ary[9][147] , \inq_ary[9][146] , \inq_ary[9][145] ,
         \inq_ary[9][144] , \inq_ary[9][143] , \inq_ary[9][142] ,
         \inq_ary[9][141] , \inq_ary[9][140] , \inq_ary[9][139] ,
         \inq_ary[9][138] , \inq_ary[9][137] , \inq_ary[9][136] ,
         \inq_ary[9][135] , \inq_ary[9][134] , \inq_ary[9][133] ,
         \inq_ary[9][132] , \inq_ary[9][131] , \inq_ary[9][130] ,
         \inq_ary[9][129] , \inq_ary[9][128] , \inq_ary[9][127] ,
         \inq_ary[9][126] , \inq_ary[9][125] , \inq_ary[9][124] ,
         \inq_ary[9][123] , \inq_ary[9][122] , \inq_ary[9][121] ,
         \inq_ary[9][120] , \inq_ary[9][119] , \inq_ary[9][118] ,
         \inq_ary[9][117] , \inq_ary[9][116] , \inq_ary[9][115] ,
         \inq_ary[9][114] , \inq_ary[9][113] , \inq_ary[9][112] ,
         \inq_ary[9][111] , \inq_ary[9][110] , \inq_ary[9][109] ,
         \inq_ary[9][108] , \inq_ary[9][107] , \inq_ary[9][106] ,
         \inq_ary[9][105] , \inq_ary[9][104] , \inq_ary[9][103] ,
         \inq_ary[9][102] , \inq_ary[9][101] , \inq_ary[9][100] ,
         \inq_ary[9][99] , \inq_ary[9][98] , \inq_ary[9][97] ,
         \inq_ary[9][96] , \inq_ary[9][95] , \inq_ary[9][94] ,
         \inq_ary[9][93] , \inq_ary[9][92] , \inq_ary[9][91] ,
         \inq_ary[9][90] , \inq_ary[9][89] , \inq_ary[9][88] ,
         \inq_ary[9][87] , \inq_ary[9][86] , \inq_ary[9][85] ,
         \inq_ary[9][84] , \inq_ary[9][83] , \inq_ary[9][82] ,
         \inq_ary[9][81] , \inq_ary[9][80] , \inq_ary[9][79] ,
         \inq_ary[9][78] , \inq_ary[9][77] , \inq_ary[9][76] ,
         \inq_ary[9][75] , \inq_ary[9][74] , \inq_ary[9][73] ,
         \inq_ary[9][72] , \inq_ary[9][71] , \inq_ary[9][70] ,
         \inq_ary[9][69] , \inq_ary[9][68] , \inq_ary[9][67] ,
         \inq_ary[9][66] , \inq_ary[9][65] , \inq_ary[9][64] ,
         \inq_ary[9][63] , \inq_ary[9][62] , \inq_ary[9][61] ,
         \inq_ary[9][60] , \inq_ary[9][59] , \inq_ary[9][58] ,
         \inq_ary[9][57] , \inq_ary[9][56] , \inq_ary[9][55] ,
         \inq_ary[9][54] , \inq_ary[9][53] , \inq_ary[9][52] ,
         \inq_ary[9][51] , \inq_ary[9][50] , \inq_ary[9][49] ,
         \inq_ary[9][48] , \inq_ary[9][47] , \inq_ary[9][46] ,
         \inq_ary[9][45] , \inq_ary[9][44] , \inq_ary[9][43] ,
         \inq_ary[9][42] , \inq_ary[9][41] , \inq_ary[9][40] ,
         \inq_ary[9][39] , \inq_ary[9][38] , \inq_ary[9][37] ,
         \inq_ary[9][36] , \inq_ary[9][35] , \inq_ary[9][34] ,
         \inq_ary[9][33] , \inq_ary[9][32] , \inq_ary[9][31] ,
         \inq_ary[9][30] , \inq_ary[9][29] , \inq_ary[9][28] ,
         \inq_ary[9][27] , \inq_ary[9][26] , \inq_ary[9][25] ,
         \inq_ary[9][24] , \inq_ary[9][23] , \inq_ary[9][22] ,
         \inq_ary[9][21] , \inq_ary[9][20] , \inq_ary[9][19] ,
         \inq_ary[9][18] , \inq_ary[9][17] , \inq_ary[9][16] ,
         \inq_ary[9][15] , \inq_ary[9][14] , \inq_ary[9][13] ,
         \inq_ary[9][12] , \inq_ary[9][11] , \inq_ary[9][10] , \inq_ary[9][9] ,
         \inq_ary[9][8] , \inq_ary[9][7] , \inq_ary[9][6] , \inq_ary[9][5] ,
         \inq_ary[8][159] , \inq_ary[8][158] , \inq_ary[8][157] ,
         \inq_ary[8][156] , \inq_ary[8][155] , \inq_ary[8][154] ,
         \inq_ary[8][153] , \inq_ary[8][152] , \inq_ary[8][151] ,
         \inq_ary[8][150] , \inq_ary[8][149] , \inq_ary[8][148] ,
         \inq_ary[8][147] , \inq_ary[8][146] , \inq_ary[8][145] ,
         \inq_ary[8][144] , \inq_ary[8][143] , \inq_ary[8][142] ,
         \inq_ary[8][141] , \inq_ary[8][140] , \inq_ary[8][139] ,
         \inq_ary[8][138] , \inq_ary[8][137] , \inq_ary[8][136] ,
         \inq_ary[8][135] , \inq_ary[8][134] , \inq_ary[8][133] ,
         \inq_ary[8][132] , \inq_ary[8][131] , \inq_ary[8][130] ,
         \inq_ary[8][129] , \inq_ary[8][128] , \inq_ary[8][127] ,
         \inq_ary[8][126] , \inq_ary[8][125] , \inq_ary[8][124] ,
         \inq_ary[8][123] , \inq_ary[8][122] , \inq_ary[8][121] ,
         \inq_ary[8][120] , \inq_ary[8][119] , \inq_ary[8][118] ,
         \inq_ary[8][117] , \inq_ary[8][116] , \inq_ary[8][115] ,
         \inq_ary[8][114] , \inq_ary[8][113] , \inq_ary[8][112] ,
         \inq_ary[8][111] , \inq_ary[8][110] , \inq_ary[8][109] ,
         \inq_ary[8][108] , \inq_ary[8][107] , \inq_ary[8][106] ,
         \inq_ary[8][105] , \inq_ary[8][104] , \inq_ary[8][103] ,
         \inq_ary[8][102] , \inq_ary[8][101] , \inq_ary[8][100] ,
         \inq_ary[8][99] , \inq_ary[8][98] , \inq_ary[8][97] ,
         \inq_ary[8][96] , \inq_ary[8][95] , \inq_ary[8][94] ,
         \inq_ary[8][93] , \inq_ary[8][92] , \inq_ary[8][91] ,
         \inq_ary[8][90] , \inq_ary[8][89] , \inq_ary[8][88] ,
         \inq_ary[8][87] , \inq_ary[8][86] , \inq_ary[8][85] ,
         \inq_ary[8][84] , \inq_ary[8][83] , \inq_ary[8][82] ,
         \inq_ary[8][81] , \inq_ary[8][80] , \inq_ary[8][79] ,
         \inq_ary[8][78] , \inq_ary[8][77] , \inq_ary[8][76] ,
         \inq_ary[8][75] , \inq_ary[8][74] , \inq_ary[8][73] ,
         \inq_ary[8][72] , \inq_ary[8][71] , \inq_ary[8][70] ,
         \inq_ary[8][69] , \inq_ary[8][68] , \inq_ary[8][67] ,
         \inq_ary[8][66] , \inq_ary[8][65] , \inq_ary[8][64] ,
         \inq_ary[8][63] , \inq_ary[8][62] , \inq_ary[8][61] ,
         \inq_ary[8][60] , \inq_ary[8][59] , \inq_ary[8][58] ,
         \inq_ary[8][57] , \inq_ary[8][56] , \inq_ary[8][55] ,
         \inq_ary[8][54] , \inq_ary[8][53] , \inq_ary[8][52] ,
         \inq_ary[8][51] , \inq_ary[8][50] , \inq_ary[8][49] ,
         \inq_ary[8][48] , \inq_ary[8][47] , \inq_ary[8][46] ,
         \inq_ary[8][45] , \inq_ary[8][44] , \inq_ary[8][43] ,
         \inq_ary[8][42] , \inq_ary[8][41] , \inq_ary[8][40] ,
         \inq_ary[8][39] , \inq_ary[8][38] , \inq_ary[8][37] ,
         \inq_ary[8][36] , \inq_ary[8][35] , \inq_ary[8][34] ,
         \inq_ary[8][33] , \inq_ary[8][32] , \inq_ary[8][31] ,
         \inq_ary[8][30] , \inq_ary[8][29] , \inq_ary[8][28] ,
         \inq_ary[8][27] , \inq_ary[8][26] , \inq_ary[8][25] ,
         \inq_ary[8][24] , \inq_ary[8][23] , \inq_ary[8][22] ,
         \inq_ary[8][21] , \inq_ary[8][20] , \inq_ary[8][19] ,
         \inq_ary[8][18] , \inq_ary[8][17] , \inq_ary[8][16] ,
         \inq_ary[8][15] , \inq_ary[8][14] , \inq_ary[8][13] ,
         \inq_ary[8][12] , \inq_ary[8][11] , \inq_ary[8][10] , \inq_ary[8][9] ,
         \inq_ary[8][8] , \inq_ary[8][7] , \inq_ary[8][6] , \inq_ary[8][5] ,
         \inq_ary[7][159] , \inq_ary[7][158] , \inq_ary[7][157] ,
         \inq_ary[7][156] , \inq_ary[7][155] , \inq_ary[7][154] ,
         \inq_ary[7][153] , \inq_ary[7][152] , \inq_ary[7][151] ,
         \inq_ary[7][150] , \inq_ary[7][149] , \inq_ary[7][148] ,
         \inq_ary[7][147] , \inq_ary[7][146] , \inq_ary[7][145] ,
         \inq_ary[7][144] , \inq_ary[7][143] , \inq_ary[7][142] ,
         \inq_ary[7][141] , \inq_ary[7][140] , \inq_ary[7][139] ,
         \inq_ary[7][138] , \inq_ary[7][137] , \inq_ary[7][136] ,
         \inq_ary[7][135] , \inq_ary[7][134] , \inq_ary[7][133] ,
         \inq_ary[7][132] , \inq_ary[7][131] , \inq_ary[7][130] ,
         \inq_ary[7][129] , \inq_ary[7][128] , \inq_ary[7][127] ,
         \inq_ary[7][126] , \inq_ary[7][125] , \inq_ary[7][124] ,
         \inq_ary[7][123] , \inq_ary[7][122] , \inq_ary[7][121] ,
         \inq_ary[7][120] , \inq_ary[7][119] , \inq_ary[7][118] ,
         \inq_ary[7][117] , \inq_ary[7][116] , \inq_ary[7][115] ,
         \inq_ary[7][114] , \inq_ary[7][113] , \inq_ary[7][112] ,
         \inq_ary[7][111] , \inq_ary[7][110] , \inq_ary[7][109] ,
         \inq_ary[7][108] , \inq_ary[7][107] , \inq_ary[7][106] ,
         \inq_ary[7][105] , \inq_ary[7][104] , \inq_ary[7][103] ,
         \inq_ary[7][102] , \inq_ary[7][101] , \inq_ary[7][100] ,
         \inq_ary[7][99] , \inq_ary[7][98] , \inq_ary[7][97] ,
         \inq_ary[7][96] , \inq_ary[7][95] , \inq_ary[7][94] ,
         \inq_ary[7][93] , \inq_ary[7][92] , \inq_ary[7][91] ,
         \inq_ary[7][90] , \inq_ary[7][89] , \inq_ary[7][88] ,
         \inq_ary[7][87] , \inq_ary[7][86] , \inq_ary[7][85] ,
         \inq_ary[7][84] , \inq_ary[7][83] , \inq_ary[7][82] ,
         \inq_ary[7][81] , \inq_ary[7][80] , \inq_ary[7][79] ,
         \inq_ary[7][78] , \inq_ary[7][77] , \inq_ary[7][76] ,
         \inq_ary[7][75] , \inq_ary[7][74] , \inq_ary[7][73] ,
         \inq_ary[7][72] , \inq_ary[7][71] , \inq_ary[7][70] ,
         \inq_ary[7][69] , \inq_ary[7][68] , \inq_ary[7][67] ,
         \inq_ary[7][66] , \inq_ary[7][65] , \inq_ary[7][64] ,
         \inq_ary[7][63] , \inq_ary[7][62] , \inq_ary[7][61] ,
         \inq_ary[7][60] , \inq_ary[7][59] , \inq_ary[7][58] ,
         \inq_ary[7][57] , \inq_ary[7][56] , \inq_ary[7][55] ,
         \inq_ary[7][54] , \inq_ary[7][53] , \inq_ary[7][52] ,
         \inq_ary[7][51] , \inq_ary[7][50] , \inq_ary[7][49] ,
         \inq_ary[7][48] , \inq_ary[7][47] , \inq_ary[7][46] ,
         \inq_ary[7][45] , \inq_ary[7][44] , \inq_ary[7][43] ,
         \inq_ary[7][42] , \inq_ary[7][41] , \inq_ary[7][40] ,
         \inq_ary[7][39] , \inq_ary[7][38] , \inq_ary[7][37] ,
         \inq_ary[7][36] , \inq_ary[7][35] , \inq_ary[7][34] ,
         \inq_ary[7][33] , \inq_ary[7][32] , \inq_ary[7][31] ,
         \inq_ary[7][30] , \inq_ary[7][29] , \inq_ary[7][28] ,
         \inq_ary[7][27] , \inq_ary[7][26] , \inq_ary[7][25] ,
         \inq_ary[7][24] , \inq_ary[7][23] , \inq_ary[7][22] ,
         \inq_ary[7][21] , \inq_ary[7][20] , \inq_ary[7][19] ,
         \inq_ary[7][18] , \inq_ary[7][17] , \inq_ary[7][16] ,
         \inq_ary[7][15] , \inq_ary[7][14] , \inq_ary[7][13] ,
         \inq_ary[7][12] , \inq_ary[7][11] , \inq_ary[7][10] , \inq_ary[7][9] ,
         \inq_ary[7][8] , \inq_ary[7][7] , \inq_ary[7][6] , \inq_ary[7][5] ,
         \inq_ary[6][159] , \inq_ary[6][158] , \inq_ary[6][157] ,
         \inq_ary[6][156] , \inq_ary[6][155] , \inq_ary[6][154] ,
         \inq_ary[6][153] , \inq_ary[6][152] , \inq_ary[6][151] ,
         \inq_ary[6][150] , \inq_ary[6][149] , \inq_ary[6][148] ,
         \inq_ary[6][147] , \inq_ary[6][146] , \inq_ary[6][145] ,
         \inq_ary[6][144] , \inq_ary[6][143] , \inq_ary[6][142] ,
         \inq_ary[6][141] , \inq_ary[6][140] , \inq_ary[6][139] ,
         \inq_ary[6][138] , \inq_ary[6][137] , \inq_ary[6][136] ,
         \inq_ary[6][135] , \inq_ary[6][134] , \inq_ary[6][133] ,
         \inq_ary[6][132] , \inq_ary[6][131] , \inq_ary[6][130] ,
         \inq_ary[6][129] , \inq_ary[6][128] , \inq_ary[6][127] ,
         \inq_ary[6][126] , \inq_ary[6][125] , \inq_ary[6][124] ,
         \inq_ary[6][123] , \inq_ary[6][122] , \inq_ary[6][121] ,
         \inq_ary[6][120] , \inq_ary[6][119] , \inq_ary[6][118] ,
         \inq_ary[6][117] , \inq_ary[6][116] , \inq_ary[6][115] ,
         \inq_ary[6][114] , \inq_ary[6][113] , \inq_ary[6][112] ,
         \inq_ary[6][111] , \inq_ary[6][110] , \inq_ary[6][109] ,
         \inq_ary[6][108] , \inq_ary[6][107] , \inq_ary[6][106] ,
         \inq_ary[6][105] , \inq_ary[6][104] , \inq_ary[6][103] ,
         \inq_ary[6][102] , \inq_ary[6][101] , \inq_ary[6][100] ,
         \inq_ary[6][99] , \inq_ary[6][98] , \inq_ary[6][97] ,
         \inq_ary[6][96] , \inq_ary[6][95] , \inq_ary[6][94] ,
         \inq_ary[6][93] , \inq_ary[6][92] , \inq_ary[6][91] ,
         \inq_ary[6][90] , \inq_ary[6][89] , \inq_ary[6][88] ,
         \inq_ary[6][87] , \inq_ary[6][86] , \inq_ary[6][85] ,
         \inq_ary[6][84] , \inq_ary[6][83] , \inq_ary[6][82] ,
         \inq_ary[6][81] , \inq_ary[6][80] , \inq_ary[6][79] ,
         \inq_ary[6][78] , \inq_ary[6][77] , \inq_ary[6][76] ,
         \inq_ary[6][75] , \inq_ary[6][74] , \inq_ary[6][73] ,
         \inq_ary[6][72] , \inq_ary[6][71] , \inq_ary[6][70] ,
         \inq_ary[6][69] , \inq_ary[6][68] , \inq_ary[6][67] ,
         \inq_ary[6][66] , \inq_ary[6][65] , \inq_ary[6][64] ,
         \inq_ary[6][63] , \inq_ary[6][62] , \inq_ary[6][61] ,
         \inq_ary[6][60] , \inq_ary[6][59] , \inq_ary[6][58] ,
         \inq_ary[6][57] , \inq_ary[6][56] , \inq_ary[6][55] ,
         \inq_ary[6][54] , \inq_ary[6][53] , \inq_ary[6][52] ,
         \inq_ary[6][51] , \inq_ary[6][50] , \inq_ary[6][49] ,
         \inq_ary[6][48] , \inq_ary[6][47] , \inq_ary[6][46] ,
         \inq_ary[6][45] , \inq_ary[6][44] , \inq_ary[6][43] ,
         \inq_ary[6][42] , \inq_ary[6][41] , \inq_ary[6][40] ,
         \inq_ary[6][39] , \inq_ary[6][38] , \inq_ary[6][37] ,
         \inq_ary[6][36] , \inq_ary[6][35] , \inq_ary[6][34] ,
         \inq_ary[6][33] , \inq_ary[6][32] , \inq_ary[6][31] ,
         \inq_ary[6][30] , \inq_ary[6][29] , \inq_ary[6][28] ,
         \inq_ary[6][27] , \inq_ary[6][26] , \inq_ary[6][25] ,
         \inq_ary[6][24] , \inq_ary[6][23] , \inq_ary[6][22] ,
         \inq_ary[6][21] , \inq_ary[6][20] , \inq_ary[6][19] ,
         \inq_ary[6][18] , \inq_ary[6][17] , \inq_ary[6][16] ,
         \inq_ary[6][15] , \inq_ary[6][14] , \inq_ary[6][13] ,
         \inq_ary[6][12] , \inq_ary[6][11] , \inq_ary[6][10] , \inq_ary[6][9] ,
         \inq_ary[6][8] , \inq_ary[6][7] , \inq_ary[6][6] , \inq_ary[6][5] ,
         \inq_ary[5][159] , \inq_ary[5][158] , \inq_ary[5][157] ,
         \inq_ary[5][156] , \inq_ary[5][155] , \inq_ary[5][154] ,
         \inq_ary[5][153] , \inq_ary[5][152] , \inq_ary[5][151] ,
         \inq_ary[5][150] , \inq_ary[5][149] , \inq_ary[5][148] ,
         \inq_ary[5][147] , \inq_ary[5][146] , \inq_ary[5][145] ,
         \inq_ary[5][144] , \inq_ary[5][143] , \inq_ary[5][142] ,
         \inq_ary[5][141] , \inq_ary[5][140] , \inq_ary[5][139] ,
         \inq_ary[5][138] , \inq_ary[5][137] , \inq_ary[5][136] ,
         \inq_ary[5][135] , \inq_ary[5][134] , \inq_ary[5][133] ,
         \inq_ary[5][132] , \inq_ary[5][131] , \inq_ary[5][130] ,
         \inq_ary[5][129] , \inq_ary[5][128] , \inq_ary[5][127] ,
         \inq_ary[5][126] , \inq_ary[5][125] , \inq_ary[5][124] ,
         \inq_ary[5][123] , \inq_ary[5][122] , \inq_ary[5][121] ,
         \inq_ary[5][120] , \inq_ary[5][119] , \inq_ary[5][118] ,
         \inq_ary[5][117] , \inq_ary[5][116] , \inq_ary[5][115] ,
         \inq_ary[5][114] , \inq_ary[5][113] , \inq_ary[5][112] ,
         \inq_ary[5][111] , \inq_ary[5][110] , \inq_ary[5][109] ,
         \inq_ary[5][108] , \inq_ary[5][107] , \inq_ary[5][106] ,
         \inq_ary[5][105] , \inq_ary[5][104] , \inq_ary[5][103] ,
         \inq_ary[5][102] , \inq_ary[5][101] , \inq_ary[5][100] ,
         \inq_ary[5][99] , \inq_ary[5][98] , \inq_ary[5][97] ,
         \inq_ary[5][96] , \inq_ary[5][95] , \inq_ary[5][94] ,
         \inq_ary[5][93] , \inq_ary[5][92] , \inq_ary[5][91] ,
         \inq_ary[5][90] , \inq_ary[5][89] , \inq_ary[5][88] ,
         \inq_ary[5][87] , \inq_ary[5][86] , \inq_ary[5][85] ,
         \inq_ary[5][84] , \inq_ary[5][83] , \inq_ary[5][82] ,
         \inq_ary[5][81] , \inq_ary[5][80] , \inq_ary[5][79] ,
         \inq_ary[5][78] , \inq_ary[5][77] , \inq_ary[5][76] ,
         \inq_ary[5][75] , \inq_ary[5][74] , \inq_ary[5][73] ,
         \inq_ary[5][72] , \inq_ary[5][71] , \inq_ary[5][70] ,
         \inq_ary[5][69] , \inq_ary[5][68] , \inq_ary[5][67] ,
         \inq_ary[5][66] , \inq_ary[5][65] , \inq_ary[5][64] ,
         \inq_ary[5][63] , \inq_ary[5][62] , \inq_ary[5][61] ,
         \inq_ary[5][60] , \inq_ary[5][59] , \inq_ary[5][58] ,
         \inq_ary[5][57] , \inq_ary[5][56] , \inq_ary[5][55] ,
         \inq_ary[5][54] , \inq_ary[5][53] , \inq_ary[5][52] ,
         \inq_ary[5][51] , \inq_ary[5][50] , \inq_ary[5][49] ,
         \inq_ary[5][48] , \inq_ary[5][47] , \inq_ary[5][46] ,
         \inq_ary[5][45] , \inq_ary[5][44] , \inq_ary[5][43] ,
         \inq_ary[5][42] , \inq_ary[5][41] , \inq_ary[5][40] ,
         \inq_ary[5][39] , \inq_ary[5][38] , \inq_ary[5][37] ,
         \inq_ary[5][36] , \inq_ary[5][35] , \inq_ary[5][34] ,
         \inq_ary[5][33] , \inq_ary[5][32] , \inq_ary[5][31] ,
         \inq_ary[5][30] , \inq_ary[5][29] , \inq_ary[5][28] ,
         \inq_ary[5][27] , \inq_ary[5][26] , \inq_ary[5][25] ,
         \inq_ary[5][24] , \inq_ary[5][23] , \inq_ary[5][22] ,
         \inq_ary[5][21] , \inq_ary[5][20] , \inq_ary[5][19] ,
         \inq_ary[5][18] , \inq_ary[5][17] , \inq_ary[5][16] ,
         \inq_ary[5][15] , \inq_ary[5][14] , \inq_ary[5][13] ,
         \inq_ary[5][12] , \inq_ary[5][11] , \inq_ary[5][10] , \inq_ary[5][9] ,
         \inq_ary[5][8] , \inq_ary[5][7] , \inq_ary[5][6] , \inq_ary[5][5] ,
         \inq_ary[4][159] , \inq_ary[4][158] , \inq_ary[4][157] ,
         \inq_ary[4][156] , \inq_ary[4][155] , \inq_ary[4][154] ,
         \inq_ary[4][153] , \inq_ary[4][152] , \inq_ary[4][151] ,
         \inq_ary[4][150] , \inq_ary[4][149] , \inq_ary[4][148] ,
         \inq_ary[4][147] , \inq_ary[4][146] , \inq_ary[4][145] ,
         \inq_ary[4][144] , \inq_ary[4][143] , \inq_ary[4][142] ,
         \inq_ary[4][141] , \inq_ary[4][140] , \inq_ary[4][139] ,
         \inq_ary[4][138] , \inq_ary[4][137] , \inq_ary[4][136] ,
         \inq_ary[4][135] , \inq_ary[4][134] , \inq_ary[4][133] ,
         \inq_ary[4][132] , \inq_ary[4][131] , \inq_ary[4][130] ,
         \inq_ary[4][129] , \inq_ary[4][128] , \inq_ary[4][127] ,
         \inq_ary[4][126] , \inq_ary[4][125] , \inq_ary[4][124] ,
         \inq_ary[4][123] , \inq_ary[4][122] , \inq_ary[4][121] ,
         \inq_ary[4][120] , \inq_ary[4][119] , \inq_ary[4][118] ,
         \inq_ary[4][117] , \inq_ary[4][116] , \inq_ary[4][115] ,
         \inq_ary[4][114] , \inq_ary[4][113] , \inq_ary[4][112] ,
         \inq_ary[4][111] , \inq_ary[4][110] , \inq_ary[4][109] ,
         \inq_ary[4][108] , \inq_ary[4][107] , \inq_ary[4][106] ,
         \inq_ary[4][105] , \inq_ary[4][104] , \inq_ary[4][103] ,
         \inq_ary[4][102] , \inq_ary[4][101] , \inq_ary[4][100] ,
         \inq_ary[4][99] , \inq_ary[4][98] , \inq_ary[4][97] ,
         \inq_ary[4][96] , \inq_ary[4][95] , \inq_ary[4][94] ,
         \inq_ary[4][93] , \inq_ary[4][92] , \inq_ary[4][91] ,
         \inq_ary[4][90] , \inq_ary[4][89] , \inq_ary[4][88] ,
         \inq_ary[4][87] , \inq_ary[4][86] , \inq_ary[4][85] ,
         \inq_ary[4][84] , \inq_ary[4][83] , \inq_ary[4][82] ,
         \inq_ary[4][81] , \inq_ary[4][80] , \inq_ary[4][79] ,
         \inq_ary[4][78] , \inq_ary[4][77] , \inq_ary[4][76] ,
         \inq_ary[4][75] , \inq_ary[4][74] , \inq_ary[4][73] ,
         \inq_ary[4][72] , \inq_ary[4][71] , \inq_ary[4][70] ,
         \inq_ary[4][69] , \inq_ary[4][68] , \inq_ary[4][67] ,
         \inq_ary[4][66] , \inq_ary[4][65] , \inq_ary[4][64] ,
         \inq_ary[4][63] , \inq_ary[4][62] , \inq_ary[4][61] ,
         \inq_ary[4][60] , \inq_ary[4][59] , \inq_ary[4][58] ,
         \inq_ary[4][57] , \inq_ary[4][56] , \inq_ary[4][55] ,
         \inq_ary[4][54] , \inq_ary[4][53] , \inq_ary[4][52] ,
         \inq_ary[4][51] , \inq_ary[4][50] , \inq_ary[4][49] ,
         \inq_ary[4][48] , \inq_ary[4][47] , \inq_ary[4][46] ,
         \inq_ary[4][45] , \inq_ary[4][44] , \inq_ary[4][43] ,
         \inq_ary[4][42] , \inq_ary[4][41] , \inq_ary[4][40] ,
         \inq_ary[4][39] , \inq_ary[4][38] , \inq_ary[4][37] ,
         \inq_ary[4][36] , \inq_ary[4][35] , \inq_ary[4][34] ,
         \inq_ary[4][33] , \inq_ary[4][32] , \inq_ary[4][31] ,
         \inq_ary[4][30] , \inq_ary[4][29] , \inq_ary[4][28] ,
         \inq_ary[4][27] , \inq_ary[4][26] , \inq_ary[4][25] ,
         \inq_ary[4][24] , \inq_ary[4][23] , \inq_ary[4][22] ,
         \inq_ary[4][21] , \inq_ary[4][20] , \inq_ary[4][19] ,
         \inq_ary[4][18] , \inq_ary[4][17] , \inq_ary[4][16] ,
         \inq_ary[4][15] , \inq_ary[4][14] , \inq_ary[4][13] ,
         \inq_ary[4][12] , \inq_ary[4][11] , \inq_ary[4][10] , \inq_ary[4][9] ,
         \inq_ary[4][8] , \inq_ary[4][7] , \inq_ary[4][6] , \inq_ary[4][5] ,
         \inq_ary[3][159] , \inq_ary[3][158] , \inq_ary[3][157] ,
         \inq_ary[3][156] , \inq_ary[3][155] , \inq_ary[3][154] ,
         \inq_ary[3][153] , \inq_ary[3][152] , \inq_ary[3][151] ,
         \inq_ary[3][150] , \inq_ary[3][149] , \inq_ary[3][148] ,
         \inq_ary[3][147] , \inq_ary[3][146] , \inq_ary[3][145] ,
         \inq_ary[3][144] , \inq_ary[3][143] , \inq_ary[3][142] ,
         \inq_ary[3][141] , \inq_ary[3][140] , \inq_ary[3][139] ,
         \inq_ary[3][138] , \inq_ary[3][137] , \inq_ary[3][136] ,
         \inq_ary[3][135] , \inq_ary[3][134] , \inq_ary[3][133] ,
         \inq_ary[3][132] , \inq_ary[3][131] , \inq_ary[3][130] ,
         \inq_ary[3][129] , \inq_ary[3][128] , \inq_ary[3][127] ,
         \inq_ary[3][126] , \inq_ary[3][125] , \inq_ary[3][124] ,
         \inq_ary[3][123] , \inq_ary[3][122] , \inq_ary[3][121] ,
         \inq_ary[3][120] , \inq_ary[3][119] , \inq_ary[3][118] ,
         \inq_ary[3][117] , \inq_ary[3][116] , \inq_ary[3][115] ,
         \inq_ary[3][114] , \inq_ary[3][113] , \inq_ary[3][112] ,
         \inq_ary[3][111] , \inq_ary[3][110] , \inq_ary[3][109] ,
         \inq_ary[3][108] , \inq_ary[3][107] , \inq_ary[3][106] ,
         \inq_ary[3][105] , \inq_ary[3][104] , \inq_ary[3][103] ,
         \inq_ary[3][102] , \inq_ary[3][101] , \inq_ary[3][100] ,
         \inq_ary[3][99] , \inq_ary[3][98] , \inq_ary[3][97] ,
         \inq_ary[3][96] , \inq_ary[3][95] , \inq_ary[3][94] ,
         \inq_ary[3][93] , \inq_ary[3][92] , \inq_ary[3][91] ,
         \inq_ary[3][90] , \inq_ary[3][89] , \inq_ary[3][88] ,
         \inq_ary[3][87] , \inq_ary[3][86] , \inq_ary[3][85] ,
         \inq_ary[3][84] , \inq_ary[3][83] , \inq_ary[3][82] ,
         \inq_ary[3][81] , \inq_ary[3][80] , \inq_ary[3][79] ,
         \inq_ary[3][78] , \inq_ary[3][77] , \inq_ary[3][76] ,
         \inq_ary[3][75] , \inq_ary[3][74] , \inq_ary[3][73] ,
         \inq_ary[3][72] , \inq_ary[3][71] , \inq_ary[3][70] ,
         \inq_ary[3][69] , \inq_ary[3][68] , \inq_ary[3][67] ,
         \inq_ary[3][66] , \inq_ary[3][65] , \inq_ary[3][64] ,
         \inq_ary[3][63] , \inq_ary[3][62] , \inq_ary[3][61] ,
         \inq_ary[3][60] , \inq_ary[3][59] , \inq_ary[3][58] ,
         \inq_ary[3][57] , \inq_ary[3][56] , \inq_ary[3][55] ,
         \inq_ary[3][54] , \inq_ary[3][53] , \inq_ary[3][52] ,
         \inq_ary[3][51] , \inq_ary[3][50] , \inq_ary[3][49] ,
         \inq_ary[3][48] , \inq_ary[3][47] , \inq_ary[3][46] ,
         \inq_ary[3][45] , \inq_ary[3][44] , \inq_ary[3][43] ,
         \inq_ary[3][42] , \inq_ary[3][41] , \inq_ary[3][40] ,
         \inq_ary[3][39] , \inq_ary[3][38] , \inq_ary[3][37] ,
         \inq_ary[3][36] , \inq_ary[3][35] , \inq_ary[3][34] ,
         \inq_ary[3][33] , \inq_ary[3][32] , \inq_ary[3][31] ,
         \inq_ary[3][30] , \inq_ary[3][29] , \inq_ary[3][28] ,
         \inq_ary[3][27] , \inq_ary[3][26] , \inq_ary[3][25] ,
         \inq_ary[3][24] , \inq_ary[3][23] , \inq_ary[3][22] ,
         \inq_ary[3][21] , \inq_ary[3][20] , \inq_ary[3][19] ,
         \inq_ary[3][18] , \inq_ary[3][17] , \inq_ary[3][16] ,
         \inq_ary[3][15] , \inq_ary[3][14] , \inq_ary[3][13] ,
         \inq_ary[3][12] , \inq_ary[3][11] , \inq_ary[3][10] , \inq_ary[3][9] ,
         \inq_ary[3][8] , \inq_ary[3][7] , \inq_ary[3][6] , \inq_ary[3][5] ,
         \inq_ary[2][159] , \inq_ary[2][158] , \inq_ary[2][157] ,
         \inq_ary[2][156] , \inq_ary[2][155] , \inq_ary[2][154] ,
         \inq_ary[2][153] , \inq_ary[2][152] , \inq_ary[2][151] ,
         \inq_ary[2][150] , \inq_ary[2][149] , \inq_ary[2][148] ,
         \inq_ary[2][147] , \inq_ary[2][146] , \inq_ary[2][145] ,
         \inq_ary[2][144] , \inq_ary[2][143] , \inq_ary[2][142] ,
         \inq_ary[2][141] , \inq_ary[2][140] , \inq_ary[2][139] ,
         \inq_ary[2][138] , \inq_ary[2][137] , \inq_ary[2][136] ,
         \inq_ary[2][135] , \inq_ary[2][134] , \inq_ary[2][133] ,
         \inq_ary[2][132] , \inq_ary[2][131] , \inq_ary[2][130] ,
         \inq_ary[2][129] , \inq_ary[2][128] , \inq_ary[2][127] ,
         \inq_ary[2][126] , \inq_ary[2][125] , \inq_ary[2][124] ,
         \inq_ary[2][123] , \inq_ary[2][122] , \inq_ary[2][121] ,
         \inq_ary[2][120] , \inq_ary[2][119] , \inq_ary[2][118] ,
         \inq_ary[2][117] , \inq_ary[2][116] , \inq_ary[2][115] ,
         \inq_ary[2][114] , \inq_ary[2][113] , \inq_ary[2][112] ,
         \inq_ary[2][111] , \inq_ary[2][110] , \inq_ary[2][109] ,
         \inq_ary[2][108] , \inq_ary[2][107] , \inq_ary[2][106] ,
         \inq_ary[2][105] , \inq_ary[2][104] , \inq_ary[2][103] ,
         \inq_ary[2][102] , \inq_ary[2][101] , \inq_ary[2][100] ,
         \inq_ary[2][99] , \inq_ary[2][98] , \inq_ary[2][97] ,
         \inq_ary[2][96] , \inq_ary[2][95] , \inq_ary[2][94] ,
         \inq_ary[2][93] , \inq_ary[2][92] , \inq_ary[2][91] ,
         \inq_ary[2][90] , \inq_ary[2][89] , \inq_ary[2][88] ,
         \inq_ary[2][87] , \inq_ary[2][86] , \inq_ary[2][85] ,
         \inq_ary[2][84] , \inq_ary[2][83] , \inq_ary[2][82] ,
         \inq_ary[2][81] , \inq_ary[2][80] , \inq_ary[2][79] ,
         \inq_ary[2][78] , \inq_ary[2][77] , \inq_ary[2][76] ,
         \inq_ary[2][75] , \inq_ary[2][74] , \inq_ary[2][73] ,
         \inq_ary[2][72] , \inq_ary[2][71] , \inq_ary[2][70] ,
         \inq_ary[2][69] , \inq_ary[2][68] , \inq_ary[2][67] ,
         \inq_ary[2][66] , \inq_ary[2][65] , \inq_ary[2][64] ,
         \inq_ary[2][63] , \inq_ary[2][62] , \inq_ary[2][61] ,
         \inq_ary[2][60] , \inq_ary[2][59] , \inq_ary[2][58] ,
         \inq_ary[2][57] , \inq_ary[2][56] , \inq_ary[2][55] ,
         \inq_ary[2][54] , \inq_ary[2][53] , \inq_ary[2][52] ,
         \inq_ary[2][51] , \inq_ary[2][50] , \inq_ary[2][49] ,
         \inq_ary[2][48] , \inq_ary[2][47] , \inq_ary[2][46] ,
         \inq_ary[2][45] , \inq_ary[2][44] , \inq_ary[2][43] ,
         \inq_ary[2][42] , \inq_ary[2][41] , \inq_ary[2][40] ,
         \inq_ary[2][39] , \inq_ary[2][38] , \inq_ary[2][37] ,
         \inq_ary[2][36] , \inq_ary[2][35] , \inq_ary[2][34] ,
         \inq_ary[2][33] , \inq_ary[2][32] , \inq_ary[2][31] ,
         \inq_ary[2][30] , \inq_ary[2][29] , \inq_ary[2][28] ,
         \inq_ary[2][27] , \inq_ary[2][26] , \inq_ary[2][25] ,
         \inq_ary[2][24] , \inq_ary[2][23] , \inq_ary[2][22] ,
         \inq_ary[2][21] , \inq_ary[2][20] , \inq_ary[2][19] ,
         \inq_ary[2][18] , \inq_ary[2][17] , \inq_ary[2][16] ,
         \inq_ary[2][15] , \inq_ary[2][14] , \inq_ary[2][13] ,
         \inq_ary[2][12] , \inq_ary[2][11] , \inq_ary[2][10] , \inq_ary[2][9] ,
         \inq_ary[2][8] , \inq_ary[2][7] , \inq_ary[2][6] , \inq_ary[2][5] ,
         \inq_ary[1][159] , \inq_ary[1][158] , \inq_ary[1][157] ,
         \inq_ary[1][156] , \inq_ary[1][155] , \inq_ary[1][154] ,
         \inq_ary[1][153] , \inq_ary[1][152] , \inq_ary[1][151] ,
         \inq_ary[1][150] , \inq_ary[1][149] , \inq_ary[1][148] ,
         \inq_ary[1][147] , \inq_ary[1][146] , \inq_ary[1][145] ,
         \inq_ary[1][144] , \inq_ary[1][143] , \inq_ary[1][142] ,
         \inq_ary[1][141] , \inq_ary[1][140] , \inq_ary[1][139] ,
         \inq_ary[1][138] , \inq_ary[1][137] , \inq_ary[1][136] ,
         \inq_ary[1][135] , \inq_ary[1][134] , \inq_ary[1][133] ,
         \inq_ary[1][132] , \inq_ary[1][131] , \inq_ary[1][130] ,
         \inq_ary[1][129] , \inq_ary[1][128] , \inq_ary[1][127] ,
         \inq_ary[1][126] , \inq_ary[1][125] , \inq_ary[1][124] ,
         \inq_ary[1][123] , \inq_ary[1][122] , \inq_ary[1][121] ,
         \inq_ary[1][120] , \inq_ary[1][119] , \inq_ary[1][118] ,
         \inq_ary[1][117] , \inq_ary[1][116] , \inq_ary[1][115] ,
         \inq_ary[1][114] , \inq_ary[1][113] , \inq_ary[1][112] ,
         \inq_ary[1][111] , \inq_ary[1][110] , \inq_ary[1][109] ,
         \inq_ary[1][108] , \inq_ary[1][107] , \inq_ary[1][106] ,
         \inq_ary[1][105] , \inq_ary[1][104] , \inq_ary[1][103] ,
         \inq_ary[1][102] , \inq_ary[1][101] , \inq_ary[1][100] ,
         \inq_ary[1][99] , \inq_ary[1][98] , \inq_ary[1][97] ,
         \inq_ary[1][96] , \inq_ary[1][95] , \inq_ary[1][94] ,
         \inq_ary[1][93] , \inq_ary[1][92] , \inq_ary[1][91] ,
         \inq_ary[1][90] , \inq_ary[1][89] , \inq_ary[1][88] ,
         \inq_ary[1][87] , \inq_ary[1][86] , \inq_ary[1][85] ,
         \inq_ary[1][84] , \inq_ary[1][83] , \inq_ary[1][82] ,
         \inq_ary[1][81] , \inq_ary[1][80] , \inq_ary[1][79] ,
         \inq_ary[1][78] , \inq_ary[1][77] , \inq_ary[1][76] ,
         \inq_ary[1][75] , \inq_ary[1][74] , \inq_ary[1][73] ,
         \inq_ary[1][72] , \inq_ary[1][71] , \inq_ary[1][70] ,
         \inq_ary[1][69] , \inq_ary[1][68] , \inq_ary[1][67] ,
         \inq_ary[1][66] , \inq_ary[1][65] , \inq_ary[1][64] ,
         \inq_ary[1][63] , \inq_ary[1][62] , \inq_ary[1][61] ,
         \inq_ary[1][60] , \inq_ary[1][59] , \inq_ary[1][58] ,
         \inq_ary[1][57] , \inq_ary[1][56] , \inq_ary[1][55] ,
         \inq_ary[1][54] , \inq_ary[1][53] , \inq_ary[1][52] ,
         \inq_ary[1][51] , \inq_ary[1][50] , \inq_ary[1][49] ,
         \inq_ary[1][48] , \inq_ary[1][47] , \inq_ary[1][46] ,
         \inq_ary[1][45] , \inq_ary[1][44] , \inq_ary[1][43] ,
         \inq_ary[1][42] , \inq_ary[1][41] , \inq_ary[1][40] ,
         \inq_ary[1][39] , \inq_ary[1][38] , \inq_ary[1][37] ,
         \inq_ary[1][36] , \inq_ary[1][35] , \inq_ary[1][34] ,
         \inq_ary[1][33] , \inq_ary[1][32] , \inq_ary[1][31] ,
         \inq_ary[1][30] , \inq_ary[1][29] , \inq_ary[1][28] ,
         \inq_ary[1][27] , \inq_ary[1][26] , \inq_ary[1][25] ,
         \inq_ary[1][24] , \inq_ary[1][23] , \inq_ary[1][22] ,
         \inq_ary[1][21] , \inq_ary[1][20] , \inq_ary[1][19] ,
         \inq_ary[1][18] , \inq_ary[1][17] , \inq_ary[1][16] ,
         \inq_ary[1][15] , \inq_ary[1][14] , \inq_ary[1][13] ,
         \inq_ary[1][12] , \inq_ary[1][11] , \inq_ary[1][10] , \inq_ary[1][9] ,
         \inq_ary[1][8] , \inq_ary[1][7] , \inq_ary[1][6] , \inq_ary[1][5] ,
         \inq_ary[0][159] , \inq_ary[0][158] , \inq_ary[0][157] ,
         \inq_ary[0][156] , \inq_ary[0][155] , \inq_ary[0][154] ,
         \inq_ary[0][153] , \inq_ary[0][152] , \inq_ary[0][151] ,
         \inq_ary[0][150] , \inq_ary[0][149] , \inq_ary[0][148] ,
         \inq_ary[0][147] , \inq_ary[0][146] , \inq_ary[0][145] ,
         \inq_ary[0][144] , \inq_ary[0][143] , \inq_ary[0][142] ,
         \inq_ary[0][141] , \inq_ary[0][140] , \inq_ary[0][139] ,
         \inq_ary[0][138] , \inq_ary[0][137] , \inq_ary[0][136] ,
         \inq_ary[0][135] , \inq_ary[0][134] , \inq_ary[0][133] ,
         \inq_ary[0][132] , \inq_ary[0][131] , \inq_ary[0][130] ,
         \inq_ary[0][129] , \inq_ary[0][128] , \inq_ary[0][127] ,
         \inq_ary[0][126] , \inq_ary[0][125] , \inq_ary[0][124] ,
         \inq_ary[0][123] , \inq_ary[0][122] , \inq_ary[0][121] ,
         \inq_ary[0][120] , \inq_ary[0][119] , \inq_ary[0][118] ,
         \inq_ary[0][117] , \inq_ary[0][116] , \inq_ary[0][115] ,
         \inq_ary[0][114] , \inq_ary[0][113] , \inq_ary[0][112] ,
         \inq_ary[0][111] , \inq_ary[0][110] , \inq_ary[0][109] ,
         \inq_ary[0][108] , \inq_ary[0][107] , \inq_ary[0][106] ,
         \inq_ary[0][105] , \inq_ary[0][104] , \inq_ary[0][103] ,
         \inq_ary[0][102] , \inq_ary[0][101] , \inq_ary[0][100] ,
         \inq_ary[0][99] , \inq_ary[0][98] , \inq_ary[0][97] ,
         \inq_ary[0][96] , \inq_ary[0][95] , \inq_ary[0][94] ,
         \inq_ary[0][93] , \inq_ary[0][92] , \inq_ary[0][91] ,
         \inq_ary[0][90] , \inq_ary[0][89] , \inq_ary[0][88] ,
         \inq_ary[0][87] , \inq_ary[0][86] , \inq_ary[0][85] ,
         \inq_ary[0][84] , \inq_ary[0][83] , \inq_ary[0][82] ,
         \inq_ary[0][81] , \inq_ary[0][80] , \inq_ary[0][79] ,
         \inq_ary[0][78] , \inq_ary[0][77] , \inq_ary[0][76] ,
         \inq_ary[0][75] , \inq_ary[0][74] , \inq_ary[0][73] ,
         \inq_ary[0][72] , \inq_ary[0][71] , \inq_ary[0][70] ,
         \inq_ary[0][69] , \inq_ary[0][68] , \inq_ary[0][67] ,
         \inq_ary[0][66] , \inq_ary[0][65] , \inq_ary[0][64] ,
         \inq_ary[0][63] , \inq_ary[0][62] , \inq_ary[0][61] ,
         \inq_ary[0][60] , \inq_ary[0][59] , \inq_ary[0][58] ,
         \inq_ary[0][57] , \inq_ary[0][56] , \inq_ary[0][55] ,
         \inq_ary[0][54] , \inq_ary[0][53] , \inq_ary[0][52] ,
         \inq_ary[0][51] , \inq_ary[0][50] , \inq_ary[0][49] ,
         \inq_ary[0][48] , \inq_ary[0][47] , \inq_ary[0][46] ,
         \inq_ary[0][45] , \inq_ary[0][44] , \inq_ary[0][43] ,
         \inq_ary[0][42] , \inq_ary[0][41] , \inq_ary[0][40] ,
         \inq_ary[0][39] , \inq_ary[0][38] , \inq_ary[0][37] ,
         \inq_ary[0][36] , \inq_ary[0][35] , \inq_ary[0][34] ,
         \inq_ary[0][33] , \inq_ary[0][32] , \inq_ary[0][31] ,
         \inq_ary[0][30] , \inq_ary[0][29] , \inq_ary[0][28] ,
         \inq_ary[0][27] , \inq_ary[0][26] , \inq_ary[0][25] ,
         \inq_ary[0][24] , \inq_ary[0][23] , \inq_ary[0][22] ,
         \inq_ary[0][21] , \inq_ary[0][20] , \inq_ary[0][19] ,
         \inq_ary[0][18] , \inq_ary[0][17] , \inq_ary[0][16] ,
         \inq_ary[0][15] , \inq_ary[0][14] , \inq_ary[0][13] ,
         \inq_ary[0][12] , \inq_ary[0][11] , \inq_ary[0][10] , \inq_ary[0][9] ,
         \inq_ary[0][8] , \inq_ary[0][7] , \inq_ary[0][6] , \inq_ary[0][5] ,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, net24660, n3574, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492;
  wire   [159:0] wrdata_d1;
  wire   [3:0] wrptr_d1;
  wire   [3:0] rdptr_d1;
  assign so_r = 1'b0;
  assign so_w = 1'b0;

  SNPS_CLOCK_GATE_HIGH_bw_r_rf16x160_0 clk_gate_byte_wen_d1_reg ( .CLK(wr_clk), 
        .EN(n3574), .ENCLK(net24660), .TE(1'b0) );
  DFFX1_RVT \wrdata_d1_reg[159]  ( .D(din[159]), .CLK(net24660), .Q(
        wrdata_d1[159]) );
  DFFX1_RVT \wrdata_d1_reg[158]  ( .D(din[158]), .CLK(net24660), .Q(
        wrdata_d1[158]) );
  DFFX1_RVT \wrdata_d1_reg[157]  ( .D(din[157]), .CLK(net24660), .Q(
        wrdata_d1[157]) );
  DFFX1_RVT \wrdata_d1_reg[156]  ( .D(din[156]), .CLK(net24660), .Q(
        wrdata_d1[156]) );
  DFFX1_RVT \wrdata_d1_reg[155]  ( .D(din[155]), .CLK(net24660), .Q(
        wrdata_d1[155]) );
  DFFX1_RVT \wrdata_d1_reg[154]  ( .D(din[154]), .CLK(net24660), .Q(
        wrdata_d1[154]) );
  DFFX1_RVT \wrdata_d1_reg[153]  ( .D(din[153]), .CLK(net24660), .Q(
        wrdata_d1[153]) );
  DFFX1_RVT \wrdata_d1_reg[152]  ( .D(din[152]), .CLK(net24660), .Q(
        wrdata_d1[152]) );
  DFFX1_RVT \wrdata_d1_reg[151]  ( .D(din[151]), .CLK(net24660), .Q(
        wrdata_d1[151]) );
  DFFX1_RVT \wrdata_d1_reg[150]  ( .D(din[150]), .CLK(net24660), .Q(
        wrdata_d1[150]) );
  DFFX1_RVT \wrdata_d1_reg[149]  ( .D(din[149]), .CLK(net24660), .Q(
        wrdata_d1[149]) );
  DFFX1_RVT \wrdata_d1_reg[148]  ( .D(din[148]), .CLK(net24660), .Q(
        wrdata_d1[148]) );
  DFFX1_RVT \wrdata_d1_reg[147]  ( .D(din[147]), .CLK(net24660), .Q(
        wrdata_d1[147]) );
  DFFX1_RVT \wrdata_d1_reg[146]  ( .D(din[146]), .CLK(net24660), .Q(
        wrdata_d1[146]) );
  DFFX1_RVT \wrdata_d1_reg[145]  ( .D(din[145]), .CLK(net24660), .Q(
        wrdata_d1[145]) );
  DFFX1_RVT \wrdata_d1_reg[144]  ( .D(din[144]), .CLK(net24660), .Q(
        wrdata_d1[144]) );
  DFFX1_RVT \wrdata_d1_reg[143]  ( .D(din[143]), .CLK(net24660), .Q(
        wrdata_d1[143]) );
  DFFX1_RVT \wrdata_d1_reg[142]  ( .D(din[142]), .CLK(net24660), .Q(
        wrdata_d1[142]) );
  DFFX1_RVT \wrdata_d1_reg[141]  ( .D(din[141]), .CLK(net24660), .Q(
        wrdata_d1[141]) );
  DFFX1_RVT \wrdata_d1_reg[140]  ( .D(din[140]), .CLK(net24660), .Q(
        wrdata_d1[140]) );
  DFFX1_RVT \wrdata_d1_reg[139]  ( .D(din[139]), .CLK(net24660), .Q(
        wrdata_d1[139]) );
  DFFX1_RVT \wrdata_d1_reg[138]  ( .D(din[138]), .CLK(net24660), .Q(
        wrdata_d1[138]) );
  DFFX1_RVT \wrdata_d1_reg[137]  ( .D(din[137]), .CLK(net24660), .Q(
        wrdata_d1[137]) );
  DFFX1_RVT \wrdata_d1_reg[136]  ( .D(din[136]), .CLK(net24660), .Q(
        wrdata_d1[136]) );
  DFFX1_RVT \wrdata_d1_reg[135]  ( .D(din[135]), .CLK(net24660), .Q(
        wrdata_d1[135]) );
  DFFX1_RVT \wrdata_d1_reg[134]  ( .D(din[134]), .CLK(net24660), .Q(
        wrdata_d1[134]) );
  DFFX1_RVT \wrdata_d1_reg[133]  ( .D(din[133]), .CLK(net24660), .Q(
        wrdata_d1[133]) );
  DFFX1_RVT \wrdata_d1_reg[132]  ( .D(din[132]), .CLK(net24660), .Q(
        wrdata_d1[132]) );
  DFFX1_RVT \wrdata_d1_reg[131]  ( .D(din[131]), .CLK(net24660), .Q(
        wrdata_d1[131]) );
  DFFX1_RVT \wrdata_d1_reg[130]  ( .D(din[130]), .CLK(net24660), .Q(
        wrdata_d1[130]) );
  DFFX1_RVT \wrdata_d1_reg[129]  ( .D(din[129]), .CLK(net24660), .Q(
        wrdata_d1[129]) );
  DFFX1_RVT \wrdata_d1_reg[128]  ( .D(din[128]), .CLK(net24660), .Q(
        wrdata_d1[128]) );
  DFFX1_RVT \wrdata_d1_reg[127]  ( .D(din[127]), .CLK(net24660), .Q(
        wrdata_d1[127]) );
  DFFX1_RVT \wrdata_d1_reg[126]  ( .D(din[126]), .CLK(net24660), .Q(
        wrdata_d1[126]) );
  DFFX1_RVT \wrdata_d1_reg[125]  ( .D(din[125]), .CLK(net24660), .Q(
        wrdata_d1[125]) );
  DFFX1_RVT \wrdata_d1_reg[124]  ( .D(din[124]), .CLK(net24660), .Q(
        wrdata_d1[124]) );
  DFFX1_RVT \wrdata_d1_reg[123]  ( .D(din[123]), .CLK(net24660), .Q(
        wrdata_d1[123]) );
  DFFX1_RVT \wrdata_d1_reg[122]  ( .D(din[122]), .CLK(net24660), .Q(
        wrdata_d1[122]) );
  DFFX1_RVT \wrdata_d1_reg[121]  ( .D(din[121]), .CLK(net24660), .Q(
        wrdata_d1[121]) );
  DFFX1_RVT \wrdata_d1_reg[120]  ( .D(din[120]), .CLK(net24660), .Q(
        wrdata_d1[120]) );
  DFFX1_RVT \wrdata_d1_reg[119]  ( .D(din[119]), .CLK(net24660), .Q(
        wrdata_d1[119]) );
  DFFX1_RVT \wrdata_d1_reg[118]  ( .D(din[118]), .CLK(net24660), .Q(
        wrdata_d1[118]) );
  DFFX1_RVT \wrdata_d1_reg[117]  ( .D(din[117]), .CLK(net24660), .Q(
        wrdata_d1[117]) );
  DFFX1_RVT \wrdata_d1_reg[116]  ( .D(din[116]), .CLK(net24660), .Q(
        wrdata_d1[116]) );
  DFFX1_RVT \wrdata_d1_reg[115]  ( .D(din[115]), .CLK(net24660), .Q(
        wrdata_d1[115]) );
  DFFX1_RVT \wrdata_d1_reg[114]  ( .D(din[114]), .CLK(net24660), .Q(
        wrdata_d1[114]) );
  DFFX1_RVT \wrdata_d1_reg[113]  ( .D(din[113]), .CLK(net24660), .Q(
        wrdata_d1[113]) );
  DFFX1_RVT \wrdata_d1_reg[112]  ( .D(din[112]), .CLK(net24660), .Q(
        wrdata_d1[112]) );
  DFFX1_RVT \wrdata_d1_reg[111]  ( .D(din[111]), .CLK(net24660), .Q(
        wrdata_d1[111]) );
  DFFX1_RVT \wrdata_d1_reg[110]  ( .D(din[110]), .CLK(net24660), .Q(
        wrdata_d1[110]) );
  DFFX1_RVT \wrdata_d1_reg[109]  ( .D(din[109]), .CLK(net24660), .Q(
        wrdata_d1[109]) );
  DFFX1_RVT \wrdata_d1_reg[108]  ( .D(din[108]), .CLK(net24660), .Q(
        wrdata_d1[108]) );
  DFFX1_RVT \wrdata_d1_reg[107]  ( .D(din[107]), .CLK(net24660), .Q(
        wrdata_d1[107]) );
  DFFX1_RVT \wrdata_d1_reg[106]  ( .D(din[106]), .CLK(net24660), .Q(
        wrdata_d1[106]) );
  DFFX1_RVT \wrdata_d1_reg[105]  ( .D(din[105]), .CLK(net24660), .Q(
        wrdata_d1[105]) );
  DFFX1_RVT \wrdata_d1_reg[104]  ( .D(din[104]), .CLK(net24660), .Q(
        wrdata_d1[104]) );
  DFFX1_RVT \wrdata_d1_reg[103]  ( .D(din[103]), .CLK(net24660), .Q(
        wrdata_d1[103]) );
  DFFX1_RVT \wrdata_d1_reg[102]  ( .D(din[102]), .CLK(net24660), .Q(
        wrdata_d1[102]) );
  DFFX1_RVT \wrdata_d1_reg[101]  ( .D(din[101]), .CLK(net24660), .Q(
        wrdata_d1[101]) );
  DFFX1_RVT \wrdata_d1_reg[100]  ( .D(din[100]), .CLK(net24660), .Q(
        wrdata_d1[100]) );
  DFFX1_RVT \wrdata_d1_reg[99]  ( .D(din[99]), .CLK(net24660), .Q(
        wrdata_d1[99]) );
  DFFX1_RVT \wrdata_d1_reg[98]  ( .D(din[98]), .CLK(net24660), .Q(
        wrdata_d1[98]) );
  DFFX1_RVT \wrdata_d1_reg[97]  ( .D(din[97]), .CLK(net24660), .Q(
        wrdata_d1[97]) );
  DFFX1_RVT \wrdata_d1_reg[96]  ( .D(din[96]), .CLK(net24660), .Q(
        wrdata_d1[96]) );
  DFFX1_RVT \wrdata_d1_reg[95]  ( .D(din[95]), .CLK(net24660), .Q(
        wrdata_d1[95]) );
  DFFX1_RVT \wrdata_d1_reg[94]  ( .D(din[94]), .CLK(net24660), .Q(
        wrdata_d1[94]) );
  DFFX1_RVT \wrdata_d1_reg[93]  ( .D(din[93]), .CLK(net24660), .Q(
        wrdata_d1[93]) );
  DFFX1_RVT \wrdata_d1_reg[92]  ( .D(din[92]), .CLK(net24660), .Q(
        wrdata_d1[92]) );
  DFFX1_RVT \wrdata_d1_reg[91]  ( .D(din[91]), .CLK(net24660), .Q(
        wrdata_d1[91]) );
  DFFX1_RVT \wrdata_d1_reg[90]  ( .D(din[90]), .CLK(net24660), .Q(
        wrdata_d1[90]) );
  DFFX1_RVT \wrdata_d1_reg[89]  ( .D(din[89]), .CLK(net24660), .Q(
        wrdata_d1[89]) );
  DFFX1_RVT \wrdata_d1_reg[88]  ( .D(din[88]), .CLK(net24660), .Q(
        wrdata_d1[88]) );
  DFFX1_RVT \wrdata_d1_reg[87]  ( .D(din[87]), .CLK(net24660), .Q(
        wrdata_d1[87]) );
  DFFX1_RVT \wrdata_d1_reg[86]  ( .D(din[86]), .CLK(net24660), .Q(
        wrdata_d1[86]) );
  DFFX1_RVT \wrdata_d1_reg[85]  ( .D(din[85]), .CLK(net24660), .Q(
        wrdata_d1[85]) );
  DFFX1_RVT \wrdata_d1_reg[84]  ( .D(din[84]), .CLK(net24660), .Q(
        wrdata_d1[84]) );
  DFFX1_RVT \wrdata_d1_reg[83]  ( .D(din[83]), .CLK(net24660), .Q(
        wrdata_d1[83]) );
  DFFX1_RVT \wrdata_d1_reg[82]  ( .D(din[82]), .CLK(net24660), .Q(
        wrdata_d1[82]) );
  DFFX1_RVT \wrdata_d1_reg[81]  ( .D(din[81]), .CLK(net24660), .Q(
        wrdata_d1[81]) );
  DFFX1_RVT \wrdata_d1_reg[80]  ( .D(din[80]), .CLK(net24660), .Q(
        wrdata_d1[80]) );
  DFFX1_RVT \wrdata_d1_reg[79]  ( .D(din[79]), .CLK(net24660), .Q(
        wrdata_d1[79]) );
  DFFX1_RVT \wrdata_d1_reg[78]  ( .D(din[78]), .CLK(net24660), .Q(
        wrdata_d1[78]) );
  DFFX1_RVT \wrdata_d1_reg[77]  ( .D(din[77]), .CLK(net24660), .Q(
        wrdata_d1[77]) );
  DFFX1_RVT \wrdata_d1_reg[76]  ( .D(din[76]), .CLK(net24660), .Q(
        wrdata_d1[76]) );
  DFFX1_RVT \wrdata_d1_reg[75]  ( .D(din[75]), .CLK(net24660), .Q(
        wrdata_d1[75]) );
  DFFX1_RVT \wrdata_d1_reg[74]  ( .D(din[74]), .CLK(net24660), .Q(
        wrdata_d1[74]) );
  DFFX1_RVT \wrdata_d1_reg[73]  ( .D(din[73]), .CLK(net24660), .Q(
        wrdata_d1[73]) );
  DFFX1_RVT \wrdata_d1_reg[72]  ( .D(din[72]), .CLK(net24660), .Q(
        wrdata_d1[72]) );
  DFFX1_RVT \wrdata_d1_reg[71]  ( .D(din[71]), .CLK(net24660), .Q(
        wrdata_d1[71]) );
  DFFX1_RVT \wrdata_d1_reg[70]  ( .D(din[70]), .CLK(net24660), .Q(
        wrdata_d1[70]) );
  DFFX1_RVT \wrdata_d1_reg[69]  ( .D(din[69]), .CLK(net24660), .Q(
        wrdata_d1[69]) );
  DFFX1_RVT \wrdata_d1_reg[68]  ( .D(din[68]), .CLK(net24660), .Q(
        wrdata_d1[68]) );
  DFFX1_RVT \wrdata_d1_reg[67]  ( .D(din[67]), .CLK(net24660), .Q(
        wrdata_d1[67]) );
  DFFX1_RVT \wrdata_d1_reg[66]  ( .D(din[66]), .CLK(net24660), .Q(
        wrdata_d1[66]) );
  DFFX1_RVT \wrdata_d1_reg[65]  ( .D(din[65]), .CLK(net24660), .Q(
        wrdata_d1[65]) );
  DFFX1_RVT \wrdata_d1_reg[64]  ( .D(din[64]), .CLK(net24660), .Q(
        wrdata_d1[64]) );
  DFFX1_RVT \wrdata_d1_reg[63]  ( .D(din[63]), .CLK(net24660), .Q(
        wrdata_d1[63]) );
  DFFX1_RVT \wrdata_d1_reg[62]  ( .D(din[62]), .CLK(net24660), .Q(
        wrdata_d1[62]) );
  DFFX1_RVT \wrdata_d1_reg[61]  ( .D(din[61]), .CLK(net24660), .Q(
        wrdata_d1[61]) );
  DFFX1_RVT \wrdata_d1_reg[60]  ( .D(din[60]), .CLK(net24660), .Q(
        wrdata_d1[60]) );
  DFFX1_RVT \wrdata_d1_reg[59]  ( .D(din[59]), .CLK(net24660), .Q(
        wrdata_d1[59]) );
  DFFX1_RVT \wrdata_d1_reg[58]  ( .D(din[58]), .CLK(net24660), .Q(
        wrdata_d1[58]) );
  DFFX1_RVT \wrdata_d1_reg[57]  ( .D(din[57]), .CLK(net24660), .Q(
        wrdata_d1[57]) );
  DFFX1_RVT \wrdata_d1_reg[56]  ( .D(din[56]), .CLK(net24660), .Q(
        wrdata_d1[56]) );
  DFFX1_RVT \wrdata_d1_reg[55]  ( .D(din[55]), .CLK(net24660), .Q(
        wrdata_d1[55]) );
  DFFX1_RVT \wrdata_d1_reg[54]  ( .D(din[54]), .CLK(net24660), .Q(
        wrdata_d1[54]) );
  DFFX1_RVT \wrdata_d1_reg[53]  ( .D(din[53]), .CLK(net24660), .Q(
        wrdata_d1[53]) );
  DFFX1_RVT \wrdata_d1_reg[52]  ( .D(din[52]), .CLK(net24660), .Q(
        wrdata_d1[52]) );
  DFFX1_RVT \wrdata_d1_reg[51]  ( .D(din[51]), .CLK(net24660), .Q(
        wrdata_d1[51]) );
  DFFX1_RVT \wrdata_d1_reg[50]  ( .D(din[50]), .CLK(net24660), .Q(
        wrdata_d1[50]) );
  DFFX1_RVT \wrdata_d1_reg[49]  ( .D(din[49]), .CLK(net24660), .Q(
        wrdata_d1[49]) );
  DFFX1_RVT \wrdata_d1_reg[48]  ( .D(din[48]), .CLK(net24660), .Q(
        wrdata_d1[48]) );
  DFFX1_RVT \wrdata_d1_reg[47]  ( .D(din[47]), .CLK(net24660), .Q(
        wrdata_d1[47]) );
  DFFX1_RVT \wrdata_d1_reg[46]  ( .D(din[46]), .CLK(net24660), .Q(
        wrdata_d1[46]) );
  DFFX1_RVT \wrdata_d1_reg[45]  ( .D(din[45]), .CLK(net24660), .Q(
        wrdata_d1[45]) );
  DFFX1_RVT \wrdata_d1_reg[44]  ( .D(din[44]), .CLK(net24660), .Q(
        wrdata_d1[44]) );
  DFFX1_RVT \wrdata_d1_reg[43]  ( .D(din[43]), .CLK(net24660), .Q(
        wrdata_d1[43]) );
  DFFX1_RVT \wrdata_d1_reg[42]  ( .D(din[42]), .CLK(net24660), .Q(
        wrdata_d1[42]) );
  DFFX1_RVT \wrdata_d1_reg[41]  ( .D(din[41]), .CLK(net24660), .Q(
        wrdata_d1[41]) );
  DFFX1_RVT \wrdata_d1_reg[40]  ( .D(din[40]), .CLK(net24660), .Q(
        wrdata_d1[40]) );
  DFFX1_RVT \wrdata_d1_reg[39]  ( .D(din[39]), .CLK(net24660), .Q(
        wrdata_d1[39]) );
  DFFX1_RVT \wrdata_d1_reg[38]  ( .D(din[38]), .CLK(net24660), .Q(
        wrdata_d1[38]) );
  DFFX1_RVT \wrdata_d1_reg[37]  ( .D(din[37]), .CLK(net24660), .Q(
        wrdata_d1[37]) );
  DFFX1_RVT \wrdata_d1_reg[36]  ( .D(din[36]), .CLK(net24660), .Q(
        wrdata_d1[36]) );
  DFFX1_RVT \wrdata_d1_reg[35]  ( .D(din[35]), .CLK(net24660), .Q(
        wrdata_d1[35]) );
  DFFX1_RVT \wrdata_d1_reg[34]  ( .D(din[34]), .CLK(net24660), .Q(
        wrdata_d1[34]) );
  DFFX1_RVT \wrdata_d1_reg[33]  ( .D(din[33]), .CLK(net24660), .Q(
        wrdata_d1[33]) );
  DFFX1_RVT \wrdata_d1_reg[32]  ( .D(din[32]), .CLK(net24660), .Q(
        wrdata_d1[32]) );
  DFFX1_RVT \wrdata_d1_reg[31]  ( .D(din[31]), .CLK(net24660), .Q(
        wrdata_d1[31]) );
  DFFX1_RVT \wrdata_d1_reg[30]  ( .D(din[30]), .CLK(net24660), .Q(
        wrdata_d1[30]) );
  DFFX1_RVT \wrdata_d1_reg[29]  ( .D(din[29]), .CLK(net24660), .Q(
        wrdata_d1[29]) );
  DFFX1_RVT \wrdata_d1_reg[28]  ( .D(din[28]), .CLK(net24660), .Q(
        wrdata_d1[28]) );
  DFFX1_RVT \wrdata_d1_reg[27]  ( .D(din[27]), .CLK(net24660), .Q(
        wrdata_d1[27]) );
  DFFX1_RVT \wrdata_d1_reg[26]  ( .D(din[26]), .CLK(net24660), .Q(
        wrdata_d1[26]) );
  DFFX1_RVT \wrdata_d1_reg[25]  ( .D(din[25]), .CLK(net24660), .Q(
        wrdata_d1[25]) );
  DFFX1_RVT \wrdata_d1_reg[24]  ( .D(din[24]), .CLK(net24660), .Q(
        wrdata_d1[24]) );
  DFFX1_RVT \wrdata_d1_reg[23]  ( .D(din[23]), .CLK(net24660), .Q(
        wrdata_d1[23]) );
  DFFX1_RVT \wrdata_d1_reg[22]  ( .D(din[22]), .CLK(net24660), .Q(
        wrdata_d1[22]) );
  DFFX1_RVT \wrdata_d1_reg[21]  ( .D(din[21]), .CLK(net24660), .Q(
        wrdata_d1[21]) );
  DFFX1_RVT \wrdata_d1_reg[20]  ( .D(din[20]), .CLK(net24660), .Q(
        wrdata_d1[20]) );
  DFFX1_RVT \wrdata_d1_reg[19]  ( .D(din[19]), .CLK(net24660), .Q(
        wrdata_d1[19]) );
  DFFX1_RVT \wrdata_d1_reg[18]  ( .D(din[18]), .CLK(net24660), .Q(
        wrdata_d1[18]) );
  DFFX1_RVT \wrdata_d1_reg[17]  ( .D(din[17]), .CLK(net24660), .Q(
        wrdata_d1[17]) );
  DFFX1_RVT \wrdata_d1_reg[16]  ( .D(din[16]), .CLK(net24660), .Q(
        wrdata_d1[16]) );
  DFFX1_RVT \wrdata_d1_reg[15]  ( .D(din[15]), .CLK(net24660), .Q(
        wrdata_d1[15]) );
  DFFX1_RVT \wrdata_d1_reg[14]  ( .D(din[14]), .CLK(net24660), .Q(
        wrdata_d1[14]) );
  DFFX1_RVT \wrdata_d1_reg[13]  ( .D(din[13]), .CLK(net24660), .Q(
        wrdata_d1[13]) );
  DFFX1_RVT \wrdata_d1_reg[12]  ( .D(din[12]), .CLK(net24660), .Q(
        wrdata_d1[12]) );
  DFFX1_RVT \wrdata_d1_reg[11]  ( .D(din[11]), .CLK(net24660), .Q(
        wrdata_d1[11]) );
  DFFX1_RVT \wrdata_d1_reg[10]  ( .D(din[10]), .CLK(net24660), .Q(
        wrdata_d1[10]) );
  DFFX1_RVT \wrdata_d1_reg[9]  ( .D(din[9]), .CLK(net24660), .Q(wrdata_d1[9])
         );
  DFFX1_RVT \wrdata_d1_reg[8]  ( .D(din[8]), .CLK(net24660), .Q(wrdata_d1[8])
         );
  DFFX1_RVT \wrdata_d1_reg[7]  ( .D(din[7]), .CLK(net24660), .Q(wrdata_d1[7])
         );
  DFFX1_RVT \wrdata_d1_reg[6]  ( .D(din[6]), .CLK(net24660), .Q(wrdata_d1[6])
         );
  DFFX1_RVT \wrdata_d1_reg[5]  ( .D(din[5]), .CLK(net24660), .Q(wrdata_d1[5])
         );
  DFFX1_RVT wr_en_d1_reg ( .D(wr_en), .CLK(net24660), .Q(wr_en_d1) );
  DFFX1_RVT \rdptr_d1_reg[2]  ( .D(rd_adr[2]), .CLK(net24660), .Q(rdptr_d1[2]), 
        .QN(n3338) );
  LATCHX1_RVT \inq_ary_reg[0][159]  ( .CLK(n3491), .D(n1761), .Q(
        \inq_ary[0][159] ) );
  LATCHX1_RVT \inq_ary_reg[1][159]  ( .CLK(n3490), .D(n1761), .Q(
        \inq_ary[1][159] ) );
  LATCHX1_RVT \inq_ary_reg[2][159]  ( .CLK(n3489), .D(n1761), .Q(
        \inq_ary[2][159] ) );
  LATCHX1_RVT \inq_ary_reg[3][159]  ( .CLK(n3488), .D(n1761), .Q(
        \inq_ary[3][159] ) );
  LATCHX1_RVT \inq_ary_reg[4][159]  ( .CLK(n3487), .D(n1761), .Q(
        \inq_ary[4][159] ) );
  LATCHX1_RVT \inq_ary_reg[5][159]  ( .CLK(n3486), .D(n1761), .Q(
        \inq_ary[5][159] ) );
  LATCHX1_RVT \inq_ary_reg[6][159]  ( .CLK(n3485), .D(n1761), .Q(
        \inq_ary[6][159] ) );
  LATCHX1_RVT \inq_ary_reg[7][159]  ( .CLK(n3484), .D(n1761), .Q(
        \inq_ary[7][159] ) );
  LATCHX1_RVT \inq_ary_reg[8][159]  ( .CLK(n3483), .D(n1761), .Q(
        \inq_ary[8][159] ) );
  LATCHX1_RVT \inq_ary_reg[9][159]  ( .CLK(n3482), .D(n1761), .Q(
        \inq_ary[9][159] ) );
  LATCHX1_RVT \inq_ary_reg[10][159]  ( .CLK(n3481), .D(n1761), .Q(
        \inq_ary[10][159] ) );
  LATCHX1_RVT \inq_ary_reg[11][159]  ( .CLK(n3480), .D(n1761), .Q(
        \inq_ary[11][159] ) );
  LATCHX1_RVT \inq_ary_reg[12][159]  ( .CLK(n3479), .D(n1761), .Q(
        \inq_ary[12][159] ) );
  LATCHX1_RVT \inq_ary_reg[13][159]  ( .CLK(n3478), .D(n1761), .Q(
        \inq_ary[13][159] ) );
  LATCHX1_RVT \inq_ary_reg[14][159]  ( .CLK(n3477), .D(n1761), .Q(
        \inq_ary[14][159] ) );
  LATCHX1_RVT \inq_ary_reg[15][159]  ( .CLK(n3476), .D(n1761), .Q(
        \inq_ary[15][159] ) );
  LATCHX1_RVT \dout_reg[159]  ( .CLK(n3492), .D(N421), .Q(dout[159]) );
  LATCHX1_RVT \inq_ary_reg[0][158]  ( .CLK(n3491), .D(n1660), .Q(
        \inq_ary[0][158] ) );
  LATCHX1_RVT \inq_ary_reg[1][158]  ( .CLK(n3490), .D(n1660), .Q(
        \inq_ary[1][158] ) );
  LATCHX1_RVT \inq_ary_reg[2][158]  ( .CLK(n3489), .D(n1660), .Q(
        \inq_ary[2][158] ) );
  LATCHX1_RVT \inq_ary_reg[3][158]  ( .CLK(n3488), .D(n1660), .Q(
        \inq_ary[3][158] ) );
  LATCHX1_RVT \inq_ary_reg[4][158]  ( .CLK(n3487), .D(n1660), .Q(
        \inq_ary[4][158] ) );
  LATCHX1_RVT \inq_ary_reg[5][158]  ( .CLK(n3486), .D(n1660), .Q(
        \inq_ary[5][158] ) );
  LATCHX1_RVT \inq_ary_reg[6][158]  ( .CLK(n3485), .D(n1660), .Q(
        \inq_ary[6][158] ) );
  LATCHX1_RVT \inq_ary_reg[7][158]  ( .CLK(n3484), .D(n1660), .Q(
        \inq_ary[7][158] ) );
  LATCHX1_RVT \inq_ary_reg[8][158]  ( .CLK(n3483), .D(n1660), .Q(
        \inq_ary[8][158] ) );
  LATCHX1_RVT \inq_ary_reg[9][158]  ( .CLK(n3482), .D(n1660), .Q(
        \inq_ary[9][158] ) );
  LATCHX1_RVT \inq_ary_reg[10][158]  ( .CLK(n3481), .D(n1660), .Q(
        \inq_ary[10][158] ) );
  LATCHX1_RVT \inq_ary_reg[11][158]  ( .CLK(n3480), .D(n1660), .Q(
        \inq_ary[11][158] ) );
  LATCHX1_RVT \inq_ary_reg[12][158]  ( .CLK(n3479), .D(n1660), .Q(
        \inq_ary[12][158] ) );
  LATCHX1_RVT \inq_ary_reg[13][158]  ( .CLK(n3478), .D(n1660), .Q(
        \inq_ary[13][158] ) );
  LATCHX1_RVT \inq_ary_reg[14][158]  ( .CLK(n3477), .D(n1660), .Q(
        \inq_ary[14][158] ) );
  LATCHX1_RVT \inq_ary_reg[15][158]  ( .CLK(n3476), .D(n1660), .Q(
        \inq_ary[15][158] ) );
  LATCHX1_RVT \dout_reg[158]  ( .CLK(n3492), .D(N420), .Q(dout[158]) );
  LATCHX1_RVT \inq_ary_reg[0][157]  ( .CLK(n3491), .D(n1648), .Q(
        \inq_ary[0][157] ) );
  LATCHX1_RVT \inq_ary_reg[1][157]  ( .CLK(n3490), .D(n1648), .Q(
        \inq_ary[1][157] ) );
  LATCHX1_RVT \inq_ary_reg[2][157]  ( .CLK(n3489), .D(n1648), .Q(
        \inq_ary[2][157] ) );
  LATCHX1_RVT \inq_ary_reg[3][157]  ( .CLK(n3488), .D(n1648), .Q(
        \inq_ary[3][157] ) );
  LATCHX1_RVT \inq_ary_reg[4][157]  ( .CLK(n3487), .D(n1648), .Q(
        \inq_ary[4][157] ) );
  LATCHX1_RVT \inq_ary_reg[5][157]  ( .CLK(n3486), .D(n1648), .Q(
        \inq_ary[5][157] ) );
  LATCHX1_RVT \inq_ary_reg[6][157]  ( .CLK(n3485), .D(n1648), .Q(
        \inq_ary[6][157] ) );
  LATCHX1_RVT \inq_ary_reg[7][157]  ( .CLK(n3484), .D(n1648), .Q(
        \inq_ary[7][157] ) );
  LATCHX1_RVT \inq_ary_reg[8][157]  ( .CLK(n3483), .D(n1648), .Q(
        \inq_ary[8][157] ) );
  LATCHX1_RVT \inq_ary_reg[9][157]  ( .CLK(n3482), .D(n1648), .Q(
        \inq_ary[9][157] ) );
  LATCHX1_RVT \inq_ary_reg[10][157]  ( .CLK(n3481), .D(n1648), .Q(
        \inq_ary[10][157] ) );
  LATCHX1_RVT \inq_ary_reg[11][157]  ( .CLK(n3480), .D(n1648), .Q(
        \inq_ary[11][157] ) );
  LATCHX1_RVT \inq_ary_reg[12][157]  ( .CLK(n3479), .D(n1648), .Q(
        \inq_ary[12][157] ) );
  LATCHX1_RVT \inq_ary_reg[13][157]  ( .CLK(n3478), .D(n1648), .Q(
        \inq_ary[13][157] ) );
  LATCHX1_RVT \inq_ary_reg[14][157]  ( .CLK(n3477), .D(n1648), .Q(
        \inq_ary[14][157] ) );
  LATCHX1_RVT \inq_ary_reg[15][157]  ( .CLK(n3476), .D(n1648), .Q(
        \inq_ary[15][157] ) );
  LATCHX1_RVT \dout_reg[157]  ( .CLK(n3492), .D(N419), .Q(dout[157]) );
  LATCHX1_RVT \inq_ary_reg[0][156]  ( .CLK(n3491), .D(n1636), .Q(
        \inq_ary[0][156] ) );
  LATCHX1_RVT \inq_ary_reg[1][156]  ( .CLK(n3490), .D(n1636), .Q(
        \inq_ary[1][156] ) );
  LATCHX1_RVT \inq_ary_reg[2][156]  ( .CLK(n3489), .D(n1636), .Q(
        \inq_ary[2][156] ) );
  LATCHX1_RVT \inq_ary_reg[3][156]  ( .CLK(n3488), .D(n1636), .Q(
        \inq_ary[3][156] ) );
  LATCHX1_RVT \inq_ary_reg[4][156]  ( .CLK(n3487), .D(n1636), .Q(
        \inq_ary[4][156] ) );
  LATCHX1_RVT \inq_ary_reg[5][156]  ( .CLK(n3486), .D(n1636), .Q(
        \inq_ary[5][156] ) );
  LATCHX1_RVT \inq_ary_reg[6][156]  ( .CLK(n3485), .D(n1636), .Q(
        \inq_ary[6][156] ) );
  LATCHX1_RVT \inq_ary_reg[7][156]  ( .CLK(n3484), .D(n1636), .Q(
        \inq_ary[7][156] ) );
  LATCHX1_RVT \inq_ary_reg[8][156]  ( .CLK(n3483), .D(n1636), .Q(
        \inq_ary[8][156] ) );
  LATCHX1_RVT \inq_ary_reg[9][156]  ( .CLK(n3482), .D(n1636), .Q(
        \inq_ary[9][156] ) );
  LATCHX1_RVT \inq_ary_reg[10][156]  ( .CLK(n3481), .D(n1636), .Q(
        \inq_ary[10][156] ) );
  LATCHX1_RVT \inq_ary_reg[11][156]  ( .CLK(n3480), .D(n1636), .Q(
        \inq_ary[11][156] ) );
  LATCHX1_RVT \inq_ary_reg[12][156]  ( .CLK(n3479), .D(n1636), .Q(
        \inq_ary[12][156] ) );
  LATCHX1_RVT \inq_ary_reg[13][156]  ( .CLK(n3478), .D(n1636), .Q(
        \inq_ary[13][156] ) );
  LATCHX1_RVT \inq_ary_reg[14][156]  ( .CLK(n3477), .D(n1636), .Q(
        \inq_ary[14][156] ) );
  LATCHX1_RVT \inq_ary_reg[15][156]  ( .CLK(n3476), .D(n1636), .Q(
        \inq_ary[15][156] ) );
  LATCHX1_RVT \dout_reg[156]  ( .CLK(n3492), .D(N418), .Q(dout[156]) );
  LATCHX1_RVT \inq_ary_reg[0][155]  ( .CLK(n3491), .D(n1624), .Q(
        \inq_ary[0][155] ) );
  LATCHX1_RVT \inq_ary_reg[1][155]  ( .CLK(n3490), .D(n1624), .Q(
        \inq_ary[1][155] ) );
  LATCHX1_RVT \inq_ary_reg[2][155]  ( .CLK(n3489), .D(n1624), .Q(
        \inq_ary[2][155] ) );
  LATCHX1_RVT \inq_ary_reg[3][155]  ( .CLK(n3488), .D(n1624), .Q(
        \inq_ary[3][155] ) );
  LATCHX1_RVT \inq_ary_reg[4][155]  ( .CLK(n3487), .D(n1624), .Q(
        \inq_ary[4][155] ) );
  LATCHX1_RVT \inq_ary_reg[5][155]  ( .CLK(n3486), .D(n1624), .Q(
        \inq_ary[5][155] ) );
  LATCHX1_RVT \inq_ary_reg[6][155]  ( .CLK(n3485), .D(n1624), .Q(
        \inq_ary[6][155] ) );
  LATCHX1_RVT \inq_ary_reg[7][155]  ( .CLK(n3484), .D(n1624), .Q(
        \inq_ary[7][155] ) );
  LATCHX1_RVT \inq_ary_reg[8][155]  ( .CLK(n3483), .D(n1624), .Q(
        \inq_ary[8][155] ) );
  LATCHX1_RVT \inq_ary_reg[9][155]  ( .CLK(n3482), .D(n1624), .Q(
        \inq_ary[9][155] ) );
  LATCHX1_RVT \inq_ary_reg[10][155]  ( .CLK(n3481), .D(n1624), .Q(
        \inq_ary[10][155] ) );
  LATCHX1_RVT \inq_ary_reg[11][155]  ( .CLK(n3480), .D(n1624), .Q(
        \inq_ary[11][155] ) );
  LATCHX1_RVT \inq_ary_reg[12][155]  ( .CLK(n3479), .D(n1624), .Q(
        \inq_ary[12][155] ) );
  LATCHX1_RVT \inq_ary_reg[13][155]  ( .CLK(n3478), .D(n1624), .Q(
        \inq_ary[13][155] ) );
  LATCHX1_RVT \inq_ary_reg[14][155]  ( .CLK(n3477), .D(n1624), .Q(
        \inq_ary[14][155] ) );
  LATCHX1_RVT \inq_ary_reg[15][155]  ( .CLK(n3476), .D(n1624), .Q(
        \inq_ary[15][155] ) );
  LATCHX1_RVT \dout_reg[155]  ( .CLK(n3492), .D(N417), .Q(dout[155]) );
  LATCHX1_RVT \inq_ary_reg[0][154]  ( .CLK(n3491), .D(n1611), .Q(
        \inq_ary[0][154] ) );
  LATCHX1_RVT \inq_ary_reg[1][154]  ( .CLK(n3490), .D(n1611), .Q(
        \inq_ary[1][154] ) );
  LATCHX1_RVT \inq_ary_reg[2][154]  ( .CLK(n3489), .D(n1611), .Q(
        \inq_ary[2][154] ) );
  LATCHX1_RVT \inq_ary_reg[3][154]  ( .CLK(n3488), .D(n1611), .Q(
        \inq_ary[3][154] ) );
  LATCHX1_RVT \inq_ary_reg[4][154]  ( .CLK(n3487), .D(n1611), .Q(
        \inq_ary[4][154] ) );
  LATCHX1_RVT \inq_ary_reg[5][154]  ( .CLK(n3486), .D(n1611), .Q(
        \inq_ary[5][154] ) );
  LATCHX1_RVT \inq_ary_reg[6][154]  ( .CLK(n3485), .D(n1611), .Q(
        \inq_ary[6][154] ) );
  LATCHX1_RVT \inq_ary_reg[7][154]  ( .CLK(n3484), .D(n1611), .Q(
        \inq_ary[7][154] ) );
  LATCHX1_RVT \inq_ary_reg[8][154]  ( .CLK(n3483), .D(n1611), .Q(
        \inq_ary[8][154] ) );
  LATCHX1_RVT \inq_ary_reg[9][154]  ( .CLK(n3482), .D(n1611), .Q(
        \inq_ary[9][154] ) );
  LATCHX1_RVT \inq_ary_reg[10][154]  ( .CLK(n3481), .D(n1611), .Q(
        \inq_ary[10][154] ) );
  LATCHX1_RVT \inq_ary_reg[11][154]  ( .CLK(n3480), .D(n1611), .Q(
        \inq_ary[11][154] ) );
  LATCHX1_RVT \inq_ary_reg[12][154]  ( .CLK(n3479), .D(n1611), .Q(
        \inq_ary[12][154] ) );
  LATCHX1_RVT \inq_ary_reg[13][154]  ( .CLK(n3478), .D(n1611), .Q(
        \inq_ary[13][154] ) );
  LATCHX1_RVT \inq_ary_reg[14][154]  ( .CLK(n3477), .D(n1611), .Q(
        \inq_ary[14][154] ) );
  LATCHX1_RVT \inq_ary_reg[15][154]  ( .CLK(n3476), .D(n1611), .Q(
        \inq_ary[15][154] ) );
  LATCHX1_RVT \dout_reg[154]  ( .CLK(n3492), .D(N416), .Q(dout[154]) );
  LATCHX1_RVT \inq_ary_reg[0][153]  ( .CLK(n3491), .D(n1737), .Q(
        \inq_ary[0][153] ) );
  LATCHX1_RVT \inq_ary_reg[1][153]  ( .CLK(n3490), .D(n1737), .Q(
        \inq_ary[1][153] ) );
  LATCHX1_RVT \inq_ary_reg[2][153]  ( .CLK(n3489), .D(n1737), .Q(
        \inq_ary[2][153] ) );
  LATCHX1_RVT \inq_ary_reg[3][153]  ( .CLK(n3488), .D(n1737), .Q(
        \inq_ary[3][153] ) );
  LATCHX1_RVT \inq_ary_reg[4][153]  ( .CLK(n3487), .D(n1737), .Q(
        \inq_ary[4][153] ) );
  LATCHX1_RVT \inq_ary_reg[5][153]  ( .CLK(n3486), .D(n1737), .Q(
        \inq_ary[5][153] ) );
  LATCHX1_RVT \inq_ary_reg[6][153]  ( .CLK(n3485), .D(n1737), .Q(
        \inq_ary[6][153] ) );
  LATCHX1_RVT \inq_ary_reg[7][153]  ( .CLK(n3484), .D(n1737), .Q(
        \inq_ary[7][153] ) );
  LATCHX1_RVT \inq_ary_reg[8][153]  ( .CLK(n3483), .D(n1737), .Q(
        \inq_ary[8][153] ) );
  LATCHX1_RVT \inq_ary_reg[9][153]  ( .CLK(n3482), .D(n1737), .Q(
        \inq_ary[9][153] ) );
  LATCHX1_RVT \inq_ary_reg[10][153]  ( .CLK(n3481), .D(n1737), .Q(
        \inq_ary[10][153] ) );
  LATCHX1_RVT \inq_ary_reg[11][153]  ( .CLK(n3480), .D(n1737), .Q(
        \inq_ary[11][153] ) );
  LATCHX1_RVT \inq_ary_reg[12][153]  ( .CLK(n3479), .D(n1737), .Q(
        \inq_ary[12][153] ) );
  LATCHX1_RVT \inq_ary_reg[13][153]  ( .CLK(n3478), .D(n1737), .Q(
        \inq_ary[13][153] ) );
  LATCHX1_RVT \inq_ary_reg[14][153]  ( .CLK(n3477), .D(n1737), .Q(
        \inq_ary[14][153] ) );
  LATCHX1_RVT \inq_ary_reg[15][153]  ( .CLK(n3476), .D(n1737), .Q(
        \inq_ary[15][153] ) );
  LATCHX1_RVT \dout_reg[153]  ( .CLK(n3492), .D(N415), .Q(dout[153]) );
  LATCHX1_RVT \inq_ary_reg[0][152]  ( .CLK(n3491), .D(n1724), .Q(
        \inq_ary[0][152] ) );
  LATCHX1_RVT \inq_ary_reg[1][152]  ( .CLK(n3490), .D(n1724), .Q(
        \inq_ary[1][152] ) );
  LATCHX1_RVT \inq_ary_reg[2][152]  ( .CLK(n3489), .D(n1724), .Q(
        \inq_ary[2][152] ) );
  LATCHX1_RVT \inq_ary_reg[3][152]  ( .CLK(n3488), .D(n1724), .Q(
        \inq_ary[3][152] ) );
  LATCHX1_RVT \inq_ary_reg[4][152]  ( .CLK(n3487), .D(n1724), .Q(
        \inq_ary[4][152] ) );
  LATCHX1_RVT \inq_ary_reg[5][152]  ( .CLK(n3486), .D(n1724), .Q(
        \inq_ary[5][152] ) );
  LATCHX1_RVT \inq_ary_reg[6][152]  ( .CLK(n3485), .D(n1724), .Q(
        \inq_ary[6][152] ) );
  LATCHX1_RVT \inq_ary_reg[7][152]  ( .CLK(n3484), .D(n1724), .Q(
        \inq_ary[7][152] ) );
  LATCHX1_RVT \inq_ary_reg[8][152]  ( .CLK(n3483), .D(n1724), .Q(
        \inq_ary[8][152] ) );
  LATCHX1_RVT \inq_ary_reg[9][152]  ( .CLK(n3482), .D(n1724), .Q(
        \inq_ary[9][152] ) );
  LATCHX1_RVT \inq_ary_reg[10][152]  ( .CLK(n3481), .D(n1724), .Q(
        \inq_ary[10][152] ) );
  LATCHX1_RVT \inq_ary_reg[11][152]  ( .CLK(n3480), .D(n1724), .Q(
        \inq_ary[11][152] ) );
  LATCHX1_RVT \inq_ary_reg[12][152]  ( .CLK(n3479), .D(n1724), .Q(
        \inq_ary[12][152] ) );
  LATCHX1_RVT \inq_ary_reg[13][152]  ( .CLK(n3478), .D(n1724), .Q(
        \inq_ary[13][152] ) );
  LATCHX1_RVT \inq_ary_reg[14][152]  ( .CLK(n3477), .D(n1724), .Q(
        \inq_ary[14][152] ) );
  LATCHX1_RVT \inq_ary_reg[15][152]  ( .CLK(n3476), .D(n1724), .Q(
        \inq_ary[15][152] ) );
  LATCHX1_RVT \dout_reg[152]  ( .CLK(n3492), .D(N414), .Q(dout[152]) );
  LATCHX1_RVT \inq_ary_reg[0][151]  ( .CLK(n3491), .D(n1710), .Q(
        \inq_ary[0][151] ) );
  LATCHX1_RVT \inq_ary_reg[1][151]  ( .CLK(n3490), .D(n1710), .Q(
        \inq_ary[1][151] ) );
  LATCHX1_RVT \inq_ary_reg[2][151]  ( .CLK(n3489), .D(n1710), .Q(
        \inq_ary[2][151] ) );
  LATCHX1_RVT \inq_ary_reg[3][151]  ( .CLK(n3488), .D(n1710), .Q(
        \inq_ary[3][151] ) );
  LATCHX1_RVT \inq_ary_reg[4][151]  ( .CLK(n3487), .D(n1710), .Q(
        \inq_ary[4][151] ) );
  LATCHX1_RVT \inq_ary_reg[5][151]  ( .CLK(n3486), .D(n1710), .Q(
        \inq_ary[5][151] ) );
  LATCHX1_RVT \inq_ary_reg[6][151]  ( .CLK(n3485), .D(n1710), .Q(
        \inq_ary[6][151] ) );
  LATCHX1_RVT \inq_ary_reg[7][151]  ( .CLK(n3484), .D(n1710), .Q(
        \inq_ary[7][151] ) );
  LATCHX1_RVT \inq_ary_reg[8][151]  ( .CLK(n3483), .D(n1710), .Q(
        \inq_ary[8][151] ) );
  LATCHX1_RVT \inq_ary_reg[9][151]  ( .CLK(n3482), .D(n1710), .Q(
        \inq_ary[9][151] ) );
  LATCHX1_RVT \inq_ary_reg[10][151]  ( .CLK(n3481), .D(n1710), .Q(
        \inq_ary[10][151] ) );
  LATCHX1_RVT \inq_ary_reg[11][151]  ( .CLK(n3480), .D(n1710), .Q(
        \inq_ary[11][151] ) );
  LATCHX1_RVT \inq_ary_reg[12][151]  ( .CLK(n3479), .D(n1710), .Q(
        \inq_ary[12][151] ) );
  LATCHX1_RVT \inq_ary_reg[13][151]  ( .CLK(n3478), .D(n1710), .Q(
        \inq_ary[13][151] ) );
  LATCHX1_RVT \inq_ary_reg[14][151]  ( .CLK(n3477), .D(n1710), .Q(
        \inq_ary[14][151] ) );
  LATCHX1_RVT \inq_ary_reg[15][151]  ( .CLK(n3476), .D(n1710), .Q(
        \inq_ary[15][151] ) );
  LATCHX1_RVT \dout_reg[151]  ( .CLK(n3492), .D(N413), .Q(dout[151]) );
  LATCHX1_RVT \inq_ary_reg[0][150]  ( .CLK(n3491), .D(n1698), .Q(
        \inq_ary[0][150] ) );
  LATCHX1_RVT \inq_ary_reg[1][150]  ( .CLK(n3490), .D(n1698), .Q(
        \inq_ary[1][150] ) );
  LATCHX1_RVT \inq_ary_reg[2][150]  ( .CLK(n3489), .D(n1698), .Q(
        \inq_ary[2][150] ) );
  LATCHX1_RVT \inq_ary_reg[3][150]  ( .CLK(n3488), .D(n1698), .Q(
        \inq_ary[3][150] ) );
  LATCHX1_RVT \inq_ary_reg[4][150]  ( .CLK(n3487), .D(n1698), .Q(
        \inq_ary[4][150] ) );
  LATCHX1_RVT \inq_ary_reg[5][150]  ( .CLK(n3486), .D(n1698), .Q(
        \inq_ary[5][150] ) );
  LATCHX1_RVT \inq_ary_reg[6][150]  ( .CLK(n3485), .D(n1698), .Q(
        \inq_ary[6][150] ) );
  LATCHX1_RVT \inq_ary_reg[7][150]  ( .CLK(n3484), .D(n1698), .Q(
        \inq_ary[7][150] ) );
  LATCHX1_RVT \inq_ary_reg[8][150]  ( .CLK(n3483), .D(n1698), .Q(
        \inq_ary[8][150] ) );
  LATCHX1_RVT \inq_ary_reg[9][150]  ( .CLK(n3482), .D(n1698), .Q(
        \inq_ary[9][150] ) );
  LATCHX1_RVT \inq_ary_reg[10][150]  ( .CLK(n3481), .D(n1698), .Q(
        \inq_ary[10][150] ) );
  LATCHX1_RVT \inq_ary_reg[11][150]  ( .CLK(n3480), .D(n1698), .Q(
        \inq_ary[11][150] ) );
  LATCHX1_RVT \inq_ary_reg[12][150]  ( .CLK(n3479), .D(n1698), .Q(
        \inq_ary[12][150] ) );
  LATCHX1_RVT \inq_ary_reg[13][150]  ( .CLK(n3478), .D(n1698), .Q(
        \inq_ary[13][150] ) );
  LATCHX1_RVT \inq_ary_reg[14][150]  ( .CLK(n3477), .D(n1698), .Q(
        \inq_ary[14][150] ) );
  LATCHX1_RVT \inq_ary_reg[15][150]  ( .CLK(n3476), .D(n1698), .Q(
        \inq_ary[15][150] ) );
  LATCHX1_RVT \dout_reg[150]  ( .CLK(n3492), .D(N412), .Q(dout[150]) );
  LATCHX1_RVT \inq_ary_reg[0][149]  ( .CLK(n3491), .D(n1685), .Q(
        \inq_ary[0][149] ) );
  LATCHX1_RVT \inq_ary_reg[1][149]  ( .CLK(n3490), .D(n1685), .Q(
        \inq_ary[1][149] ) );
  LATCHX1_RVT \inq_ary_reg[2][149]  ( .CLK(n3489), .D(n1685), .Q(
        \inq_ary[2][149] ) );
  LATCHX1_RVT \inq_ary_reg[3][149]  ( .CLK(n3488), .D(n1685), .Q(
        \inq_ary[3][149] ) );
  LATCHX1_RVT \inq_ary_reg[4][149]  ( .CLK(n3487), .D(n1685), .Q(
        \inq_ary[4][149] ) );
  LATCHX1_RVT \inq_ary_reg[5][149]  ( .CLK(n3486), .D(n1685), .Q(
        \inq_ary[5][149] ) );
  LATCHX1_RVT \inq_ary_reg[6][149]  ( .CLK(n3485), .D(n1685), .Q(
        \inq_ary[6][149] ) );
  LATCHX1_RVT \inq_ary_reg[7][149]  ( .CLK(n3484), .D(n1685), .Q(
        \inq_ary[7][149] ) );
  LATCHX1_RVT \inq_ary_reg[8][149]  ( .CLK(n3483), .D(n1685), .Q(
        \inq_ary[8][149] ) );
  LATCHX1_RVT \inq_ary_reg[9][149]  ( .CLK(n3482), .D(n1685), .Q(
        \inq_ary[9][149] ) );
  LATCHX1_RVT \inq_ary_reg[10][149]  ( .CLK(n3481), .D(n1685), .Q(
        \inq_ary[10][149] ) );
  LATCHX1_RVT \inq_ary_reg[11][149]  ( .CLK(n3480), .D(n1685), .Q(
        \inq_ary[11][149] ) );
  LATCHX1_RVT \inq_ary_reg[12][149]  ( .CLK(n3479), .D(n1685), .Q(
        \inq_ary[12][149] ) );
  LATCHX1_RVT \inq_ary_reg[13][149]  ( .CLK(n3478), .D(n1685), .Q(
        \inq_ary[13][149] ) );
  LATCHX1_RVT \inq_ary_reg[14][149]  ( .CLK(n3477), .D(n1685), .Q(
        \inq_ary[14][149] ) );
  LATCHX1_RVT \inq_ary_reg[15][149]  ( .CLK(n3476), .D(n1685), .Q(
        \inq_ary[15][149] ) );
  LATCHX1_RVT \dout_reg[149]  ( .CLK(n3492), .D(N411), .Q(dout[149]) );
  LATCHX1_RVT \inq_ary_reg[0][148]  ( .CLK(n3491), .D(n1672), .Q(
        \inq_ary[0][148] ) );
  LATCHX1_RVT \inq_ary_reg[1][148]  ( .CLK(n3490), .D(n1672), .Q(
        \inq_ary[1][148] ) );
  LATCHX1_RVT \inq_ary_reg[2][148]  ( .CLK(n3489), .D(n1672), .Q(
        \inq_ary[2][148] ) );
  LATCHX1_RVT \inq_ary_reg[3][148]  ( .CLK(n3488), .D(n1672), .Q(
        \inq_ary[3][148] ) );
  LATCHX1_RVT \inq_ary_reg[4][148]  ( .CLK(n3487), .D(n1672), .Q(
        \inq_ary[4][148] ) );
  LATCHX1_RVT \inq_ary_reg[5][148]  ( .CLK(n3486), .D(n1672), .Q(
        \inq_ary[5][148] ) );
  LATCHX1_RVT \inq_ary_reg[6][148]  ( .CLK(n3485), .D(n1672), .Q(
        \inq_ary[6][148] ) );
  LATCHX1_RVT \inq_ary_reg[7][148]  ( .CLK(n3484), .D(n1672), .Q(
        \inq_ary[7][148] ) );
  LATCHX1_RVT \inq_ary_reg[8][148]  ( .CLK(n3483), .D(n1672), .Q(
        \inq_ary[8][148] ) );
  LATCHX1_RVT \inq_ary_reg[9][148]  ( .CLK(n3482), .D(n1672), .Q(
        \inq_ary[9][148] ) );
  LATCHX1_RVT \inq_ary_reg[10][148]  ( .CLK(n3481), .D(n1672), .Q(
        \inq_ary[10][148] ) );
  LATCHX1_RVT \inq_ary_reg[11][148]  ( .CLK(n3480), .D(n1672), .Q(
        \inq_ary[11][148] ) );
  LATCHX1_RVT \inq_ary_reg[12][148]  ( .CLK(n3479), .D(n1672), .Q(
        \inq_ary[12][148] ) );
  LATCHX1_RVT \inq_ary_reg[13][148]  ( .CLK(n3478), .D(n1672), .Q(
        \inq_ary[13][148] ) );
  LATCHX1_RVT \inq_ary_reg[14][148]  ( .CLK(n3477), .D(n1672), .Q(
        \inq_ary[14][148] ) );
  LATCHX1_RVT \inq_ary_reg[15][148]  ( .CLK(n3476), .D(n1672), .Q(
        \inq_ary[15][148] ) );
  LATCHX1_RVT \dout_reg[148]  ( .CLK(n3492), .D(N410), .Q(dout[148]) );
  LATCHX1_RVT \inq_ary_reg[0][147]  ( .CLK(n3491), .D(n3475), .Q(
        \inq_ary[0][147] ) );
  LATCHX1_RVT \inq_ary_reg[1][147]  ( .CLK(n3490), .D(n3475), .Q(
        \inq_ary[1][147] ) );
  LATCHX1_RVT \inq_ary_reg[2][147]  ( .CLK(n3489), .D(n3475), .Q(
        \inq_ary[2][147] ) );
  LATCHX1_RVT \inq_ary_reg[3][147]  ( .CLK(n3488), .D(n3475), .Q(
        \inq_ary[3][147] ) );
  LATCHX1_RVT \inq_ary_reg[4][147]  ( .CLK(n3487), .D(n3475), .Q(
        \inq_ary[4][147] ) );
  LATCHX1_RVT \inq_ary_reg[5][147]  ( .CLK(n3486), .D(n3475), .Q(
        \inq_ary[5][147] ) );
  LATCHX1_RVT \inq_ary_reg[6][147]  ( .CLK(n3485), .D(n3475), .Q(
        \inq_ary[6][147] ) );
  LATCHX1_RVT \inq_ary_reg[7][147]  ( .CLK(n3484), .D(n3475), .Q(
        \inq_ary[7][147] ) );
  LATCHX1_RVT \inq_ary_reg[8][147]  ( .CLK(n3483), .D(n3475), .Q(
        \inq_ary[8][147] ) );
  LATCHX1_RVT \inq_ary_reg[9][147]  ( .CLK(n3482), .D(n3475), .Q(
        \inq_ary[9][147] ) );
  LATCHX1_RVT \inq_ary_reg[10][147]  ( .CLK(n3481), .D(n3475), .Q(
        \inq_ary[10][147] ) );
  LATCHX1_RVT \inq_ary_reg[11][147]  ( .CLK(n3480), .D(n3475), .Q(
        \inq_ary[11][147] ) );
  LATCHX1_RVT \inq_ary_reg[12][147]  ( .CLK(n3479), .D(n3475), .Q(
        \inq_ary[12][147] ) );
  LATCHX1_RVT \inq_ary_reg[13][147]  ( .CLK(n3478), .D(n3475), .Q(
        \inq_ary[13][147] ) );
  LATCHX1_RVT \inq_ary_reg[14][147]  ( .CLK(n3477), .D(n3475), .Q(
        \inq_ary[14][147] ) );
  LATCHX1_RVT \inq_ary_reg[15][147]  ( .CLK(n3476), .D(n3475), .Q(
        \inq_ary[15][147] ) );
  LATCHX1_RVT \dout_reg[147]  ( .CLK(n3492), .D(N409), .Q(dout[147]) );
  LATCHX1_RVT \inq_ary_reg[0][146]  ( .CLK(n3491), .D(n3474), .Q(
        \inq_ary[0][146] ) );
  LATCHX1_RVT \inq_ary_reg[1][146]  ( .CLK(n3490), .D(n3474), .Q(
        \inq_ary[1][146] ) );
  LATCHX1_RVT \inq_ary_reg[2][146]  ( .CLK(n3489), .D(n3474), .Q(
        \inq_ary[2][146] ) );
  LATCHX1_RVT \inq_ary_reg[3][146]  ( .CLK(n3488), .D(n3474), .Q(
        \inq_ary[3][146] ) );
  LATCHX1_RVT \inq_ary_reg[4][146]  ( .CLK(n3487), .D(n3474), .Q(
        \inq_ary[4][146] ) );
  LATCHX1_RVT \inq_ary_reg[5][146]  ( .CLK(n3486), .D(n3474), .Q(
        \inq_ary[5][146] ) );
  LATCHX1_RVT \inq_ary_reg[6][146]  ( .CLK(n3485), .D(n3474), .Q(
        \inq_ary[6][146] ) );
  LATCHX1_RVT \inq_ary_reg[7][146]  ( .CLK(n3484), .D(n3474), .Q(
        \inq_ary[7][146] ) );
  LATCHX1_RVT \inq_ary_reg[8][146]  ( .CLK(n3483), .D(n3474), .Q(
        \inq_ary[8][146] ) );
  LATCHX1_RVT \inq_ary_reg[9][146]  ( .CLK(n3482), .D(n3474), .Q(
        \inq_ary[9][146] ) );
  LATCHX1_RVT \inq_ary_reg[10][146]  ( .CLK(n3481), .D(n3474), .Q(
        \inq_ary[10][146] ) );
  LATCHX1_RVT \inq_ary_reg[11][146]  ( .CLK(n3480), .D(n3474), .Q(
        \inq_ary[11][146] ) );
  LATCHX1_RVT \inq_ary_reg[12][146]  ( .CLK(n3479), .D(n3474), .Q(
        \inq_ary[12][146] ) );
  LATCHX1_RVT \inq_ary_reg[13][146]  ( .CLK(n3478), .D(n3474), .Q(
        \inq_ary[13][146] ) );
  LATCHX1_RVT \inq_ary_reg[14][146]  ( .CLK(n3477), .D(n3474), .Q(
        \inq_ary[14][146] ) );
  LATCHX1_RVT \inq_ary_reg[15][146]  ( .CLK(n3476), .D(n3474), .Q(
        \inq_ary[15][146] ) );
  LATCHX1_RVT \dout_reg[146]  ( .CLK(n3492), .D(N408), .Q(dout[146]) );
  LATCHX1_RVT \inq_ary_reg[0][145]  ( .CLK(n3491), .D(n3473), .Q(
        \inq_ary[0][145] ) );
  LATCHX1_RVT \inq_ary_reg[1][145]  ( .CLK(n3490), .D(n3473), .Q(
        \inq_ary[1][145] ) );
  LATCHX1_RVT \inq_ary_reg[2][145]  ( .CLK(n3489), .D(n3473), .Q(
        \inq_ary[2][145] ) );
  LATCHX1_RVT \inq_ary_reg[3][145]  ( .CLK(n3488), .D(n3473), .Q(
        \inq_ary[3][145] ) );
  LATCHX1_RVT \inq_ary_reg[4][145]  ( .CLK(n3487), .D(n3473), .Q(
        \inq_ary[4][145] ) );
  LATCHX1_RVT \inq_ary_reg[5][145]  ( .CLK(n3486), .D(n3473), .Q(
        \inq_ary[5][145] ) );
  LATCHX1_RVT \inq_ary_reg[6][145]  ( .CLK(n3485), .D(n3473), .Q(
        \inq_ary[6][145] ) );
  LATCHX1_RVT \inq_ary_reg[7][145]  ( .CLK(n3484), .D(n3473), .Q(
        \inq_ary[7][145] ) );
  LATCHX1_RVT \inq_ary_reg[8][145]  ( .CLK(n3483), .D(n3473), .Q(
        \inq_ary[8][145] ) );
  LATCHX1_RVT \inq_ary_reg[9][145]  ( .CLK(n3482), .D(n3473), .Q(
        \inq_ary[9][145] ) );
  LATCHX1_RVT \inq_ary_reg[10][145]  ( .CLK(n3481), .D(n3473), .Q(
        \inq_ary[10][145] ) );
  LATCHX1_RVT \inq_ary_reg[11][145]  ( .CLK(n3480), .D(n3473), .Q(
        \inq_ary[11][145] ) );
  LATCHX1_RVT \inq_ary_reg[12][145]  ( .CLK(n3479), .D(n3473), .Q(
        \inq_ary[12][145] ) );
  LATCHX1_RVT \inq_ary_reg[13][145]  ( .CLK(n3478), .D(n3473), .Q(
        \inq_ary[13][145] ) );
  LATCHX1_RVT \inq_ary_reg[14][145]  ( .CLK(n3477), .D(n3473), .Q(
        \inq_ary[14][145] ) );
  LATCHX1_RVT \inq_ary_reg[15][145]  ( .CLK(n3476), .D(n3473), .Q(
        \inq_ary[15][145] ) );
  LATCHX1_RVT \dout_reg[145]  ( .CLK(n3492), .D(N407), .Q(dout[145]) );
  LATCHX1_RVT \inq_ary_reg[0][144]  ( .CLK(n3491), .D(n3472), .Q(
        \inq_ary[0][144] ) );
  LATCHX1_RVT \inq_ary_reg[1][144]  ( .CLK(n3490), .D(n3472), .Q(
        \inq_ary[1][144] ) );
  LATCHX1_RVT \inq_ary_reg[2][144]  ( .CLK(n3489), .D(n3472), .Q(
        \inq_ary[2][144] ) );
  LATCHX1_RVT \inq_ary_reg[3][144]  ( .CLK(n3488), .D(n3472), .Q(
        \inq_ary[3][144] ) );
  LATCHX1_RVT \inq_ary_reg[4][144]  ( .CLK(n3487), .D(n3472), .Q(
        \inq_ary[4][144] ) );
  LATCHX1_RVT \inq_ary_reg[5][144]  ( .CLK(n3486), .D(n3472), .Q(
        \inq_ary[5][144] ) );
  LATCHX1_RVT \inq_ary_reg[6][144]  ( .CLK(n3485), .D(n3472), .Q(
        \inq_ary[6][144] ) );
  LATCHX1_RVT \inq_ary_reg[7][144]  ( .CLK(n3484), .D(n3472), .Q(
        \inq_ary[7][144] ) );
  LATCHX1_RVT \inq_ary_reg[8][144]  ( .CLK(n3483), .D(n3472), .Q(
        \inq_ary[8][144] ) );
  LATCHX1_RVT \inq_ary_reg[9][144]  ( .CLK(n3482), .D(n3472), .Q(
        \inq_ary[9][144] ) );
  LATCHX1_RVT \inq_ary_reg[10][144]  ( .CLK(n3481), .D(n3472), .Q(
        \inq_ary[10][144] ) );
  LATCHX1_RVT \inq_ary_reg[11][144]  ( .CLK(n3480), .D(n3472), .Q(
        \inq_ary[11][144] ) );
  LATCHX1_RVT \inq_ary_reg[12][144]  ( .CLK(n3479), .D(n3472), .Q(
        \inq_ary[12][144] ) );
  LATCHX1_RVT \inq_ary_reg[13][144]  ( .CLK(n3478), .D(n3472), .Q(
        \inq_ary[13][144] ) );
  LATCHX1_RVT \inq_ary_reg[14][144]  ( .CLK(n3477), .D(n3472), .Q(
        \inq_ary[14][144] ) );
  LATCHX1_RVT \inq_ary_reg[15][144]  ( .CLK(n3476), .D(n3472), .Q(
        \inq_ary[15][144] ) );
  LATCHX1_RVT \dout_reg[144]  ( .CLK(n3492), .D(N406), .Q(dout[144]) );
  LATCHX1_RVT \inq_ary_reg[0][143]  ( .CLK(n3491), .D(n3470), .Q(
        \inq_ary[0][143] ) );
  LATCHX1_RVT \inq_ary_reg[1][143]  ( .CLK(n3490), .D(n3470), .Q(
        \inq_ary[1][143] ) );
  LATCHX1_RVT \inq_ary_reg[2][143]  ( .CLK(n3489), .D(n3470), .Q(
        \inq_ary[2][143] ) );
  LATCHX1_RVT \inq_ary_reg[3][143]  ( .CLK(n3488), .D(n3470), .Q(
        \inq_ary[3][143] ) );
  LATCHX1_RVT \inq_ary_reg[4][143]  ( .CLK(n3487), .D(n3470), .Q(
        \inq_ary[4][143] ) );
  LATCHX1_RVT \inq_ary_reg[5][143]  ( .CLK(n3486), .D(n3470), .Q(
        \inq_ary[5][143] ) );
  LATCHX1_RVT \inq_ary_reg[6][143]  ( .CLK(n3485), .D(n3470), .Q(
        \inq_ary[6][143] ) );
  LATCHX1_RVT \inq_ary_reg[7][143]  ( .CLK(n3484), .D(n3470), .Q(
        \inq_ary[7][143] ) );
  LATCHX1_RVT \inq_ary_reg[8][143]  ( .CLK(n3483), .D(n3470), .Q(
        \inq_ary[8][143] ) );
  LATCHX1_RVT \inq_ary_reg[9][143]  ( .CLK(n3482), .D(n3470), .Q(
        \inq_ary[9][143] ) );
  LATCHX1_RVT \inq_ary_reg[10][143]  ( .CLK(n3481), .D(n3470), .Q(
        \inq_ary[10][143] ) );
  LATCHX1_RVT \inq_ary_reg[11][143]  ( .CLK(n3480), .D(n3470), .Q(
        \inq_ary[11][143] ) );
  LATCHX1_RVT \inq_ary_reg[12][143]  ( .CLK(n3479), .D(n3470), .Q(
        \inq_ary[12][143] ) );
  LATCHX1_RVT \inq_ary_reg[13][143]  ( .CLK(n3478), .D(n3470), .Q(
        \inq_ary[13][143] ) );
  LATCHX1_RVT \inq_ary_reg[14][143]  ( .CLK(n3477), .D(n3470), .Q(
        \inq_ary[14][143] ) );
  LATCHX1_RVT \inq_ary_reg[15][143]  ( .CLK(n3476), .D(n3470), .Q(
        \inq_ary[15][143] ) );
  LATCHX1_RVT \dout_reg[143]  ( .CLK(n3492), .D(N405), .Q(dout[143]) );
  LATCHX1_RVT \inq_ary_reg[0][142]  ( .CLK(n3491), .D(n3468), .Q(
        \inq_ary[0][142] ) );
  LATCHX1_RVT \inq_ary_reg[1][142]  ( .CLK(n3490), .D(n3468), .Q(
        \inq_ary[1][142] ) );
  LATCHX1_RVT \inq_ary_reg[2][142]  ( .CLK(n3489), .D(n3468), .Q(
        \inq_ary[2][142] ) );
  LATCHX1_RVT \inq_ary_reg[3][142]  ( .CLK(n3488), .D(n3468), .Q(
        \inq_ary[3][142] ) );
  LATCHX1_RVT \inq_ary_reg[4][142]  ( .CLK(n3487), .D(n3468), .Q(
        \inq_ary[4][142] ) );
  LATCHX1_RVT \inq_ary_reg[5][142]  ( .CLK(n3486), .D(n3468), .Q(
        \inq_ary[5][142] ) );
  LATCHX1_RVT \inq_ary_reg[6][142]  ( .CLK(n3485), .D(n3468), .Q(
        \inq_ary[6][142] ) );
  LATCHX1_RVT \inq_ary_reg[7][142]  ( .CLK(n3484), .D(n3468), .Q(
        \inq_ary[7][142] ) );
  LATCHX1_RVT \inq_ary_reg[8][142]  ( .CLK(n3483), .D(n3468), .Q(
        \inq_ary[8][142] ) );
  LATCHX1_RVT \inq_ary_reg[9][142]  ( .CLK(n3482), .D(n3468), .Q(
        \inq_ary[9][142] ) );
  LATCHX1_RVT \inq_ary_reg[10][142]  ( .CLK(n3481), .D(n3468), .Q(
        \inq_ary[10][142] ) );
  LATCHX1_RVT \inq_ary_reg[11][142]  ( .CLK(n3480), .D(n3468), .Q(
        \inq_ary[11][142] ) );
  LATCHX1_RVT \inq_ary_reg[12][142]  ( .CLK(n3479), .D(n3468), .Q(
        \inq_ary[12][142] ) );
  LATCHX1_RVT \inq_ary_reg[13][142]  ( .CLK(n3478), .D(n3468), .Q(
        \inq_ary[13][142] ) );
  LATCHX1_RVT \inq_ary_reg[14][142]  ( .CLK(n3477), .D(n3468), .Q(
        \inq_ary[14][142] ) );
  LATCHX1_RVT \inq_ary_reg[15][142]  ( .CLK(n3476), .D(n3468), .Q(
        \inq_ary[15][142] ) );
  LATCHX1_RVT \dout_reg[142]  ( .CLK(n3492), .D(N404), .Q(dout[142]) );
  LATCHX1_RVT \inq_ary_reg[0][141]  ( .CLK(n3491), .D(n3466), .Q(
        \inq_ary[0][141] ) );
  LATCHX1_RVT \inq_ary_reg[1][141]  ( .CLK(n3490), .D(n3466), .Q(
        \inq_ary[1][141] ) );
  LATCHX1_RVT \inq_ary_reg[2][141]  ( .CLK(n3489), .D(n3466), .Q(
        \inq_ary[2][141] ) );
  LATCHX1_RVT \inq_ary_reg[3][141]  ( .CLK(n3488), .D(n3466), .Q(
        \inq_ary[3][141] ) );
  LATCHX1_RVT \inq_ary_reg[4][141]  ( .CLK(n3487), .D(n3466), .Q(
        \inq_ary[4][141] ) );
  LATCHX1_RVT \inq_ary_reg[5][141]  ( .CLK(n3486), .D(n3466), .Q(
        \inq_ary[5][141] ) );
  LATCHX1_RVT \inq_ary_reg[6][141]  ( .CLK(n3485), .D(n3466), .Q(
        \inq_ary[6][141] ) );
  LATCHX1_RVT \inq_ary_reg[7][141]  ( .CLK(n3484), .D(n3466), .Q(
        \inq_ary[7][141] ) );
  LATCHX1_RVT \inq_ary_reg[8][141]  ( .CLK(n3483), .D(n3466), .Q(
        \inq_ary[8][141] ) );
  LATCHX1_RVT \inq_ary_reg[9][141]  ( .CLK(n3482), .D(n3466), .Q(
        \inq_ary[9][141] ) );
  LATCHX1_RVT \inq_ary_reg[10][141]  ( .CLK(n3481), .D(n3466), .Q(
        \inq_ary[10][141] ) );
  LATCHX1_RVT \inq_ary_reg[11][141]  ( .CLK(n3480), .D(n3466), .Q(
        \inq_ary[11][141] ) );
  LATCHX1_RVT \inq_ary_reg[12][141]  ( .CLK(n3479), .D(n3466), .Q(
        \inq_ary[12][141] ) );
  LATCHX1_RVT \inq_ary_reg[13][141]  ( .CLK(n3478), .D(n3466), .Q(
        \inq_ary[13][141] ) );
  LATCHX1_RVT \inq_ary_reg[14][141]  ( .CLK(n3477), .D(n3466), .Q(
        \inq_ary[14][141] ) );
  LATCHX1_RVT \inq_ary_reg[15][141]  ( .CLK(n3476), .D(n3466), .Q(
        \inq_ary[15][141] ) );
  LATCHX1_RVT \dout_reg[141]  ( .CLK(n3492), .D(N403), .Q(dout[141]) );
  LATCHX1_RVT \inq_ary_reg[0][140]  ( .CLK(n3491), .D(n3464), .Q(
        \inq_ary[0][140] ) );
  LATCHX1_RVT \inq_ary_reg[1][140]  ( .CLK(n3490), .D(n3464), .Q(
        \inq_ary[1][140] ) );
  LATCHX1_RVT \inq_ary_reg[2][140]  ( .CLK(n3489), .D(n3464), .Q(
        \inq_ary[2][140] ) );
  LATCHX1_RVT \inq_ary_reg[3][140]  ( .CLK(n3488), .D(n3464), .Q(
        \inq_ary[3][140] ) );
  LATCHX1_RVT \inq_ary_reg[4][140]  ( .CLK(n3487), .D(n3464), .Q(
        \inq_ary[4][140] ) );
  LATCHX1_RVT \inq_ary_reg[5][140]  ( .CLK(n3486), .D(n3464), .Q(
        \inq_ary[5][140] ) );
  LATCHX1_RVT \inq_ary_reg[6][140]  ( .CLK(n3485), .D(n3464), .Q(
        \inq_ary[6][140] ) );
  LATCHX1_RVT \inq_ary_reg[7][140]  ( .CLK(n3484), .D(n3464), .Q(
        \inq_ary[7][140] ) );
  LATCHX1_RVT \inq_ary_reg[8][140]  ( .CLK(n3483), .D(n3464), .Q(
        \inq_ary[8][140] ) );
  LATCHX1_RVT \inq_ary_reg[9][140]  ( .CLK(n3482), .D(n3464), .Q(
        \inq_ary[9][140] ) );
  LATCHX1_RVT \inq_ary_reg[10][140]  ( .CLK(n3481), .D(n3464), .Q(
        \inq_ary[10][140] ) );
  LATCHX1_RVT \inq_ary_reg[11][140]  ( .CLK(n3480), .D(n3464), .Q(
        \inq_ary[11][140] ) );
  LATCHX1_RVT \inq_ary_reg[12][140]  ( .CLK(n3479), .D(n3464), .Q(
        \inq_ary[12][140] ) );
  LATCHX1_RVT \inq_ary_reg[13][140]  ( .CLK(n3478), .D(n3464), .Q(
        \inq_ary[13][140] ) );
  LATCHX1_RVT \inq_ary_reg[14][140]  ( .CLK(n3477), .D(n3464), .Q(
        \inq_ary[14][140] ) );
  LATCHX1_RVT \inq_ary_reg[15][140]  ( .CLK(n3476), .D(n3464), .Q(
        \inq_ary[15][140] ) );
  LATCHX1_RVT \dout_reg[140]  ( .CLK(n3492), .D(N402), .Q(dout[140]) );
  LATCHX1_RVT \inq_ary_reg[0][139]  ( .CLK(n3491), .D(n3471), .Q(
        \inq_ary[0][139] ) );
  LATCHX1_RVT \inq_ary_reg[1][139]  ( .CLK(n3490), .D(n3471), .Q(
        \inq_ary[1][139] ) );
  LATCHX1_RVT \inq_ary_reg[2][139]  ( .CLK(n3489), .D(n3471), .Q(
        \inq_ary[2][139] ) );
  LATCHX1_RVT \inq_ary_reg[3][139]  ( .CLK(n3488), .D(n3471), .Q(
        \inq_ary[3][139] ) );
  LATCHX1_RVT \inq_ary_reg[4][139]  ( .CLK(n3487), .D(n3471), .Q(
        \inq_ary[4][139] ) );
  LATCHX1_RVT \inq_ary_reg[5][139]  ( .CLK(n3486), .D(n3471), .Q(
        \inq_ary[5][139] ) );
  LATCHX1_RVT \inq_ary_reg[6][139]  ( .CLK(n3485), .D(n3471), .Q(
        \inq_ary[6][139] ) );
  LATCHX1_RVT \inq_ary_reg[7][139]  ( .CLK(n3484), .D(n3471), .Q(
        \inq_ary[7][139] ) );
  LATCHX1_RVT \inq_ary_reg[8][139]  ( .CLK(n3483), .D(n3471), .Q(
        \inq_ary[8][139] ) );
  LATCHX1_RVT \inq_ary_reg[9][139]  ( .CLK(n3482), .D(n3471), .Q(
        \inq_ary[9][139] ) );
  LATCHX1_RVT \inq_ary_reg[10][139]  ( .CLK(n3481), .D(n3471), .Q(
        \inq_ary[10][139] ) );
  LATCHX1_RVT \inq_ary_reg[11][139]  ( .CLK(n3480), .D(n3471), .Q(
        \inq_ary[11][139] ) );
  LATCHX1_RVT \inq_ary_reg[12][139]  ( .CLK(n3479), .D(n3471), .Q(
        \inq_ary[12][139] ) );
  LATCHX1_RVT \inq_ary_reg[13][139]  ( .CLK(n3478), .D(n3471), .Q(
        \inq_ary[13][139] ) );
  LATCHX1_RVT \inq_ary_reg[14][139]  ( .CLK(n3477), .D(n3471), .Q(
        \inq_ary[14][139] ) );
  LATCHX1_RVT \inq_ary_reg[15][139]  ( .CLK(n3476), .D(n3471), .Q(
        \inq_ary[15][139] ) );
  LATCHX1_RVT \dout_reg[139]  ( .CLK(n3492), .D(N401), .Q(dout[139]) );
  LATCHX1_RVT \inq_ary_reg[0][138]  ( .CLK(n3491), .D(n3469), .Q(
        \inq_ary[0][138] ) );
  LATCHX1_RVT \inq_ary_reg[1][138]  ( .CLK(n3490), .D(n3469), .Q(
        \inq_ary[1][138] ) );
  LATCHX1_RVT \inq_ary_reg[2][138]  ( .CLK(n3489), .D(n3469), .Q(
        \inq_ary[2][138] ) );
  LATCHX1_RVT \inq_ary_reg[3][138]  ( .CLK(n3488), .D(n3469), .Q(
        \inq_ary[3][138] ) );
  LATCHX1_RVT \inq_ary_reg[4][138]  ( .CLK(n3487), .D(n3469), .Q(
        \inq_ary[4][138] ) );
  LATCHX1_RVT \inq_ary_reg[5][138]  ( .CLK(n3486), .D(n3469), .Q(
        \inq_ary[5][138] ) );
  LATCHX1_RVT \inq_ary_reg[6][138]  ( .CLK(n3485), .D(n3469), .Q(
        \inq_ary[6][138] ) );
  LATCHX1_RVT \inq_ary_reg[7][138]  ( .CLK(n3484), .D(n3469), .Q(
        \inq_ary[7][138] ) );
  LATCHX1_RVT \inq_ary_reg[8][138]  ( .CLK(n3483), .D(n3469), .Q(
        \inq_ary[8][138] ) );
  LATCHX1_RVT \inq_ary_reg[9][138]  ( .CLK(n3482), .D(n3469), .Q(
        \inq_ary[9][138] ) );
  LATCHX1_RVT \inq_ary_reg[10][138]  ( .CLK(n3481), .D(n3469), .Q(
        \inq_ary[10][138] ) );
  LATCHX1_RVT \inq_ary_reg[11][138]  ( .CLK(n3480), .D(n3469), .Q(
        \inq_ary[11][138] ) );
  LATCHX1_RVT \inq_ary_reg[12][138]  ( .CLK(n3479), .D(n3469), .Q(
        \inq_ary[12][138] ) );
  LATCHX1_RVT \inq_ary_reg[13][138]  ( .CLK(n3478), .D(n3469), .Q(
        \inq_ary[13][138] ) );
  LATCHX1_RVT \inq_ary_reg[14][138]  ( .CLK(n3477), .D(n3469), .Q(
        \inq_ary[14][138] ) );
  LATCHX1_RVT \inq_ary_reg[15][138]  ( .CLK(n3476), .D(n3469), .Q(
        \inq_ary[15][138] ) );
  LATCHX1_RVT \dout_reg[138]  ( .CLK(n3492), .D(N400), .Q(dout[138]) );
  LATCHX1_RVT \inq_ary_reg[0][137]  ( .CLK(n3491), .D(n3467), .Q(
        \inq_ary[0][137] ) );
  LATCHX1_RVT \inq_ary_reg[1][137]  ( .CLK(n3490), .D(n3467), .Q(
        \inq_ary[1][137] ) );
  LATCHX1_RVT \inq_ary_reg[2][137]  ( .CLK(n3489), .D(n3467), .Q(
        \inq_ary[2][137] ) );
  LATCHX1_RVT \inq_ary_reg[3][137]  ( .CLK(n3488), .D(n3467), .Q(
        \inq_ary[3][137] ) );
  LATCHX1_RVT \inq_ary_reg[4][137]  ( .CLK(n3487), .D(n3467), .Q(
        \inq_ary[4][137] ) );
  LATCHX1_RVT \inq_ary_reg[5][137]  ( .CLK(n3486), .D(n3467), .Q(
        \inq_ary[5][137] ) );
  LATCHX1_RVT \inq_ary_reg[6][137]  ( .CLK(n3485), .D(n3467), .Q(
        \inq_ary[6][137] ) );
  LATCHX1_RVT \inq_ary_reg[7][137]  ( .CLK(n3484), .D(n3467), .Q(
        \inq_ary[7][137] ) );
  LATCHX1_RVT \inq_ary_reg[8][137]  ( .CLK(n3483), .D(n3467), .Q(
        \inq_ary[8][137] ) );
  LATCHX1_RVT \inq_ary_reg[9][137]  ( .CLK(n3482), .D(n3467), .Q(
        \inq_ary[9][137] ) );
  LATCHX1_RVT \inq_ary_reg[10][137]  ( .CLK(n3481), .D(n3467), .Q(
        \inq_ary[10][137] ) );
  LATCHX1_RVT \inq_ary_reg[11][137]  ( .CLK(n3480), .D(n3467), .Q(
        \inq_ary[11][137] ) );
  LATCHX1_RVT \inq_ary_reg[12][137]  ( .CLK(n3479), .D(n3467), .Q(
        \inq_ary[12][137] ) );
  LATCHX1_RVT \inq_ary_reg[13][137]  ( .CLK(n3478), .D(n3467), .Q(
        \inq_ary[13][137] ) );
  LATCHX1_RVT \inq_ary_reg[14][137]  ( .CLK(n3477), .D(n3467), .Q(
        \inq_ary[14][137] ) );
  LATCHX1_RVT \inq_ary_reg[15][137]  ( .CLK(n3476), .D(n3467), .Q(
        \inq_ary[15][137] ) );
  LATCHX1_RVT \dout_reg[137]  ( .CLK(n3492), .D(N399), .Q(dout[137]) );
  LATCHX1_RVT \inq_ary_reg[0][136]  ( .CLK(n3491), .D(n3465), .Q(
        \inq_ary[0][136] ) );
  LATCHX1_RVT \inq_ary_reg[1][136]  ( .CLK(n3490), .D(n3465), .Q(
        \inq_ary[1][136] ) );
  LATCHX1_RVT \inq_ary_reg[2][136]  ( .CLK(n3489), .D(n3465), .Q(
        \inq_ary[2][136] ) );
  LATCHX1_RVT \inq_ary_reg[3][136]  ( .CLK(n3488), .D(n3465), .Q(
        \inq_ary[3][136] ) );
  LATCHX1_RVT \inq_ary_reg[4][136]  ( .CLK(n3487), .D(n3465), .Q(
        \inq_ary[4][136] ) );
  LATCHX1_RVT \inq_ary_reg[5][136]  ( .CLK(n3486), .D(n3465), .Q(
        \inq_ary[5][136] ) );
  LATCHX1_RVT \inq_ary_reg[6][136]  ( .CLK(n3485), .D(n3465), .Q(
        \inq_ary[6][136] ) );
  LATCHX1_RVT \inq_ary_reg[7][136]  ( .CLK(n3484), .D(n3465), .Q(
        \inq_ary[7][136] ) );
  LATCHX1_RVT \inq_ary_reg[8][136]  ( .CLK(n3483), .D(n3465), .Q(
        \inq_ary[8][136] ) );
  LATCHX1_RVT \inq_ary_reg[9][136]  ( .CLK(n3482), .D(n3465), .Q(
        \inq_ary[9][136] ) );
  LATCHX1_RVT \inq_ary_reg[10][136]  ( .CLK(n3481), .D(n3465), .Q(
        \inq_ary[10][136] ) );
  LATCHX1_RVT \inq_ary_reg[11][136]  ( .CLK(n3480), .D(n3465), .Q(
        \inq_ary[11][136] ) );
  LATCHX1_RVT \inq_ary_reg[12][136]  ( .CLK(n3479), .D(n3465), .Q(
        \inq_ary[12][136] ) );
  LATCHX1_RVT \inq_ary_reg[13][136]  ( .CLK(n3478), .D(n3465), .Q(
        \inq_ary[13][136] ) );
  LATCHX1_RVT \inq_ary_reg[14][136]  ( .CLK(n3477), .D(n3465), .Q(
        \inq_ary[14][136] ) );
  LATCHX1_RVT \inq_ary_reg[15][136]  ( .CLK(n3476), .D(n3465), .Q(
        \inq_ary[15][136] ) );
  LATCHX1_RVT \dout_reg[136]  ( .CLK(n3492), .D(N398), .Q(dout[136]) );
  LATCHX1_RVT \inq_ary_reg[0][135]  ( .CLK(n3491), .D(n3462), .Q(
        \inq_ary[0][135] ) );
  LATCHX1_RVT \inq_ary_reg[1][135]  ( .CLK(n3490), .D(n3462), .Q(
        \inq_ary[1][135] ) );
  LATCHX1_RVT \inq_ary_reg[2][135]  ( .CLK(n3489), .D(n3462), .Q(
        \inq_ary[2][135] ) );
  LATCHX1_RVT \inq_ary_reg[3][135]  ( .CLK(n3488), .D(n3462), .Q(
        \inq_ary[3][135] ) );
  LATCHX1_RVT \inq_ary_reg[4][135]  ( .CLK(n3487), .D(n3462), .Q(
        \inq_ary[4][135] ) );
  LATCHX1_RVT \inq_ary_reg[5][135]  ( .CLK(n3486), .D(n3462), .Q(
        \inq_ary[5][135] ) );
  LATCHX1_RVT \inq_ary_reg[6][135]  ( .CLK(n3485), .D(n3462), .Q(
        \inq_ary[6][135] ) );
  LATCHX1_RVT \inq_ary_reg[7][135]  ( .CLK(n3484), .D(n3462), .Q(
        \inq_ary[7][135] ) );
  LATCHX1_RVT \inq_ary_reg[8][135]  ( .CLK(n3483), .D(n3462), .Q(
        \inq_ary[8][135] ) );
  LATCHX1_RVT \inq_ary_reg[9][135]  ( .CLK(n3482), .D(n3462), .Q(
        \inq_ary[9][135] ) );
  LATCHX1_RVT \inq_ary_reg[10][135]  ( .CLK(n3481), .D(n3462), .Q(
        \inq_ary[10][135] ) );
  LATCHX1_RVT \inq_ary_reg[11][135]  ( .CLK(n3480), .D(n3462), .Q(
        \inq_ary[11][135] ) );
  LATCHX1_RVT \inq_ary_reg[12][135]  ( .CLK(n3479), .D(n3462), .Q(
        \inq_ary[12][135] ) );
  LATCHX1_RVT \inq_ary_reg[13][135]  ( .CLK(n3478), .D(n3462), .Q(
        \inq_ary[13][135] ) );
  LATCHX1_RVT \inq_ary_reg[14][135]  ( .CLK(n3477), .D(n3462), .Q(
        \inq_ary[14][135] ) );
  LATCHX1_RVT \inq_ary_reg[15][135]  ( .CLK(n3476), .D(n3462), .Q(
        \inq_ary[15][135] ) );
  LATCHX1_RVT \dout_reg[135]  ( .CLK(n3492), .D(N397), .Q(dout[135]) );
  LATCHX1_RVT \inq_ary_reg[0][134]  ( .CLK(n3491), .D(n3460), .Q(
        \inq_ary[0][134] ) );
  LATCHX1_RVT \inq_ary_reg[1][134]  ( .CLK(n3490), .D(n3460), .Q(
        \inq_ary[1][134] ) );
  LATCHX1_RVT \inq_ary_reg[2][134]  ( .CLK(n3489), .D(n3460), .Q(
        \inq_ary[2][134] ) );
  LATCHX1_RVT \inq_ary_reg[3][134]  ( .CLK(n3488), .D(n3460), .Q(
        \inq_ary[3][134] ) );
  LATCHX1_RVT \inq_ary_reg[4][134]  ( .CLK(n3487), .D(n3460), .Q(
        \inq_ary[4][134] ) );
  LATCHX1_RVT \inq_ary_reg[5][134]  ( .CLK(n3486), .D(n3460), .Q(
        \inq_ary[5][134] ) );
  LATCHX1_RVT \inq_ary_reg[6][134]  ( .CLK(n3485), .D(n3460), .Q(
        \inq_ary[6][134] ) );
  LATCHX1_RVT \inq_ary_reg[7][134]  ( .CLK(n3484), .D(n3460), .Q(
        \inq_ary[7][134] ) );
  LATCHX1_RVT \inq_ary_reg[8][134]  ( .CLK(n3483), .D(n3460), .Q(
        \inq_ary[8][134] ) );
  LATCHX1_RVT \inq_ary_reg[9][134]  ( .CLK(n3482), .D(n3460), .Q(
        \inq_ary[9][134] ) );
  LATCHX1_RVT \inq_ary_reg[10][134]  ( .CLK(n3481), .D(n3460), .Q(
        \inq_ary[10][134] ) );
  LATCHX1_RVT \inq_ary_reg[11][134]  ( .CLK(n3480), .D(n3460), .Q(
        \inq_ary[11][134] ) );
  LATCHX1_RVT \inq_ary_reg[12][134]  ( .CLK(n3479), .D(n3460), .Q(
        \inq_ary[12][134] ) );
  LATCHX1_RVT \inq_ary_reg[13][134]  ( .CLK(n3478), .D(n3460), .Q(
        \inq_ary[13][134] ) );
  LATCHX1_RVT \inq_ary_reg[14][134]  ( .CLK(n3477), .D(n3460), .Q(
        \inq_ary[14][134] ) );
  LATCHX1_RVT \inq_ary_reg[15][134]  ( .CLK(n3476), .D(n3460), .Q(
        \inq_ary[15][134] ) );
  LATCHX1_RVT \dout_reg[134]  ( .CLK(n3492), .D(N396), .Q(dout[134]) );
  LATCHX1_RVT \inq_ary_reg[0][133]  ( .CLK(n3491), .D(n3458), .Q(
        \inq_ary[0][133] ) );
  LATCHX1_RVT \inq_ary_reg[1][133]  ( .CLK(n3490), .D(n3458), .Q(
        \inq_ary[1][133] ) );
  LATCHX1_RVT \inq_ary_reg[2][133]  ( .CLK(n3489), .D(n3458), .Q(
        \inq_ary[2][133] ) );
  LATCHX1_RVT \inq_ary_reg[3][133]  ( .CLK(n3488), .D(n3458), .Q(
        \inq_ary[3][133] ) );
  LATCHX1_RVT \inq_ary_reg[4][133]  ( .CLK(n3487), .D(n3458), .Q(
        \inq_ary[4][133] ) );
  LATCHX1_RVT \inq_ary_reg[5][133]  ( .CLK(n3486), .D(n3458), .Q(
        \inq_ary[5][133] ) );
  LATCHX1_RVT \inq_ary_reg[6][133]  ( .CLK(n3485), .D(n3458), .Q(
        \inq_ary[6][133] ) );
  LATCHX1_RVT \inq_ary_reg[7][133]  ( .CLK(n3484), .D(n3458), .Q(
        \inq_ary[7][133] ) );
  LATCHX1_RVT \inq_ary_reg[8][133]  ( .CLK(n3483), .D(n3458), .Q(
        \inq_ary[8][133] ) );
  LATCHX1_RVT \inq_ary_reg[9][133]  ( .CLK(n3482), .D(n3458), .Q(
        \inq_ary[9][133] ) );
  LATCHX1_RVT \inq_ary_reg[10][133]  ( .CLK(n3481), .D(n3458), .Q(
        \inq_ary[10][133] ) );
  LATCHX1_RVT \inq_ary_reg[11][133]  ( .CLK(n3480), .D(n3458), .Q(
        \inq_ary[11][133] ) );
  LATCHX1_RVT \inq_ary_reg[12][133]  ( .CLK(n3479), .D(n3458), .Q(
        \inq_ary[12][133] ) );
  LATCHX1_RVT \inq_ary_reg[13][133]  ( .CLK(n3478), .D(n3458), .Q(
        \inq_ary[13][133] ) );
  LATCHX1_RVT \inq_ary_reg[14][133]  ( .CLK(n3477), .D(n3458), .Q(
        \inq_ary[14][133] ) );
  LATCHX1_RVT \inq_ary_reg[15][133]  ( .CLK(n3476), .D(n3458), .Q(
        \inq_ary[15][133] ) );
  LATCHX1_RVT \dout_reg[133]  ( .CLK(n3492), .D(N395), .Q(dout[133]) );
  LATCHX1_RVT \inq_ary_reg[0][132]  ( .CLK(n3491), .D(n3456), .Q(
        \inq_ary[0][132] ) );
  LATCHX1_RVT \inq_ary_reg[1][132]  ( .CLK(n3490), .D(n3456), .Q(
        \inq_ary[1][132] ) );
  LATCHX1_RVT \inq_ary_reg[2][132]  ( .CLK(n3489), .D(n3456), .Q(
        \inq_ary[2][132] ) );
  LATCHX1_RVT \inq_ary_reg[3][132]  ( .CLK(n3488), .D(n3456), .Q(
        \inq_ary[3][132] ) );
  LATCHX1_RVT \inq_ary_reg[4][132]  ( .CLK(n3487), .D(n3456), .Q(
        \inq_ary[4][132] ) );
  LATCHX1_RVT \inq_ary_reg[5][132]  ( .CLK(n3486), .D(n3456), .Q(
        \inq_ary[5][132] ) );
  LATCHX1_RVT \inq_ary_reg[6][132]  ( .CLK(n3485), .D(n3456), .Q(
        \inq_ary[6][132] ) );
  LATCHX1_RVT \inq_ary_reg[7][132]  ( .CLK(n3484), .D(n3456), .Q(
        \inq_ary[7][132] ) );
  LATCHX1_RVT \inq_ary_reg[8][132]  ( .CLK(n3483), .D(n3456), .Q(
        \inq_ary[8][132] ) );
  LATCHX1_RVT \inq_ary_reg[9][132]  ( .CLK(n3482), .D(n3456), .Q(
        \inq_ary[9][132] ) );
  LATCHX1_RVT \inq_ary_reg[10][132]  ( .CLK(n3481), .D(n3456), .Q(
        \inq_ary[10][132] ) );
  LATCHX1_RVT \inq_ary_reg[11][132]  ( .CLK(n3480), .D(n3456), .Q(
        \inq_ary[11][132] ) );
  LATCHX1_RVT \inq_ary_reg[12][132]  ( .CLK(n3479), .D(n3456), .Q(
        \inq_ary[12][132] ) );
  LATCHX1_RVT \inq_ary_reg[13][132]  ( .CLK(n3478), .D(n3456), .Q(
        \inq_ary[13][132] ) );
  LATCHX1_RVT \inq_ary_reg[14][132]  ( .CLK(n3477), .D(n3456), .Q(
        \inq_ary[14][132] ) );
  LATCHX1_RVT \inq_ary_reg[15][132]  ( .CLK(n3476), .D(n3456), .Q(
        \inq_ary[15][132] ) );
  LATCHX1_RVT \dout_reg[132]  ( .CLK(n3492), .D(N394), .Q(dout[132]) );
  LATCHX1_RVT \inq_ary_reg[0][131]  ( .CLK(n3491), .D(n3463), .Q(
        \inq_ary[0][131] ) );
  LATCHX1_RVT \inq_ary_reg[1][131]  ( .CLK(n3490), .D(n3463), .Q(
        \inq_ary[1][131] ) );
  LATCHX1_RVT \inq_ary_reg[2][131]  ( .CLK(n3489), .D(n3463), .Q(
        \inq_ary[2][131] ) );
  LATCHX1_RVT \inq_ary_reg[3][131]  ( .CLK(n3488), .D(n3463), .Q(
        \inq_ary[3][131] ) );
  LATCHX1_RVT \inq_ary_reg[4][131]  ( .CLK(n3487), .D(n3463), .Q(
        \inq_ary[4][131] ) );
  LATCHX1_RVT \inq_ary_reg[5][131]  ( .CLK(n3486), .D(n3463), .Q(
        \inq_ary[5][131] ) );
  LATCHX1_RVT \inq_ary_reg[6][131]  ( .CLK(n3485), .D(n3463), .Q(
        \inq_ary[6][131] ) );
  LATCHX1_RVT \inq_ary_reg[7][131]  ( .CLK(n3484), .D(n3463), .Q(
        \inq_ary[7][131] ) );
  LATCHX1_RVT \inq_ary_reg[8][131]  ( .CLK(n3483), .D(n3463), .Q(
        \inq_ary[8][131] ) );
  LATCHX1_RVT \inq_ary_reg[9][131]  ( .CLK(n3482), .D(n3463), .Q(
        \inq_ary[9][131] ) );
  LATCHX1_RVT \inq_ary_reg[10][131]  ( .CLK(n3481), .D(n3463), .Q(
        \inq_ary[10][131] ) );
  LATCHX1_RVT \inq_ary_reg[11][131]  ( .CLK(n3480), .D(n3463), .Q(
        \inq_ary[11][131] ) );
  LATCHX1_RVT \inq_ary_reg[12][131]  ( .CLK(n3479), .D(n3463), .Q(
        \inq_ary[12][131] ) );
  LATCHX1_RVT \inq_ary_reg[13][131]  ( .CLK(n3478), .D(n3463), .Q(
        \inq_ary[13][131] ) );
  LATCHX1_RVT \inq_ary_reg[14][131]  ( .CLK(n3477), .D(n3463), .Q(
        \inq_ary[14][131] ) );
  LATCHX1_RVT \inq_ary_reg[15][131]  ( .CLK(n3476), .D(n3463), .Q(
        \inq_ary[15][131] ) );
  LATCHX1_RVT \dout_reg[131]  ( .CLK(n3492), .D(N393), .Q(dout[131]) );
  LATCHX1_RVT \inq_ary_reg[0][130]  ( .CLK(n3491), .D(n3461), .Q(
        \inq_ary[0][130] ) );
  LATCHX1_RVT \inq_ary_reg[1][130]  ( .CLK(n3490), .D(n3461), .Q(
        \inq_ary[1][130] ) );
  LATCHX1_RVT \inq_ary_reg[2][130]  ( .CLK(n3489), .D(n3461), .Q(
        \inq_ary[2][130] ) );
  LATCHX1_RVT \inq_ary_reg[3][130]  ( .CLK(n3488), .D(n3461), .Q(
        \inq_ary[3][130] ) );
  LATCHX1_RVT \inq_ary_reg[4][130]  ( .CLK(n3487), .D(n3461), .Q(
        \inq_ary[4][130] ) );
  LATCHX1_RVT \inq_ary_reg[5][130]  ( .CLK(n3486), .D(n3461), .Q(
        \inq_ary[5][130] ) );
  LATCHX1_RVT \inq_ary_reg[6][130]  ( .CLK(n3485), .D(n3461), .Q(
        \inq_ary[6][130] ) );
  LATCHX1_RVT \inq_ary_reg[7][130]  ( .CLK(n3484), .D(n3461), .Q(
        \inq_ary[7][130] ) );
  LATCHX1_RVT \inq_ary_reg[8][130]  ( .CLK(n3483), .D(n3461), .Q(
        \inq_ary[8][130] ) );
  LATCHX1_RVT \inq_ary_reg[9][130]  ( .CLK(n3482), .D(n3461), .Q(
        \inq_ary[9][130] ) );
  LATCHX1_RVT \inq_ary_reg[10][130]  ( .CLK(n3481), .D(n3461), .Q(
        \inq_ary[10][130] ) );
  LATCHX1_RVT \inq_ary_reg[11][130]  ( .CLK(n3480), .D(n3461), .Q(
        \inq_ary[11][130] ) );
  LATCHX1_RVT \inq_ary_reg[12][130]  ( .CLK(n3479), .D(n3461), .Q(
        \inq_ary[12][130] ) );
  LATCHX1_RVT \inq_ary_reg[13][130]  ( .CLK(n3478), .D(n3461), .Q(
        \inq_ary[13][130] ) );
  LATCHX1_RVT \inq_ary_reg[14][130]  ( .CLK(n3477), .D(n3461), .Q(
        \inq_ary[14][130] ) );
  LATCHX1_RVT \inq_ary_reg[15][130]  ( .CLK(n3476), .D(n3461), .Q(
        \inq_ary[15][130] ) );
  LATCHX1_RVT \dout_reg[130]  ( .CLK(n3492), .D(N392), .Q(dout[130]) );
  LATCHX1_RVT \inq_ary_reg[0][129]  ( .CLK(n3491), .D(n3459), .Q(
        \inq_ary[0][129] ) );
  LATCHX1_RVT \inq_ary_reg[1][129]  ( .CLK(n3490), .D(n3459), .Q(
        \inq_ary[1][129] ) );
  LATCHX1_RVT \inq_ary_reg[2][129]  ( .CLK(n3489), .D(n3459), .Q(
        \inq_ary[2][129] ) );
  LATCHX1_RVT \inq_ary_reg[3][129]  ( .CLK(n3488), .D(n3459), .Q(
        \inq_ary[3][129] ) );
  LATCHX1_RVT \inq_ary_reg[4][129]  ( .CLK(n3487), .D(n3459), .Q(
        \inq_ary[4][129] ) );
  LATCHX1_RVT \inq_ary_reg[5][129]  ( .CLK(n3486), .D(n3459), .Q(
        \inq_ary[5][129] ) );
  LATCHX1_RVT \inq_ary_reg[6][129]  ( .CLK(n3485), .D(n3459), .Q(
        \inq_ary[6][129] ) );
  LATCHX1_RVT \inq_ary_reg[7][129]  ( .CLK(n3484), .D(n3459), .Q(
        \inq_ary[7][129] ) );
  LATCHX1_RVT \inq_ary_reg[8][129]  ( .CLK(n3483), .D(n3459), .Q(
        \inq_ary[8][129] ) );
  LATCHX1_RVT \inq_ary_reg[9][129]  ( .CLK(n3482), .D(n3459), .Q(
        \inq_ary[9][129] ) );
  LATCHX1_RVT \inq_ary_reg[10][129]  ( .CLK(n3481), .D(n3459), .Q(
        \inq_ary[10][129] ) );
  LATCHX1_RVT \inq_ary_reg[11][129]  ( .CLK(n3480), .D(n3459), .Q(
        \inq_ary[11][129] ) );
  LATCHX1_RVT \inq_ary_reg[12][129]  ( .CLK(n3479), .D(n3459), .Q(
        \inq_ary[12][129] ) );
  LATCHX1_RVT \inq_ary_reg[13][129]  ( .CLK(n3478), .D(n3459), .Q(
        \inq_ary[13][129] ) );
  LATCHX1_RVT \inq_ary_reg[14][129]  ( .CLK(n3477), .D(n3459), .Q(
        \inq_ary[14][129] ) );
  LATCHX1_RVT \inq_ary_reg[15][129]  ( .CLK(n3476), .D(n3459), .Q(
        \inq_ary[15][129] ) );
  LATCHX1_RVT \dout_reg[129]  ( .CLK(n3492), .D(N391), .Q(dout[129]) );
  LATCHX1_RVT \inq_ary_reg[0][128]  ( .CLK(n3491), .D(n3457), .Q(
        \inq_ary[0][128] ) );
  LATCHX1_RVT \inq_ary_reg[1][128]  ( .CLK(n3490), .D(n3457), .Q(
        \inq_ary[1][128] ) );
  LATCHX1_RVT \inq_ary_reg[2][128]  ( .CLK(n3489), .D(n3457), .Q(
        \inq_ary[2][128] ) );
  LATCHX1_RVT \inq_ary_reg[3][128]  ( .CLK(n3488), .D(n3457), .Q(
        \inq_ary[3][128] ) );
  LATCHX1_RVT \inq_ary_reg[4][128]  ( .CLK(n3487), .D(n3457), .Q(
        \inq_ary[4][128] ) );
  LATCHX1_RVT \inq_ary_reg[5][128]  ( .CLK(n3486), .D(n3457), .Q(
        \inq_ary[5][128] ) );
  LATCHX1_RVT \inq_ary_reg[6][128]  ( .CLK(n3485), .D(n3457), .Q(
        \inq_ary[6][128] ) );
  LATCHX1_RVT \inq_ary_reg[7][128]  ( .CLK(n3484), .D(n3457), .Q(
        \inq_ary[7][128] ) );
  LATCHX1_RVT \inq_ary_reg[8][128]  ( .CLK(n3483), .D(n3457), .Q(
        \inq_ary[8][128] ) );
  LATCHX1_RVT \inq_ary_reg[9][128]  ( .CLK(n3482), .D(n3457), .Q(
        \inq_ary[9][128] ) );
  LATCHX1_RVT \inq_ary_reg[10][128]  ( .CLK(n3481), .D(n3457), .Q(
        \inq_ary[10][128] ) );
  LATCHX1_RVT \inq_ary_reg[11][128]  ( .CLK(n3480), .D(n3457), .Q(
        \inq_ary[11][128] ) );
  LATCHX1_RVT \inq_ary_reg[12][128]  ( .CLK(n3479), .D(n3457), .Q(
        \inq_ary[12][128] ) );
  LATCHX1_RVT \inq_ary_reg[13][128]  ( .CLK(n3478), .D(n3457), .Q(
        \inq_ary[13][128] ) );
  LATCHX1_RVT \inq_ary_reg[14][128]  ( .CLK(n3477), .D(n3457), .Q(
        \inq_ary[14][128] ) );
  LATCHX1_RVT \inq_ary_reg[15][128]  ( .CLK(n3476), .D(n3457), .Q(
        \inq_ary[15][128] ) );
  LATCHX1_RVT \dout_reg[128]  ( .CLK(n3492), .D(N390), .Q(dout[128]) );
  LATCHX1_RVT \inq_ary_reg[0][127]  ( .CLK(n3491), .D(n3454), .Q(
        \inq_ary[0][127] ) );
  LATCHX1_RVT \inq_ary_reg[1][127]  ( .CLK(n3490), .D(n3454), .Q(
        \inq_ary[1][127] ) );
  LATCHX1_RVT \inq_ary_reg[2][127]  ( .CLK(n3489), .D(n3454), .Q(
        \inq_ary[2][127] ) );
  LATCHX1_RVT \inq_ary_reg[3][127]  ( .CLK(n3488), .D(n3454), .Q(
        \inq_ary[3][127] ) );
  LATCHX1_RVT \inq_ary_reg[4][127]  ( .CLK(n3487), .D(n3454), .Q(
        \inq_ary[4][127] ) );
  LATCHX1_RVT \inq_ary_reg[5][127]  ( .CLK(n3486), .D(n3454), .Q(
        \inq_ary[5][127] ) );
  LATCHX1_RVT \inq_ary_reg[6][127]  ( .CLK(n3485), .D(n3454), .Q(
        \inq_ary[6][127] ) );
  LATCHX1_RVT \inq_ary_reg[7][127]  ( .CLK(n3484), .D(n3454), .Q(
        \inq_ary[7][127] ) );
  LATCHX1_RVT \inq_ary_reg[8][127]  ( .CLK(n3483), .D(n3454), .Q(
        \inq_ary[8][127] ) );
  LATCHX1_RVT \inq_ary_reg[9][127]  ( .CLK(n3482), .D(n3454), .Q(
        \inq_ary[9][127] ) );
  LATCHX1_RVT \inq_ary_reg[10][127]  ( .CLK(n3481), .D(n3454), .Q(
        \inq_ary[10][127] ) );
  LATCHX1_RVT \inq_ary_reg[11][127]  ( .CLK(n3480), .D(n3454), .Q(
        \inq_ary[11][127] ) );
  LATCHX1_RVT \inq_ary_reg[12][127]  ( .CLK(n3479), .D(n3454), .Q(
        \inq_ary[12][127] ) );
  LATCHX1_RVT \inq_ary_reg[13][127]  ( .CLK(n3478), .D(n3454), .Q(
        \inq_ary[13][127] ) );
  LATCHX1_RVT \inq_ary_reg[14][127]  ( .CLK(n3477), .D(n3454), .Q(
        \inq_ary[14][127] ) );
  LATCHX1_RVT \inq_ary_reg[15][127]  ( .CLK(n3476), .D(n3454), .Q(
        \inq_ary[15][127] ) );
  LATCHX1_RVT \dout_reg[127]  ( .CLK(n3492), .D(N389), .Q(dout[127]) );
  LATCHX1_RVT \inq_ary_reg[0][126]  ( .CLK(n3491), .D(n3452), .Q(
        \inq_ary[0][126] ) );
  LATCHX1_RVT \inq_ary_reg[1][126]  ( .CLK(n3490), .D(n3452), .Q(
        \inq_ary[1][126] ) );
  LATCHX1_RVT \inq_ary_reg[2][126]  ( .CLK(n3489), .D(n3452), .Q(
        \inq_ary[2][126] ) );
  LATCHX1_RVT \inq_ary_reg[3][126]  ( .CLK(n3488), .D(n3452), .Q(
        \inq_ary[3][126] ) );
  LATCHX1_RVT \inq_ary_reg[4][126]  ( .CLK(n3487), .D(n3452), .Q(
        \inq_ary[4][126] ) );
  LATCHX1_RVT \inq_ary_reg[5][126]  ( .CLK(n3486), .D(n3452), .Q(
        \inq_ary[5][126] ) );
  LATCHX1_RVT \inq_ary_reg[6][126]  ( .CLK(n3485), .D(n3452), .Q(
        \inq_ary[6][126] ) );
  LATCHX1_RVT \inq_ary_reg[7][126]  ( .CLK(n3484), .D(n3452), .Q(
        \inq_ary[7][126] ) );
  LATCHX1_RVT \inq_ary_reg[8][126]  ( .CLK(n3483), .D(n3452), .Q(
        \inq_ary[8][126] ) );
  LATCHX1_RVT \inq_ary_reg[9][126]  ( .CLK(n3482), .D(n3452), .Q(
        \inq_ary[9][126] ) );
  LATCHX1_RVT \inq_ary_reg[10][126]  ( .CLK(n3481), .D(n3452), .Q(
        \inq_ary[10][126] ) );
  LATCHX1_RVT \inq_ary_reg[11][126]  ( .CLK(n3480), .D(n3452), .Q(
        \inq_ary[11][126] ) );
  LATCHX1_RVT \inq_ary_reg[12][126]  ( .CLK(n3479), .D(n3452), .Q(
        \inq_ary[12][126] ) );
  LATCHX1_RVT \inq_ary_reg[13][126]  ( .CLK(n3478), .D(n3452), .Q(
        \inq_ary[13][126] ) );
  LATCHX1_RVT \inq_ary_reg[14][126]  ( .CLK(n3477), .D(n3452), .Q(
        \inq_ary[14][126] ) );
  LATCHX1_RVT \inq_ary_reg[15][126]  ( .CLK(n3476), .D(n3452), .Q(
        \inq_ary[15][126] ) );
  LATCHX1_RVT \dout_reg[126]  ( .CLK(n3492), .D(N388), .Q(dout[126]) );
  LATCHX1_RVT \inq_ary_reg[0][125]  ( .CLK(n3491), .D(n3450), .Q(
        \inq_ary[0][125] ) );
  LATCHX1_RVT \inq_ary_reg[1][125]  ( .CLK(n3490), .D(n3450), .Q(
        \inq_ary[1][125] ) );
  LATCHX1_RVT \inq_ary_reg[2][125]  ( .CLK(n3489), .D(n3450), .Q(
        \inq_ary[2][125] ) );
  LATCHX1_RVT \inq_ary_reg[3][125]  ( .CLK(n3488), .D(n3450), .Q(
        \inq_ary[3][125] ) );
  LATCHX1_RVT \inq_ary_reg[4][125]  ( .CLK(n3487), .D(n3450), .Q(
        \inq_ary[4][125] ) );
  LATCHX1_RVT \inq_ary_reg[5][125]  ( .CLK(n3486), .D(n3450), .Q(
        \inq_ary[5][125] ) );
  LATCHX1_RVT \inq_ary_reg[6][125]  ( .CLK(n3485), .D(n3450), .Q(
        \inq_ary[6][125] ) );
  LATCHX1_RVT \inq_ary_reg[7][125]  ( .CLK(n3484), .D(n3450), .Q(
        \inq_ary[7][125] ) );
  LATCHX1_RVT \inq_ary_reg[8][125]  ( .CLK(n3483), .D(n3450), .Q(
        \inq_ary[8][125] ) );
  LATCHX1_RVT \inq_ary_reg[9][125]  ( .CLK(n3482), .D(n3450), .Q(
        \inq_ary[9][125] ) );
  LATCHX1_RVT \inq_ary_reg[10][125]  ( .CLK(n3481), .D(n3450), .Q(
        \inq_ary[10][125] ) );
  LATCHX1_RVT \inq_ary_reg[11][125]  ( .CLK(n3480), .D(n3450), .Q(
        \inq_ary[11][125] ) );
  LATCHX1_RVT \inq_ary_reg[12][125]  ( .CLK(n3479), .D(n3450), .Q(
        \inq_ary[12][125] ) );
  LATCHX1_RVT \inq_ary_reg[13][125]  ( .CLK(n3478), .D(n3450), .Q(
        \inq_ary[13][125] ) );
  LATCHX1_RVT \inq_ary_reg[14][125]  ( .CLK(n3477), .D(n3450), .Q(
        \inq_ary[14][125] ) );
  LATCHX1_RVT \inq_ary_reg[15][125]  ( .CLK(n3476), .D(n3450), .Q(
        \inq_ary[15][125] ) );
  LATCHX1_RVT \dout_reg[125]  ( .CLK(n3492), .D(N387), .Q(dout[125]) );
  LATCHX1_RVT \inq_ary_reg[0][124]  ( .CLK(n3491), .D(n3448), .Q(
        \inq_ary[0][124] ) );
  LATCHX1_RVT \inq_ary_reg[1][124]  ( .CLK(n3490), .D(n3448), .Q(
        \inq_ary[1][124] ) );
  LATCHX1_RVT \inq_ary_reg[2][124]  ( .CLK(n3489), .D(n3448), .Q(
        \inq_ary[2][124] ) );
  LATCHX1_RVT \inq_ary_reg[3][124]  ( .CLK(n3488), .D(n3448), .Q(
        \inq_ary[3][124] ) );
  LATCHX1_RVT \inq_ary_reg[4][124]  ( .CLK(n3487), .D(n3448), .Q(
        \inq_ary[4][124] ) );
  LATCHX1_RVT \inq_ary_reg[5][124]  ( .CLK(n3486), .D(n3448), .Q(
        \inq_ary[5][124] ) );
  LATCHX1_RVT \inq_ary_reg[6][124]  ( .CLK(n3485), .D(n3448), .Q(
        \inq_ary[6][124] ) );
  LATCHX1_RVT \inq_ary_reg[7][124]  ( .CLK(n3484), .D(n3448), .Q(
        \inq_ary[7][124] ) );
  LATCHX1_RVT \inq_ary_reg[8][124]  ( .CLK(n3483), .D(n3448), .Q(
        \inq_ary[8][124] ) );
  LATCHX1_RVT \inq_ary_reg[9][124]  ( .CLK(n3482), .D(n3448), .Q(
        \inq_ary[9][124] ) );
  LATCHX1_RVT \inq_ary_reg[10][124]  ( .CLK(n3481), .D(n3448), .Q(
        \inq_ary[10][124] ) );
  LATCHX1_RVT \inq_ary_reg[11][124]  ( .CLK(n3480), .D(n3448), .Q(
        \inq_ary[11][124] ) );
  LATCHX1_RVT \inq_ary_reg[12][124]  ( .CLK(n3479), .D(n3448), .Q(
        \inq_ary[12][124] ) );
  LATCHX1_RVT \inq_ary_reg[13][124]  ( .CLK(n3478), .D(n3448), .Q(
        \inq_ary[13][124] ) );
  LATCHX1_RVT \inq_ary_reg[14][124]  ( .CLK(n3477), .D(n3448), .Q(
        \inq_ary[14][124] ) );
  LATCHX1_RVT \inq_ary_reg[15][124]  ( .CLK(n3476), .D(n3448), .Q(
        \inq_ary[15][124] ) );
  LATCHX1_RVT \dout_reg[124]  ( .CLK(n3492), .D(N386), .Q(dout[124]) );
  LATCHX1_RVT \inq_ary_reg[0][123]  ( .CLK(n3491), .D(n3455), .Q(
        \inq_ary[0][123] ) );
  LATCHX1_RVT \inq_ary_reg[1][123]  ( .CLK(n3490), .D(n3455), .Q(
        \inq_ary[1][123] ) );
  LATCHX1_RVT \inq_ary_reg[2][123]  ( .CLK(n3489), .D(n3455), .Q(
        \inq_ary[2][123] ) );
  LATCHX1_RVT \inq_ary_reg[3][123]  ( .CLK(n3488), .D(n3455), .Q(
        \inq_ary[3][123] ) );
  LATCHX1_RVT \inq_ary_reg[4][123]  ( .CLK(n3487), .D(n3455), .Q(
        \inq_ary[4][123] ) );
  LATCHX1_RVT \inq_ary_reg[5][123]  ( .CLK(n3486), .D(n3455), .Q(
        \inq_ary[5][123] ) );
  LATCHX1_RVT \inq_ary_reg[6][123]  ( .CLK(n3485), .D(n3455), .Q(
        \inq_ary[6][123] ) );
  LATCHX1_RVT \inq_ary_reg[7][123]  ( .CLK(n3484), .D(n3455), .Q(
        \inq_ary[7][123] ) );
  LATCHX1_RVT \inq_ary_reg[8][123]  ( .CLK(n3483), .D(n3455), .Q(
        \inq_ary[8][123] ) );
  LATCHX1_RVT \inq_ary_reg[9][123]  ( .CLK(n3482), .D(n3455), .Q(
        \inq_ary[9][123] ) );
  LATCHX1_RVT \inq_ary_reg[10][123]  ( .CLK(n3481), .D(n3455), .Q(
        \inq_ary[10][123] ) );
  LATCHX1_RVT \inq_ary_reg[11][123]  ( .CLK(n3480), .D(n3455), .Q(
        \inq_ary[11][123] ) );
  LATCHX1_RVT \inq_ary_reg[12][123]  ( .CLK(n3479), .D(n3455), .Q(
        \inq_ary[12][123] ) );
  LATCHX1_RVT \inq_ary_reg[13][123]  ( .CLK(n3478), .D(n3455), .Q(
        \inq_ary[13][123] ) );
  LATCHX1_RVT \inq_ary_reg[14][123]  ( .CLK(n3477), .D(n3455), .Q(
        \inq_ary[14][123] ) );
  LATCHX1_RVT \inq_ary_reg[15][123]  ( .CLK(n3476), .D(n3455), .Q(
        \inq_ary[15][123] ) );
  LATCHX1_RVT \dout_reg[123]  ( .CLK(n3492), .D(N385), .Q(dout[123]) );
  LATCHX1_RVT \inq_ary_reg[0][122]  ( .CLK(n3491), .D(n3453), .Q(
        \inq_ary[0][122] ) );
  LATCHX1_RVT \inq_ary_reg[1][122]  ( .CLK(n3490), .D(n3453), .Q(
        \inq_ary[1][122] ) );
  LATCHX1_RVT \inq_ary_reg[2][122]  ( .CLK(n3489), .D(n3453), .Q(
        \inq_ary[2][122] ) );
  LATCHX1_RVT \inq_ary_reg[3][122]  ( .CLK(n3488), .D(n3453), .Q(
        \inq_ary[3][122] ) );
  LATCHX1_RVT \inq_ary_reg[4][122]  ( .CLK(n3487), .D(n3453), .Q(
        \inq_ary[4][122] ) );
  LATCHX1_RVT \inq_ary_reg[5][122]  ( .CLK(n3486), .D(n3453), .Q(
        \inq_ary[5][122] ) );
  LATCHX1_RVT \inq_ary_reg[6][122]  ( .CLK(n3485), .D(n3453), .Q(
        \inq_ary[6][122] ) );
  LATCHX1_RVT \inq_ary_reg[7][122]  ( .CLK(n3484), .D(n3453), .Q(
        \inq_ary[7][122] ) );
  LATCHX1_RVT \inq_ary_reg[8][122]  ( .CLK(n3483), .D(n3453), .Q(
        \inq_ary[8][122] ) );
  LATCHX1_RVT \inq_ary_reg[9][122]  ( .CLK(n3482), .D(n3453), .Q(
        \inq_ary[9][122] ) );
  LATCHX1_RVT \inq_ary_reg[10][122]  ( .CLK(n3481), .D(n3453), .Q(
        \inq_ary[10][122] ) );
  LATCHX1_RVT \inq_ary_reg[11][122]  ( .CLK(n3480), .D(n3453), .Q(
        \inq_ary[11][122] ) );
  LATCHX1_RVT \inq_ary_reg[12][122]  ( .CLK(n3479), .D(n3453), .Q(
        \inq_ary[12][122] ) );
  LATCHX1_RVT \inq_ary_reg[13][122]  ( .CLK(n3478), .D(n3453), .Q(
        \inq_ary[13][122] ) );
  LATCHX1_RVT \inq_ary_reg[14][122]  ( .CLK(n3477), .D(n3453), .Q(
        \inq_ary[14][122] ) );
  LATCHX1_RVT \inq_ary_reg[15][122]  ( .CLK(n3476), .D(n3453), .Q(
        \inq_ary[15][122] ) );
  LATCHX1_RVT \dout_reg[122]  ( .CLK(n3492), .D(N384), .Q(dout[122]) );
  LATCHX1_RVT \inq_ary_reg[0][121]  ( .CLK(n3491), .D(n3451), .Q(
        \inq_ary[0][121] ) );
  LATCHX1_RVT \inq_ary_reg[1][121]  ( .CLK(n3490), .D(n3451), .Q(
        \inq_ary[1][121] ) );
  LATCHX1_RVT \inq_ary_reg[2][121]  ( .CLK(n3489), .D(n3451), .Q(
        \inq_ary[2][121] ) );
  LATCHX1_RVT \inq_ary_reg[3][121]  ( .CLK(n3488), .D(n3451), .Q(
        \inq_ary[3][121] ) );
  LATCHX1_RVT \inq_ary_reg[4][121]  ( .CLK(n3487), .D(n3451), .Q(
        \inq_ary[4][121] ) );
  LATCHX1_RVT \inq_ary_reg[5][121]  ( .CLK(n3486), .D(n3451), .Q(
        \inq_ary[5][121] ) );
  LATCHX1_RVT \inq_ary_reg[6][121]  ( .CLK(n3485), .D(n3451), .Q(
        \inq_ary[6][121] ) );
  LATCHX1_RVT \inq_ary_reg[7][121]  ( .CLK(n3484), .D(n3451), .Q(
        \inq_ary[7][121] ) );
  LATCHX1_RVT \inq_ary_reg[8][121]  ( .CLK(n3483), .D(n3451), .Q(
        \inq_ary[8][121] ) );
  LATCHX1_RVT \inq_ary_reg[9][121]  ( .CLK(n3482), .D(n3451), .Q(
        \inq_ary[9][121] ) );
  LATCHX1_RVT \inq_ary_reg[10][121]  ( .CLK(n3481), .D(n3451), .Q(
        \inq_ary[10][121] ) );
  LATCHX1_RVT \inq_ary_reg[11][121]  ( .CLK(n3480), .D(n3451), .Q(
        \inq_ary[11][121] ) );
  LATCHX1_RVT \inq_ary_reg[12][121]  ( .CLK(n3479), .D(n3451), .Q(
        \inq_ary[12][121] ) );
  LATCHX1_RVT \inq_ary_reg[13][121]  ( .CLK(n3478), .D(n3451), .Q(
        \inq_ary[13][121] ) );
  LATCHX1_RVT \inq_ary_reg[14][121]  ( .CLK(n3477), .D(n3451), .Q(
        \inq_ary[14][121] ) );
  LATCHX1_RVT \inq_ary_reg[15][121]  ( .CLK(n3476), .D(n3451), .Q(
        \inq_ary[15][121] ) );
  LATCHX1_RVT \dout_reg[121]  ( .CLK(n3492), .D(N383), .Q(dout[121]) );
  LATCHX1_RVT \inq_ary_reg[0][120]  ( .CLK(n3491), .D(n3449), .Q(
        \inq_ary[0][120] ) );
  LATCHX1_RVT \inq_ary_reg[1][120]  ( .CLK(n3490), .D(n3449), .Q(
        \inq_ary[1][120] ) );
  LATCHX1_RVT \inq_ary_reg[2][120]  ( .CLK(n3489), .D(n3449), .Q(
        \inq_ary[2][120] ) );
  LATCHX1_RVT \inq_ary_reg[3][120]  ( .CLK(n3488), .D(n3449), .Q(
        \inq_ary[3][120] ) );
  LATCHX1_RVT \inq_ary_reg[4][120]  ( .CLK(n3487), .D(n3449), .Q(
        \inq_ary[4][120] ) );
  LATCHX1_RVT \inq_ary_reg[5][120]  ( .CLK(n3486), .D(n3449), .Q(
        \inq_ary[5][120] ) );
  LATCHX1_RVT \inq_ary_reg[6][120]  ( .CLK(n3485), .D(n3449), .Q(
        \inq_ary[6][120] ) );
  LATCHX1_RVT \inq_ary_reg[7][120]  ( .CLK(n3484), .D(n3449), .Q(
        \inq_ary[7][120] ) );
  LATCHX1_RVT \inq_ary_reg[8][120]  ( .CLK(n3483), .D(n3449), .Q(
        \inq_ary[8][120] ) );
  LATCHX1_RVT \inq_ary_reg[9][120]  ( .CLK(n3482), .D(n3449), .Q(
        \inq_ary[9][120] ) );
  LATCHX1_RVT \inq_ary_reg[10][120]  ( .CLK(n3481), .D(n3449), .Q(
        \inq_ary[10][120] ) );
  LATCHX1_RVT \inq_ary_reg[11][120]  ( .CLK(n3480), .D(n3449), .Q(
        \inq_ary[11][120] ) );
  LATCHX1_RVT \inq_ary_reg[12][120]  ( .CLK(n3479), .D(n3449), .Q(
        \inq_ary[12][120] ) );
  LATCHX1_RVT \inq_ary_reg[13][120]  ( .CLK(n3478), .D(n3449), .Q(
        \inq_ary[13][120] ) );
  LATCHX1_RVT \inq_ary_reg[14][120]  ( .CLK(n3477), .D(n3449), .Q(
        \inq_ary[14][120] ) );
  LATCHX1_RVT \inq_ary_reg[15][120]  ( .CLK(n3476), .D(n3449), .Q(
        \inq_ary[15][120] ) );
  LATCHX1_RVT \dout_reg[120]  ( .CLK(n3492), .D(N382), .Q(dout[120]) );
  LATCHX1_RVT \inq_ary_reg[0][119]  ( .CLK(n3491), .D(n3446), .Q(
        \inq_ary[0][119] ) );
  LATCHX1_RVT \inq_ary_reg[1][119]  ( .CLK(n3490), .D(n3446), .Q(
        \inq_ary[1][119] ) );
  LATCHX1_RVT \inq_ary_reg[2][119]  ( .CLK(n3489), .D(n3446), .Q(
        \inq_ary[2][119] ) );
  LATCHX1_RVT \inq_ary_reg[3][119]  ( .CLK(n3488), .D(n3446), .Q(
        \inq_ary[3][119] ) );
  LATCHX1_RVT \inq_ary_reg[4][119]  ( .CLK(n3487), .D(n3446), .Q(
        \inq_ary[4][119] ) );
  LATCHX1_RVT \inq_ary_reg[5][119]  ( .CLK(n3486), .D(n3446), .Q(
        \inq_ary[5][119] ) );
  LATCHX1_RVT \inq_ary_reg[6][119]  ( .CLK(n3485), .D(n3446), .Q(
        \inq_ary[6][119] ) );
  LATCHX1_RVT \inq_ary_reg[7][119]  ( .CLK(n3484), .D(n3446), .Q(
        \inq_ary[7][119] ) );
  LATCHX1_RVT \inq_ary_reg[8][119]  ( .CLK(n3483), .D(n3446), .Q(
        \inq_ary[8][119] ) );
  LATCHX1_RVT \inq_ary_reg[9][119]  ( .CLK(n3482), .D(n3446), .Q(
        \inq_ary[9][119] ) );
  LATCHX1_RVT \inq_ary_reg[10][119]  ( .CLK(n3481), .D(n3446), .Q(
        \inq_ary[10][119] ) );
  LATCHX1_RVT \inq_ary_reg[11][119]  ( .CLK(n3480), .D(n3446), .Q(
        \inq_ary[11][119] ) );
  LATCHX1_RVT \inq_ary_reg[12][119]  ( .CLK(n3479), .D(n3446), .Q(
        \inq_ary[12][119] ) );
  LATCHX1_RVT \inq_ary_reg[13][119]  ( .CLK(n3478), .D(n3446), .Q(
        \inq_ary[13][119] ) );
  LATCHX1_RVT \inq_ary_reg[14][119]  ( .CLK(n3477), .D(n3446), .Q(
        \inq_ary[14][119] ) );
  LATCHX1_RVT \inq_ary_reg[15][119]  ( .CLK(n3476), .D(n3446), .Q(
        \inq_ary[15][119] ) );
  LATCHX1_RVT \dout_reg[119]  ( .CLK(n3492), .D(N381), .Q(dout[119]) );
  LATCHX1_RVT \inq_ary_reg[0][118]  ( .CLK(n3491), .D(n3444), .Q(
        \inq_ary[0][118] ) );
  LATCHX1_RVT \inq_ary_reg[1][118]  ( .CLK(n3490), .D(n3444), .Q(
        \inq_ary[1][118] ) );
  LATCHX1_RVT \inq_ary_reg[2][118]  ( .CLK(n3489), .D(n3444), .Q(
        \inq_ary[2][118] ) );
  LATCHX1_RVT \inq_ary_reg[3][118]  ( .CLK(n3488), .D(n3444), .Q(
        \inq_ary[3][118] ) );
  LATCHX1_RVT \inq_ary_reg[4][118]  ( .CLK(n3487), .D(n3444), .Q(
        \inq_ary[4][118] ) );
  LATCHX1_RVT \inq_ary_reg[5][118]  ( .CLK(n3486), .D(n3444), .Q(
        \inq_ary[5][118] ) );
  LATCHX1_RVT \inq_ary_reg[6][118]  ( .CLK(n3485), .D(n3444), .Q(
        \inq_ary[6][118] ) );
  LATCHX1_RVT \inq_ary_reg[7][118]  ( .CLK(n3484), .D(n3444), .Q(
        \inq_ary[7][118] ) );
  LATCHX1_RVT \inq_ary_reg[8][118]  ( .CLK(n3483), .D(n3444), .Q(
        \inq_ary[8][118] ) );
  LATCHX1_RVT \inq_ary_reg[9][118]  ( .CLK(n3482), .D(n3444), .Q(
        \inq_ary[9][118] ) );
  LATCHX1_RVT \inq_ary_reg[10][118]  ( .CLK(n3481), .D(n3444), .Q(
        \inq_ary[10][118] ) );
  LATCHX1_RVT \inq_ary_reg[11][118]  ( .CLK(n3480), .D(n3444), .Q(
        \inq_ary[11][118] ) );
  LATCHX1_RVT \inq_ary_reg[12][118]  ( .CLK(n3479), .D(n3444), .Q(
        \inq_ary[12][118] ) );
  LATCHX1_RVT \inq_ary_reg[13][118]  ( .CLK(n3478), .D(n3444), .Q(
        \inq_ary[13][118] ) );
  LATCHX1_RVT \inq_ary_reg[14][118]  ( .CLK(n3477), .D(n3444), .Q(
        \inq_ary[14][118] ) );
  LATCHX1_RVT \inq_ary_reg[15][118]  ( .CLK(n3476), .D(n3444), .Q(
        \inq_ary[15][118] ) );
  LATCHX1_RVT \dout_reg[118]  ( .CLK(n3492), .D(N380), .Q(dout[118]) );
  LATCHX1_RVT \inq_ary_reg[0][117]  ( .CLK(n3491), .D(n3442), .Q(
        \inq_ary[0][117] ) );
  LATCHX1_RVT \inq_ary_reg[1][117]  ( .CLK(n3490), .D(n3442), .Q(
        \inq_ary[1][117] ) );
  LATCHX1_RVT \inq_ary_reg[2][117]  ( .CLK(n3489), .D(n3442), .Q(
        \inq_ary[2][117] ) );
  LATCHX1_RVT \inq_ary_reg[3][117]  ( .CLK(n3488), .D(n3442), .Q(
        \inq_ary[3][117] ) );
  LATCHX1_RVT \inq_ary_reg[4][117]  ( .CLK(n3487), .D(n3442), .Q(
        \inq_ary[4][117] ) );
  LATCHX1_RVT \inq_ary_reg[5][117]  ( .CLK(n3486), .D(n3442), .Q(
        \inq_ary[5][117] ) );
  LATCHX1_RVT \inq_ary_reg[6][117]  ( .CLK(n3485), .D(n3442), .Q(
        \inq_ary[6][117] ) );
  LATCHX1_RVT \inq_ary_reg[7][117]  ( .CLK(n3484), .D(n3442), .Q(
        \inq_ary[7][117] ) );
  LATCHX1_RVT \inq_ary_reg[8][117]  ( .CLK(n3483), .D(n3442), .Q(
        \inq_ary[8][117] ) );
  LATCHX1_RVT \inq_ary_reg[9][117]  ( .CLK(n3482), .D(n3442), .Q(
        \inq_ary[9][117] ) );
  LATCHX1_RVT \inq_ary_reg[10][117]  ( .CLK(n3481), .D(n3442), .Q(
        \inq_ary[10][117] ) );
  LATCHX1_RVT \inq_ary_reg[11][117]  ( .CLK(n3480), .D(n3442), .Q(
        \inq_ary[11][117] ) );
  LATCHX1_RVT \inq_ary_reg[12][117]  ( .CLK(n3479), .D(n3442), .Q(
        \inq_ary[12][117] ) );
  LATCHX1_RVT \inq_ary_reg[13][117]  ( .CLK(n3478), .D(n3442), .Q(
        \inq_ary[13][117] ) );
  LATCHX1_RVT \inq_ary_reg[14][117]  ( .CLK(n3477), .D(n3442), .Q(
        \inq_ary[14][117] ) );
  LATCHX1_RVT \inq_ary_reg[15][117]  ( .CLK(n3476), .D(n3442), .Q(
        \inq_ary[15][117] ) );
  LATCHX1_RVT \dout_reg[117]  ( .CLK(n3492), .D(N379), .Q(dout[117]) );
  LATCHX1_RVT \inq_ary_reg[0][116]  ( .CLK(n3491), .D(n3440), .Q(
        \inq_ary[0][116] ) );
  LATCHX1_RVT \inq_ary_reg[1][116]  ( .CLK(n3490), .D(n3440), .Q(
        \inq_ary[1][116] ) );
  LATCHX1_RVT \inq_ary_reg[2][116]  ( .CLK(n3489), .D(n3440), .Q(
        \inq_ary[2][116] ) );
  LATCHX1_RVT \inq_ary_reg[3][116]  ( .CLK(n3488), .D(n3440), .Q(
        \inq_ary[3][116] ) );
  LATCHX1_RVT \inq_ary_reg[4][116]  ( .CLK(n3487), .D(n3440), .Q(
        \inq_ary[4][116] ) );
  LATCHX1_RVT \inq_ary_reg[5][116]  ( .CLK(n3486), .D(n3440), .Q(
        \inq_ary[5][116] ) );
  LATCHX1_RVT \inq_ary_reg[6][116]  ( .CLK(n3485), .D(n3440), .Q(
        \inq_ary[6][116] ) );
  LATCHX1_RVT \inq_ary_reg[7][116]  ( .CLK(n3484), .D(n3440), .Q(
        \inq_ary[7][116] ) );
  LATCHX1_RVT \inq_ary_reg[8][116]  ( .CLK(n3483), .D(n3440), .Q(
        \inq_ary[8][116] ) );
  LATCHX1_RVT \inq_ary_reg[9][116]  ( .CLK(n3482), .D(n3440), .Q(
        \inq_ary[9][116] ) );
  LATCHX1_RVT \inq_ary_reg[10][116]  ( .CLK(n3481), .D(n3440), .Q(
        \inq_ary[10][116] ) );
  LATCHX1_RVT \inq_ary_reg[11][116]  ( .CLK(n3480), .D(n3440), .Q(
        \inq_ary[11][116] ) );
  LATCHX1_RVT \inq_ary_reg[12][116]  ( .CLK(n3479), .D(n3440), .Q(
        \inq_ary[12][116] ) );
  LATCHX1_RVT \inq_ary_reg[13][116]  ( .CLK(n3478), .D(n3440), .Q(
        \inq_ary[13][116] ) );
  LATCHX1_RVT \inq_ary_reg[14][116]  ( .CLK(n3477), .D(n3440), .Q(
        \inq_ary[14][116] ) );
  LATCHX1_RVT \inq_ary_reg[15][116]  ( .CLK(n3476), .D(n3440), .Q(
        \inq_ary[15][116] ) );
  LATCHX1_RVT \dout_reg[116]  ( .CLK(n3492), .D(N378), .Q(dout[116]) );
  LATCHX1_RVT \inq_ary_reg[0][115]  ( .CLK(n3491), .D(n3447), .Q(
        \inq_ary[0][115] ) );
  LATCHX1_RVT \inq_ary_reg[1][115]  ( .CLK(n3490), .D(n3447), .Q(
        \inq_ary[1][115] ) );
  LATCHX1_RVT \inq_ary_reg[2][115]  ( .CLK(n3489), .D(n3447), .Q(
        \inq_ary[2][115] ) );
  LATCHX1_RVT \inq_ary_reg[3][115]  ( .CLK(n3488), .D(n3447), .Q(
        \inq_ary[3][115] ) );
  LATCHX1_RVT \inq_ary_reg[4][115]  ( .CLK(n3487), .D(n3447), .Q(
        \inq_ary[4][115] ) );
  LATCHX1_RVT \inq_ary_reg[5][115]  ( .CLK(n3486), .D(n3447), .Q(
        \inq_ary[5][115] ) );
  LATCHX1_RVT \inq_ary_reg[6][115]  ( .CLK(n3485), .D(n3447), .Q(
        \inq_ary[6][115] ) );
  LATCHX1_RVT \inq_ary_reg[7][115]  ( .CLK(n3484), .D(n3447), .Q(
        \inq_ary[7][115] ) );
  LATCHX1_RVT \inq_ary_reg[8][115]  ( .CLK(n3483), .D(n3447), .Q(
        \inq_ary[8][115] ) );
  LATCHX1_RVT \inq_ary_reg[9][115]  ( .CLK(n3482), .D(n3447), .Q(
        \inq_ary[9][115] ) );
  LATCHX1_RVT \inq_ary_reg[10][115]  ( .CLK(n3481), .D(n3447), .Q(
        \inq_ary[10][115] ) );
  LATCHX1_RVT \inq_ary_reg[11][115]  ( .CLK(n3480), .D(n3447), .Q(
        \inq_ary[11][115] ) );
  LATCHX1_RVT \inq_ary_reg[12][115]  ( .CLK(n3479), .D(n3447), .Q(
        \inq_ary[12][115] ) );
  LATCHX1_RVT \inq_ary_reg[13][115]  ( .CLK(n3478), .D(n3447), .Q(
        \inq_ary[13][115] ) );
  LATCHX1_RVT \inq_ary_reg[14][115]  ( .CLK(n3477), .D(n3447), .Q(
        \inq_ary[14][115] ) );
  LATCHX1_RVT \inq_ary_reg[15][115]  ( .CLK(n3476), .D(n3447), .Q(
        \inq_ary[15][115] ) );
  LATCHX1_RVT \dout_reg[115]  ( .CLK(n3492), .D(N377), .Q(dout[115]) );
  LATCHX1_RVT \inq_ary_reg[0][114]  ( .CLK(n3491), .D(n3445), .Q(
        \inq_ary[0][114] ) );
  LATCHX1_RVT \inq_ary_reg[1][114]  ( .CLK(n3490), .D(n3445), .Q(
        \inq_ary[1][114] ) );
  LATCHX1_RVT \inq_ary_reg[2][114]  ( .CLK(n3489), .D(n3445), .Q(
        \inq_ary[2][114] ) );
  LATCHX1_RVT \inq_ary_reg[3][114]  ( .CLK(n3488), .D(n3445), .Q(
        \inq_ary[3][114] ) );
  LATCHX1_RVT \inq_ary_reg[4][114]  ( .CLK(n3487), .D(n3445), .Q(
        \inq_ary[4][114] ) );
  LATCHX1_RVT \inq_ary_reg[5][114]  ( .CLK(n3486), .D(n3445), .Q(
        \inq_ary[5][114] ) );
  LATCHX1_RVT \inq_ary_reg[6][114]  ( .CLK(n3485), .D(n3445), .Q(
        \inq_ary[6][114] ) );
  LATCHX1_RVT \inq_ary_reg[7][114]  ( .CLK(n3484), .D(n3445), .Q(
        \inq_ary[7][114] ) );
  LATCHX1_RVT \inq_ary_reg[8][114]  ( .CLK(n3483), .D(n3445), .Q(
        \inq_ary[8][114] ) );
  LATCHX1_RVT \inq_ary_reg[9][114]  ( .CLK(n3482), .D(n3445), .Q(
        \inq_ary[9][114] ) );
  LATCHX1_RVT \inq_ary_reg[10][114]  ( .CLK(n3481), .D(n3445), .Q(
        \inq_ary[10][114] ) );
  LATCHX1_RVT \inq_ary_reg[11][114]  ( .CLK(n3480), .D(n3445), .Q(
        \inq_ary[11][114] ) );
  LATCHX1_RVT \inq_ary_reg[12][114]  ( .CLK(n3479), .D(n3445), .Q(
        \inq_ary[12][114] ) );
  LATCHX1_RVT \inq_ary_reg[13][114]  ( .CLK(n3478), .D(n3445), .Q(
        \inq_ary[13][114] ) );
  LATCHX1_RVT \inq_ary_reg[14][114]  ( .CLK(n3477), .D(n3445), .Q(
        \inq_ary[14][114] ) );
  LATCHX1_RVT \inq_ary_reg[15][114]  ( .CLK(n3476), .D(n3445), .Q(
        \inq_ary[15][114] ) );
  LATCHX1_RVT \dout_reg[114]  ( .CLK(n3492), .D(N376), .Q(dout[114]) );
  LATCHX1_RVT \inq_ary_reg[0][113]  ( .CLK(n3491), .D(n3443), .Q(
        \inq_ary[0][113] ) );
  LATCHX1_RVT \inq_ary_reg[1][113]  ( .CLK(n3490), .D(n3443), .Q(
        \inq_ary[1][113] ) );
  LATCHX1_RVT \inq_ary_reg[2][113]  ( .CLK(n3489), .D(n3443), .Q(
        \inq_ary[2][113] ) );
  LATCHX1_RVT \inq_ary_reg[3][113]  ( .CLK(n3488), .D(n3443), .Q(
        \inq_ary[3][113] ) );
  LATCHX1_RVT \inq_ary_reg[4][113]  ( .CLK(n3487), .D(n3443), .Q(
        \inq_ary[4][113] ) );
  LATCHX1_RVT \inq_ary_reg[5][113]  ( .CLK(n3486), .D(n3443), .Q(
        \inq_ary[5][113] ) );
  LATCHX1_RVT \inq_ary_reg[6][113]  ( .CLK(n3485), .D(n3443), .Q(
        \inq_ary[6][113] ) );
  LATCHX1_RVT \inq_ary_reg[7][113]  ( .CLK(n3484), .D(n3443), .Q(
        \inq_ary[7][113] ) );
  LATCHX1_RVT \inq_ary_reg[8][113]  ( .CLK(n3483), .D(n3443), .Q(
        \inq_ary[8][113] ) );
  LATCHX1_RVT \inq_ary_reg[9][113]  ( .CLK(n3482), .D(n3443), .Q(
        \inq_ary[9][113] ) );
  LATCHX1_RVT \inq_ary_reg[10][113]  ( .CLK(n3481), .D(n3443), .Q(
        \inq_ary[10][113] ) );
  LATCHX1_RVT \inq_ary_reg[11][113]  ( .CLK(n3480), .D(n3443), .Q(
        \inq_ary[11][113] ) );
  LATCHX1_RVT \inq_ary_reg[12][113]  ( .CLK(n3479), .D(n3443), .Q(
        \inq_ary[12][113] ) );
  LATCHX1_RVT \inq_ary_reg[13][113]  ( .CLK(n3478), .D(n3443), .Q(
        \inq_ary[13][113] ) );
  LATCHX1_RVT \inq_ary_reg[14][113]  ( .CLK(n3477), .D(n3443), .Q(
        \inq_ary[14][113] ) );
  LATCHX1_RVT \inq_ary_reg[15][113]  ( .CLK(n3476), .D(n3443), .Q(
        \inq_ary[15][113] ) );
  LATCHX1_RVT \dout_reg[113]  ( .CLK(n3492), .D(N375), .Q(dout[113]) );
  LATCHX1_RVT \inq_ary_reg[0][112]  ( .CLK(n3491), .D(n3441), .Q(
        \inq_ary[0][112] ) );
  LATCHX1_RVT \inq_ary_reg[1][112]  ( .CLK(n3490), .D(n3441), .Q(
        \inq_ary[1][112] ) );
  LATCHX1_RVT \inq_ary_reg[2][112]  ( .CLK(n3489), .D(n3441), .Q(
        \inq_ary[2][112] ) );
  LATCHX1_RVT \inq_ary_reg[3][112]  ( .CLK(n3488), .D(n3441), .Q(
        \inq_ary[3][112] ) );
  LATCHX1_RVT \inq_ary_reg[4][112]  ( .CLK(n3487), .D(n3441), .Q(
        \inq_ary[4][112] ) );
  LATCHX1_RVT \inq_ary_reg[5][112]  ( .CLK(n3486), .D(n3441), .Q(
        \inq_ary[5][112] ) );
  LATCHX1_RVT \inq_ary_reg[6][112]  ( .CLK(n3485), .D(n3441), .Q(
        \inq_ary[6][112] ) );
  LATCHX1_RVT \inq_ary_reg[7][112]  ( .CLK(n3484), .D(n3441), .Q(
        \inq_ary[7][112] ) );
  LATCHX1_RVT \inq_ary_reg[8][112]  ( .CLK(n3483), .D(n3441), .Q(
        \inq_ary[8][112] ) );
  LATCHX1_RVT \inq_ary_reg[9][112]  ( .CLK(n3482), .D(n3441), .Q(
        \inq_ary[9][112] ) );
  LATCHX1_RVT \inq_ary_reg[10][112]  ( .CLK(n3481), .D(n3441), .Q(
        \inq_ary[10][112] ) );
  LATCHX1_RVT \inq_ary_reg[11][112]  ( .CLK(n3480), .D(n3441), .Q(
        \inq_ary[11][112] ) );
  LATCHX1_RVT \inq_ary_reg[12][112]  ( .CLK(n3479), .D(n3441), .Q(
        \inq_ary[12][112] ) );
  LATCHX1_RVT \inq_ary_reg[13][112]  ( .CLK(n3478), .D(n3441), .Q(
        \inq_ary[13][112] ) );
  LATCHX1_RVT \inq_ary_reg[14][112]  ( .CLK(n3477), .D(n3441), .Q(
        \inq_ary[14][112] ) );
  LATCHX1_RVT \inq_ary_reg[15][112]  ( .CLK(n3476), .D(n3441), .Q(
        \inq_ary[15][112] ) );
  LATCHX1_RVT \dout_reg[112]  ( .CLK(n3492), .D(N374), .Q(dout[112]) );
  LATCHX1_RVT \inq_ary_reg[0][111]  ( .CLK(n3491), .D(n3438), .Q(
        \inq_ary[0][111] ) );
  LATCHX1_RVT \inq_ary_reg[1][111]  ( .CLK(n3490), .D(n3438), .Q(
        \inq_ary[1][111] ) );
  LATCHX1_RVT \inq_ary_reg[2][111]  ( .CLK(n3489), .D(n3438), .Q(
        \inq_ary[2][111] ) );
  LATCHX1_RVT \inq_ary_reg[3][111]  ( .CLK(n3488), .D(n3438), .Q(
        \inq_ary[3][111] ) );
  LATCHX1_RVT \inq_ary_reg[4][111]  ( .CLK(n3487), .D(n3438), .Q(
        \inq_ary[4][111] ) );
  LATCHX1_RVT \inq_ary_reg[5][111]  ( .CLK(n3486), .D(n3438), .Q(
        \inq_ary[5][111] ) );
  LATCHX1_RVT \inq_ary_reg[6][111]  ( .CLK(n3485), .D(n3438), .Q(
        \inq_ary[6][111] ) );
  LATCHX1_RVT \inq_ary_reg[7][111]  ( .CLK(n3484), .D(n3438), .Q(
        \inq_ary[7][111] ) );
  LATCHX1_RVT \inq_ary_reg[8][111]  ( .CLK(n3483), .D(n3438), .Q(
        \inq_ary[8][111] ) );
  LATCHX1_RVT \inq_ary_reg[9][111]  ( .CLK(n3482), .D(n3438), .Q(
        \inq_ary[9][111] ) );
  LATCHX1_RVT \inq_ary_reg[10][111]  ( .CLK(n3481), .D(n3438), .Q(
        \inq_ary[10][111] ) );
  LATCHX1_RVT \inq_ary_reg[11][111]  ( .CLK(n3480), .D(n3438), .Q(
        \inq_ary[11][111] ) );
  LATCHX1_RVT \inq_ary_reg[12][111]  ( .CLK(n3479), .D(n3438), .Q(
        \inq_ary[12][111] ) );
  LATCHX1_RVT \inq_ary_reg[13][111]  ( .CLK(n3478), .D(n3438), .Q(
        \inq_ary[13][111] ) );
  LATCHX1_RVT \inq_ary_reg[14][111]  ( .CLK(n3477), .D(n3438), .Q(
        \inq_ary[14][111] ) );
  LATCHX1_RVT \inq_ary_reg[15][111]  ( .CLK(n3476), .D(n3438), .Q(
        \inq_ary[15][111] ) );
  LATCHX1_RVT \dout_reg[111]  ( .CLK(n3492), .D(N373), .Q(dout[111]) );
  LATCHX1_RVT \inq_ary_reg[0][110]  ( .CLK(n3491), .D(n3436), .Q(
        \inq_ary[0][110] ) );
  LATCHX1_RVT \inq_ary_reg[1][110]  ( .CLK(n3490), .D(n3436), .Q(
        \inq_ary[1][110] ) );
  LATCHX1_RVT \inq_ary_reg[2][110]  ( .CLK(n3489), .D(n3436), .Q(
        \inq_ary[2][110] ) );
  LATCHX1_RVT \inq_ary_reg[3][110]  ( .CLK(n3488), .D(n3436), .Q(
        \inq_ary[3][110] ) );
  LATCHX1_RVT \inq_ary_reg[4][110]  ( .CLK(n3487), .D(n3436), .Q(
        \inq_ary[4][110] ) );
  LATCHX1_RVT \inq_ary_reg[5][110]  ( .CLK(n3486), .D(n3436), .Q(
        \inq_ary[5][110] ) );
  LATCHX1_RVT \inq_ary_reg[6][110]  ( .CLK(n3485), .D(n3436), .Q(
        \inq_ary[6][110] ) );
  LATCHX1_RVT \inq_ary_reg[7][110]  ( .CLK(n3484), .D(n3436), .Q(
        \inq_ary[7][110] ) );
  LATCHX1_RVT \inq_ary_reg[8][110]  ( .CLK(n3483), .D(n3436), .Q(
        \inq_ary[8][110] ) );
  LATCHX1_RVT \inq_ary_reg[9][110]  ( .CLK(n3482), .D(n3436), .Q(
        \inq_ary[9][110] ) );
  LATCHX1_RVT \inq_ary_reg[10][110]  ( .CLK(n3481), .D(n3436), .Q(
        \inq_ary[10][110] ) );
  LATCHX1_RVT \inq_ary_reg[11][110]  ( .CLK(n3480), .D(n3436), .Q(
        \inq_ary[11][110] ) );
  LATCHX1_RVT \inq_ary_reg[12][110]  ( .CLK(n3479), .D(n3436), .Q(
        \inq_ary[12][110] ) );
  LATCHX1_RVT \inq_ary_reg[13][110]  ( .CLK(n3478), .D(n3436), .Q(
        \inq_ary[13][110] ) );
  LATCHX1_RVT \inq_ary_reg[14][110]  ( .CLK(n3477), .D(n3436), .Q(
        \inq_ary[14][110] ) );
  LATCHX1_RVT \inq_ary_reg[15][110]  ( .CLK(n3476), .D(n3436), .Q(
        \inq_ary[15][110] ) );
  LATCHX1_RVT \dout_reg[110]  ( .CLK(n3492), .D(N372), .Q(dout[110]) );
  LATCHX1_RVT \inq_ary_reg[0][109]  ( .CLK(n3491), .D(n3434), .Q(
        \inq_ary[0][109] ) );
  LATCHX1_RVT \inq_ary_reg[1][109]  ( .CLK(n3490), .D(n3434), .Q(
        \inq_ary[1][109] ) );
  LATCHX1_RVT \inq_ary_reg[2][109]  ( .CLK(n3489), .D(n3434), .Q(
        \inq_ary[2][109] ) );
  LATCHX1_RVT \inq_ary_reg[3][109]  ( .CLK(n3488), .D(n3434), .Q(
        \inq_ary[3][109] ) );
  LATCHX1_RVT \inq_ary_reg[4][109]  ( .CLK(n3487), .D(n3434), .Q(
        \inq_ary[4][109] ) );
  LATCHX1_RVT \inq_ary_reg[5][109]  ( .CLK(n3486), .D(n3434), .Q(
        \inq_ary[5][109] ) );
  LATCHX1_RVT \inq_ary_reg[6][109]  ( .CLK(n3485), .D(n3434), .Q(
        \inq_ary[6][109] ) );
  LATCHX1_RVT \inq_ary_reg[7][109]  ( .CLK(n3484), .D(n3434), .Q(
        \inq_ary[7][109] ) );
  LATCHX1_RVT \inq_ary_reg[8][109]  ( .CLK(n3483), .D(n3434), .Q(
        \inq_ary[8][109] ) );
  LATCHX1_RVT \inq_ary_reg[9][109]  ( .CLK(n3482), .D(n3434), .Q(
        \inq_ary[9][109] ) );
  LATCHX1_RVT \inq_ary_reg[10][109]  ( .CLK(n3481), .D(n3434), .Q(
        \inq_ary[10][109] ) );
  LATCHX1_RVT \inq_ary_reg[11][109]  ( .CLK(n3480), .D(n3434), .Q(
        \inq_ary[11][109] ) );
  LATCHX1_RVT \inq_ary_reg[12][109]  ( .CLK(n3479), .D(n3434), .Q(
        \inq_ary[12][109] ) );
  LATCHX1_RVT \inq_ary_reg[13][109]  ( .CLK(n3478), .D(n3434), .Q(
        \inq_ary[13][109] ) );
  LATCHX1_RVT \inq_ary_reg[14][109]  ( .CLK(n3477), .D(n3434), .Q(
        \inq_ary[14][109] ) );
  LATCHX1_RVT \inq_ary_reg[15][109]  ( .CLK(n3476), .D(n3434), .Q(
        \inq_ary[15][109] ) );
  LATCHX1_RVT \dout_reg[109]  ( .CLK(n3492), .D(N371), .Q(dout[109]) );
  LATCHX1_RVT \inq_ary_reg[0][108]  ( .CLK(n3491), .D(n3432), .Q(
        \inq_ary[0][108] ) );
  LATCHX1_RVT \inq_ary_reg[1][108]  ( .CLK(n3490), .D(n3432), .Q(
        \inq_ary[1][108] ) );
  LATCHX1_RVT \inq_ary_reg[2][108]  ( .CLK(n3489), .D(n3432), .Q(
        \inq_ary[2][108] ) );
  LATCHX1_RVT \inq_ary_reg[3][108]  ( .CLK(n3488), .D(n3432), .Q(
        \inq_ary[3][108] ) );
  LATCHX1_RVT \inq_ary_reg[4][108]  ( .CLK(n3487), .D(n3432), .Q(
        \inq_ary[4][108] ) );
  LATCHX1_RVT \inq_ary_reg[5][108]  ( .CLK(n3486), .D(n3432), .Q(
        \inq_ary[5][108] ) );
  LATCHX1_RVT \inq_ary_reg[6][108]  ( .CLK(n3485), .D(n3432), .Q(
        \inq_ary[6][108] ) );
  LATCHX1_RVT \inq_ary_reg[7][108]  ( .CLK(n3484), .D(n3432), .Q(
        \inq_ary[7][108] ) );
  LATCHX1_RVT \inq_ary_reg[8][108]  ( .CLK(n3483), .D(n3432), .Q(
        \inq_ary[8][108] ) );
  LATCHX1_RVT \inq_ary_reg[9][108]  ( .CLK(n3482), .D(n3432), .Q(
        \inq_ary[9][108] ) );
  LATCHX1_RVT \inq_ary_reg[10][108]  ( .CLK(n3481), .D(n3432), .Q(
        \inq_ary[10][108] ) );
  LATCHX1_RVT \inq_ary_reg[11][108]  ( .CLK(n3480), .D(n3432), .Q(
        \inq_ary[11][108] ) );
  LATCHX1_RVT \inq_ary_reg[12][108]  ( .CLK(n3479), .D(n3432), .Q(
        \inq_ary[12][108] ) );
  LATCHX1_RVT \inq_ary_reg[13][108]  ( .CLK(n3478), .D(n3432), .Q(
        \inq_ary[13][108] ) );
  LATCHX1_RVT \inq_ary_reg[14][108]  ( .CLK(n3477), .D(n3432), .Q(
        \inq_ary[14][108] ) );
  LATCHX1_RVT \inq_ary_reg[15][108]  ( .CLK(n3476), .D(n3432), .Q(
        \inq_ary[15][108] ) );
  LATCHX1_RVT \dout_reg[108]  ( .CLK(n3492), .D(N370), .Q(dout[108]) );
  LATCHX1_RVT \inq_ary_reg[0][107]  ( .CLK(n3491), .D(n3439), .Q(
        \inq_ary[0][107] ) );
  LATCHX1_RVT \inq_ary_reg[1][107]  ( .CLK(n3490), .D(n3439), .Q(
        \inq_ary[1][107] ) );
  LATCHX1_RVT \inq_ary_reg[2][107]  ( .CLK(n3489), .D(n3439), .Q(
        \inq_ary[2][107] ) );
  LATCHX1_RVT \inq_ary_reg[3][107]  ( .CLK(n3488), .D(n3439), .Q(
        \inq_ary[3][107] ) );
  LATCHX1_RVT \inq_ary_reg[4][107]  ( .CLK(n3487), .D(n3439), .Q(
        \inq_ary[4][107] ) );
  LATCHX1_RVT \inq_ary_reg[5][107]  ( .CLK(n3486), .D(n3439), .Q(
        \inq_ary[5][107] ) );
  LATCHX1_RVT \inq_ary_reg[6][107]  ( .CLK(n3485), .D(n3439), .Q(
        \inq_ary[6][107] ) );
  LATCHX1_RVT \inq_ary_reg[7][107]  ( .CLK(n3484), .D(n3439), .Q(
        \inq_ary[7][107] ) );
  LATCHX1_RVT \inq_ary_reg[8][107]  ( .CLK(n3483), .D(n3439), .Q(
        \inq_ary[8][107] ) );
  LATCHX1_RVT \inq_ary_reg[9][107]  ( .CLK(n3482), .D(n3439), .Q(
        \inq_ary[9][107] ) );
  LATCHX1_RVT \inq_ary_reg[10][107]  ( .CLK(n3481), .D(n3439), .Q(
        \inq_ary[10][107] ) );
  LATCHX1_RVT \inq_ary_reg[11][107]  ( .CLK(n3480), .D(n3439), .Q(
        \inq_ary[11][107] ) );
  LATCHX1_RVT \inq_ary_reg[12][107]  ( .CLK(n3479), .D(n3439), .Q(
        \inq_ary[12][107] ) );
  LATCHX1_RVT \inq_ary_reg[13][107]  ( .CLK(n3478), .D(n3439), .Q(
        \inq_ary[13][107] ) );
  LATCHX1_RVT \inq_ary_reg[14][107]  ( .CLK(n3477), .D(n3439), .Q(
        \inq_ary[14][107] ) );
  LATCHX1_RVT \inq_ary_reg[15][107]  ( .CLK(n3476), .D(n3439), .Q(
        \inq_ary[15][107] ) );
  LATCHX1_RVT \dout_reg[107]  ( .CLK(n3492), .D(N369), .Q(dout[107]) );
  LATCHX1_RVT \inq_ary_reg[0][106]  ( .CLK(n3491), .D(n3437), .Q(
        \inq_ary[0][106] ) );
  LATCHX1_RVT \inq_ary_reg[1][106]  ( .CLK(n3490), .D(n3437), .Q(
        \inq_ary[1][106] ) );
  LATCHX1_RVT \inq_ary_reg[2][106]  ( .CLK(n3489), .D(n3437), .Q(
        \inq_ary[2][106] ) );
  LATCHX1_RVT \inq_ary_reg[3][106]  ( .CLK(n3488), .D(n3437), .Q(
        \inq_ary[3][106] ) );
  LATCHX1_RVT \inq_ary_reg[4][106]  ( .CLK(n3487), .D(n3437), .Q(
        \inq_ary[4][106] ) );
  LATCHX1_RVT \inq_ary_reg[5][106]  ( .CLK(n3486), .D(n3437), .Q(
        \inq_ary[5][106] ) );
  LATCHX1_RVT \inq_ary_reg[6][106]  ( .CLK(n3485), .D(n3437), .Q(
        \inq_ary[6][106] ) );
  LATCHX1_RVT \inq_ary_reg[7][106]  ( .CLK(n3484), .D(n3437), .Q(
        \inq_ary[7][106] ) );
  LATCHX1_RVT \inq_ary_reg[8][106]  ( .CLK(n3483), .D(n3437), .Q(
        \inq_ary[8][106] ) );
  LATCHX1_RVT \inq_ary_reg[9][106]  ( .CLK(n3482), .D(n3437), .Q(
        \inq_ary[9][106] ) );
  LATCHX1_RVT \inq_ary_reg[10][106]  ( .CLK(n3481), .D(n3437), .Q(
        \inq_ary[10][106] ) );
  LATCHX1_RVT \inq_ary_reg[11][106]  ( .CLK(n3480), .D(n3437), .Q(
        \inq_ary[11][106] ) );
  LATCHX1_RVT \inq_ary_reg[12][106]  ( .CLK(n3479), .D(n3437), .Q(
        \inq_ary[12][106] ) );
  LATCHX1_RVT \inq_ary_reg[13][106]  ( .CLK(n3478), .D(n3437), .Q(
        \inq_ary[13][106] ) );
  LATCHX1_RVT \inq_ary_reg[14][106]  ( .CLK(n3477), .D(n3437), .Q(
        \inq_ary[14][106] ) );
  LATCHX1_RVT \inq_ary_reg[15][106]  ( .CLK(n3476), .D(n3437), .Q(
        \inq_ary[15][106] ) );
  LATCHX1_RVT \dout_reg[106]  ( .CLK(n3492), .D(N368), .Q(dout[106]) );
  LATCHX1_RVT \inq_ary_reg[0][105]  ( .CLK(n3491), .D(n3435), .Q(
        \inq_ary[0][105] ) );
  LATCHX1_RVT \inq_ary_reg[1][105]  ( .CLK(n3490), .D(n3435), .Q(
        \inq_ary[1][105] ) );
  LATCHX1_RVT \inq_ary_reg[2][105]  ( .CLK(n3489), .D(n3435), .Q(
        \inq_ary[2][105] ) );
  LATCHX1_RVT \inq_ary_reg[3][105]  ( .CLK(n3488), .D(n3435), .Q(
        \inq_ary[3][105] ) );
  LATCHX1_RVT \inq_ary_reg[4][105]  ( .CLK(n3487), .D(n3435), .Q(
        \inq_ary[4][105] ) );
  LATCHX1_RVT \inq_ary_reg[5][105]  ( .CLK(n3486), .D(n3435), .Q(
        \inq_ary[5][105] ) );
  LATCHX1_RVT \inq_ary_reg[6][105]  ( .CLK(n3485), .D(n3435), .Q(
        \inq_ary[6][105] ) );
  LATCHX1_RVT \inq_ary_reg[7][105]  ( .CLK(n3484), .D(n3435), .Q(
        \inq_ary[7][105] ) );
  LATCHX1_RVT \inq_ary_reg[8][105]  ( .CLK(n3483), .D(n3435), .Q(
        \inq_ary[8][105] ) );
  LATCHX1_RVT \inq_ary_reg[9][105]  ( .CLK(n3482), .D(n3435), .Q(
        \inq_ary[9][105] ) );
  LATCHX1_RVT \inq_ary_reg[10][105]  ( .CLK(n3481), .D(n3435), .Q(
        \inq_ary[10][105] ) );
  LATCHX1_RVT \inq_ary_reg[11][105]  ( .CLK(n3480), .D(n3435), .Q(
        \inq_ary[11][105] ) );
  LATCHX1_RVT \inq_ary_reg[12][105]  ( .CLK(n3479), .D(n3435), .Q(
        \inq_ary[12][105] ) );
  LATCHX1_RVT \inq_ary_reg[13][105]  ( .CLK(n3478), .D(n3435), .Q(
        \inq_ary[13][105] ) );
  LATCHX1_RVT \inq_ary_reg[14][105]  ( .CLK(n3477), .D(n3435), .Q(
        \inq_ary[14][105] ) );
  LATCHX1_RVT \inq_ary_reg[15][105]  ( .CLK(n3476), .D(n3435), .Q(
        \inq_ary[15][105] ) );
  LATCHX1_RVT \dout_reg[105]  ( .CLK(n3492), .D(N367), .Q(dout[105]) );
  LATCHX1_RVT \inq_ary_reg[0][104]  ( .CLK(n3491), .D(n3433), .Q(
        \inq_ary[0][104] ) );
  LATCHX1_RVT \inq_ary_reg[1][104]  ( .CLK(n3490), .D(n3433), .Q(
        \inq_ary[1][104] ) );
  LATCHX1_RVT \inq_ary_reg[2][104]  ( .CLK(n3489), .D(n3433), .Q(
        \inq_ary[2][104] ) );
  LATCHX1_RVT \inq_ary_reg[3][104]  ( .CLK(n3488), .D(n3433), .Q(
        \inq_ary[3][104] ) );
  LATCHX1_RVT \inq_ary_reg[4][104]  ( .CLK(n3487), .D(n3433), .Q(
        \inq_ary[4][104] ) );
  LATCHX1_RVT \inq_ary_reg[5][104]  ( .CLK(n3486), .D(n3433), .Q(
        \inq_ary[5][104] ) );
  LATCHX1_RVT \inq_ary_reg[6][104]  ( .CLK(n3485), .D(n3433), .Q(
        \inq_ary[6][104] ) );
  LATCHX1_RVT \inq_ary_reg[7][104]  ( .CLK(n3484), .D(n3433), .Q(
        \inq_ary[7][104] ) );
  LATCHX1_RVT \inq_ary_reg[8][104]  ( .CLK(n3483), .D(n3433), .Q(
        \inq_ary[8][104] ) );
  LATCHX1_RVT \inq_ary_reg[9][104]  ( .CLK(n3482), .D(n3433), .Q(
        \inq_ary[9][104] ) );
  LATCHX1_RVT \inq_ary_reg[10][104]  ( .CLK(n3481), .D(n3433), .Q(
        \inq_ary[10][104] ) );
  LATCHX1_RVT \inq_ary_reg[11][104]  ( .CLK(n3480), .D(n3433), .Q(
        \inq_ary[11][104] ) );
  LATCHX1_RVT \inq_ary_reg[12][104]  ( .CLK(n3479), .D(n3433), .Q(
        \inq_ary[12][104] ) );
  LATCHX1_RVT \inq_ary_reg[13][104]  ( .CLK(n3478), .D(n3433), .Q(
        \inq_ary[13][104] ) );
  LATCHX1_RVT \inq_ary_reg[14][104]  ( .CLK(n3477), .D(n3433), .Q(
        \inq_ary[14][104] ) );
  LATCHX1_RVT \inq_ary_reg[15][104]  ( .CLK(n3476), .D(n3433), .Q(
        \inq_ary[15][104] ) );
  LATCHX1_RVT \dout_reg[104]  ( .CLK(n3492), .D(N366), .Q(dout[104]) );
  LATCHX1_RVT \inq_ary_reg[0][103]  ( .CLK(n3491), .D(n3430), .Q(
        \inq_ary[0][103] ) );
  LATCHX1_RVT \inq_ary_reg[1][103]  ( .CLK(n3490), .D(n3430), .Q(
        \inq_ary[1][103] ) );
  LATCHX1_RVT \inq_ary_reg[2][103]  ( .CLK(n3489), .D(n3430), .Q(
        \inq_ary[2][103] ) );
  LATCHX1_RVT \inq_ary_reg[3][103]  ( .CLK(n3488), .D(n3430), .Q(
        \inq_ary[3][103] ) );
  LATCHX1_RVT \inq_ary_reg[4][103]  ( .CLK(n3487), .D(n3430), .Q(
        \inq_ary[4][103] ) );
  LATCHX1_RVT \inq_ary_reg[5][103]  ( .CLK(n3486), .D(n3430), .Q(
        \inq_ary[5][103] ) );
  LATCHX1_RVT \inq_ary_reg[6][103]  ( .CLK(n3485), .D(n3430), .Q(
        \inq_ary[6][103] ) );
  LATCHX1_RVT \inq_ary_reg[7][103]  ( .CLK(n3484), .D(n3430), .Q(
        \inq_ary[7][103] ) );
  LATCHX1_RVT \inq_ary_reg[8][103]  ( .CLK(n3483), .D(n3430), .Q(
        \inq_ary[8][103] ) );
  LATCHX1_RVT \inq_ary_reg[9][103]  ( .CLK(n3482), .D(n3430), .Q(
        \inq_ary[9][103] ) );
  LATCHX1_RVT \inq_ary_reg[10][103]  ( .CLK(n3481), .D(n3430), .Q(
        \inq_ary[10][103] ) );
  LATCHX1_RVT \inq_ary_reg[11][103]  ( .CLK(n3480), .D(n3430), .Q(
        \inq_ary[11][103] ) );
  LATCHX1_RVT \inq_ary_reg[12][103]  ( .CLK(n3479), .D(n3430), .Q(
        \inq_ary[12][103] ) );
  LATCHX1_RVT \inq_ary_reg[13][103]  ( .CLK(n3478), .D(n3430), .Q(
        \inq_ary[13][103] ) );
  LATCHX1_RVT \inq_ary_reg[14][103]  ( .CLK(n3477), .D(n3430), .Q(
        \inq_ary[14][103] ) );
  LATCHX1_RVT \inq_ary_reg[15][103]  ( .CLK(n3476), .D(n3430), .Q(
        \inq_ary[15][103] ) );
  LATCHX1_RVT \dout_reg[103]  ( .CLK(n3492), .D(N365), .Q(dout[103]) );
  LATCHX1_RVT \inq_ary_reg[0][102]  ( .CLK(n3491), .D(n3428), .Q(
        \inq_ary[0][102] ) );
  LATCHX1_RVT \inq_ary_reg[1][102]  ( .CLK(n3490), .D(n3428), .Q(
        \inq_ary[1][102] ) );
  LATCHX1_RVT \inq_ary_reg[2][102]  ( .CLK(n3489), .D(n3428), .Q(
        \inq_ary[2][102] ) );
  LATCHX1_RVT \inq_ary_reg[3][102]  ( .CLK(n3488), .D(n3428), .Q(
        \inq_ary[3][102] ) );
  LATCHX1_RVT \inq_ary_reg[4][102]  ( .CLK(n3487), .D(n3428), .Q(
        \inq_ary[4][102] ) );
  LATCHX1_RVT \inq_ary_reg[5][102]  ( .CLK(n3486), .D(n3428), .Q(
        \inq_ary[5][102] ) );
  LATCHX1_RVT \inq_ary_reg[6][102]  ( .CLK(n3485), .D(n3428), .Q(
        \inq_ary[6][102] ) );
  LATCHX1_RVT \inq_ary_reg[7][102]  ( .CLK(n3484), .D(n3428), .Q(
        \inq_ary[7][102] ) );
  LATCHX1_RVT \inq_ary_reg[8][102]  ( .CLK(n3483), .D(n3428), .Q(
        \inq_ary[8][102] ) );
  LATCHX1_RVT \inq_ary_reg[9][102]  ( .CLK(n3482), .D(n3428), .Q(
        \inq_ary[9][102] ) );
  LATCHX1_RVT \inq_ary_reg[10][102]  ( .CLK(n3481), .D(n3428), .Q(
        \inq_ary[10][102] ) );
  LATCHX1_RVT \inq_ary_reg[11][102]  ( .CLK(n3480), .D(n3428), .Q(
        \inq_ary[11][102] ) );
  LATCHX1_RVT \inq_ary_reg[12][102]  ( .CLK(n3479), .D(n3428), .Q(
        \inq_ary[12][102] ) );
  LATCHX1_RVT \inq_ary_reg[13][102]  ( .CLK(n3478), .D(n3428), .Q(
        \inq_ary[13][102] ) );
  LATCHX1_RVT \inq_ary_reg[14][102]  ( .CLK(n3477), .D(n3428), .Q(
        \inq_ary[14][102] ) );
  LATCHX1_RVT \inq_ary_reg[15][102]  ( .CLK(n3476), .D(n3428), .Q(
        \inq_ary[15][102] ) );
  LATCHX1_RVT \dout_reg[102]  ( .CLK(n3492), .D(N364), .Q(dout[102]) );
  LATCHX1_RVT \inq_ary_reg[0][101]  ( .CLK(n3491), .D(n3426), .Q(
        \inq_ary[0][101] ) );
  LATCHX1_RVT \inq_ary_reg[1][101]  ( .CLK(n3490), .D(n3426), .Q(
        \inq_ary[1][101] ) );
  LATCHX1_RVT \inq_ary_reg[2][101]  ( .CLK(n3489), .D(n3426), .Q(
        \inq_ary[2][101] ) );
  LATCHX1_RVT \inq_ary_reg[3][101]  ( .CLK(n3488), .D(n3426), .Q(
        \inq_ary[3][101] ) );
  LATCHX1_RVT \inq_ary_reg[4][101]  ( .CLK(n3487), .D(n3426), .Q(
        \inq_ary[4][101] ) );
  LATCHX1_RVT \inq_ary_reg[5][101]  ( .CLK(n3486), .D(n3426), .Q(
        \inq_ary[5][101] ) );
  LATCHX1_RVT \inq_ary_reg[6][101]  ( .CLK(n3485), .D(n3426), .Q(
        \inq_ary[6][101] ) );
  LATCHX1_RVT \inq_ary_reg[7][101]  ( .CLK(n3484), .D(n3426), .Q(
        \inq_ary[7][101] ) );
  LATCHX1_RVT \inq_ary_reg[8][101]  ( .CLK(n3483), .D(n3426), .Q(
        \inq_ary[8][101] ) );
  LATCHX1_RVT \inq_ary_reg[9][101]  ( .CLK(n3482), .D(n3426), .Q(
        \inq_ary[9][101] ) );
  LATCHX1_RVT \inq_ary_reg[10][101]  ( .CLK(n3481), .D(n3426), .Q(
        \inq_ary[10][101] ) );
  LATCHX1_RVT \inq_ary_reg[11][101]  ( .CLK(n3480), .D(n3426), .Q(
        \inq_ary[11][101] ) );
  LATCHX1_RVT \inq_ary_reg[12][101]  ( .CLK(n3479), .D(n3426), .Q(
        \inq_ary[12][101] ) );
  LATCHX1_RVT \inq_ary_reg[13][101]  ( .CLK(n3478), .D(n3426), .Q(
        \inq_ary[13][101] ) );
  LATCHX1_RVT \inq_ary_reg[14][101]  ( .CLK(n3477), .D(n3426), .Q(
        \inq_ary[14][101] ) );
  LATCHX1_RVT \inq_ary_reg[15][101]  ( .CLK(n3476), .D(n3426), .Q(
        \inq_ary[15][101] ) );
  LATCHX1_RVT \dout_reg[101]  ( .CLK(n3492), .D(N363), .Q(dout[101]) );
  LATCHX1_RVT \inq_ary_reg[0][100]  ( .CLK(n3491), .D(n3424), .Q(
        \inq_ary[0][100] ) );
  LATCHX1_RVT \inq_ary_reg[1][100]  ( .CLK(n3490), .D(n3424), .Q(
        \inq_ary[1][100] ) );
  LATCHX1_RVT \inq_ary_reg[2][100]  ( .CLK(n3489), .D(n3424), .Q(
        \inq_ary[2][100] ) );
  LATCHX1_RVT \inq_ary_reg[3][100]  ( .CLK(n3488), .D(n3424), .Q(
        \inq_ary[3][100] ) );
  LATCHX1_RVT \inq_ary_reg[4][100]  ( .CLK(n3487), .D(n3424), .Q(
        \inq_ary[4][100] ) );
  LATCHX1_RVT \inq_ary_reg[5][100]  ( .CLK(n3486), .D(n3424), .Q(
        \inq_ary[5][100] ) );
  LATCHX1_RVT \inq_ary_reg[6][100]  ( .CLK(n3485), .D(n3424), .Q(
        \inq_ary[6][100] ) );
  LATCHX1_RVT \inq_ary_reg[7][100]  ( .CLK(n3484), .D(n3424), .Q(
        \inq_ary[7][100] ) );
  LATCHX1_RVT \inq_ary_reg[8][100]  ( .CLK(n3483), .D(n3424), .Q(
        \inq_ary[8][100] ) );
  LATCHX1_RVT \inq_ary_reg[9][100]  ( .CLK(n3482), .D(n3424), .Q(
        \inq_ary[9][100] ) );
  LATCHX1_RVT \inq_ary_reg[10][100]  ( .CLK(n3481), .D(n3424), .Q(
        \inq_ary[10][100] ) );
  LATCHX1_RVT \inq_ary_reg[11][100]  ( .CLK(n3480), .D(n3424), .Q(
        \inq_ary[11][100] ) );
  LATCHX1_RVT \inq_ary_reg[12][100]  ( .CLK(n3479), .D(n3424), .Q(
        \inq_ary[12][100] ) );
  LATCHX1_RVT \inq_ary_reg[13][100]  ( .CLK(n3478), .D(n3424), .Q(
        \inq_ary[13][100] ) );
  LATCHX1_RVT \inq_ary_reg[14][100]  ( .CLK(n3477), .D(n3424), .Q(
        \inq_ary[14][100] ) );
  LATCHX1_RVT \inq_ary_reg[15][100]  ( .CLK(n3476), .D(n3424), .Q(
        \inq_ary[15][100] ) );
  LATCHX1_RVT \dout_reg[100]  ( .CLK(n3492), .D(N362), .Q(dout[100]) );
  LATCHX1_RVT \inq_ary_reg[0][99]  ( .CLK(n3491), .D(n3431), .Q(
        \inq_ary[0][99] ) );
  LATCHX1_RVT \inq_ary_reg[1][99]  ( .CLK(n3490), .D(n3431), .Q(
        \inq_ary[1][99] ) );
  LATCHX1_RVT \inq_ary_reg[2][99]  ( .CLK(n3489), .D(n3431), .Q(
        \inq_ary[2][99] ) );
  LATCHX1_RVT \inq_ary_reg[3][99]  ( .CLK(n3488), .D(n3431), .Q(
        \inq_ary[3][99] ) );
  LATCHX1_RVT \inq_ary_reg[4][99]  ( .CLK(n3487), .D(n3431), .Q(
        \inq_ary[4][99] ) );
  LATCHX1_RVT \inq_ary_reg[5][99]  ( .CLK(n3486), .D(n3431), .Q(
        \inq_ary[5][99] ) );
  LATCHX1_RVT \inq_ary_reg[6][99]  ( .CLK(n3485), .D(n3431), .Q(
        \inq_ary[6][99] ) );
  LATCHX1_RVT \inq_ary_reg[7][99]  ( .CLK(n3484), .D(n3431), .Q(
        \inq_ary[7][99] ) );
  LATCHX1_RVT \inq_ary_reg[8][99]  ( .CLK(n3483), .D(n3431), .Q(
        \inq_ary[8][99] ) );
  LATCHX1_RVT \inq_ary_reg[9][99]  ( .CLK(n3482), .D(n3431), .Q(
        \inq_ary[9][99] ) );
  LATCHX1_RVT \inq_ary_reg[10][99]  ( .CLK(n3481), .D(n3431), .Q(
        \inq_ary[10][99] ) );
  LATCHX1_RVT \inq_ary_reg[11][99]  ( .CLK(n3480), .D(n3431), .Q(
        \inq_ary[11][99] ) );
  LATCHX1_RVT \inq_ary_reg[12][99]  ( .CLK(n3479), .D(n3431), .Q(
        \inq_ary[12][99] ) );
  LATCHX1_RVT \inq_ary_reg[13][99]  ( .CLK(n3478), .D(n3431), .Q(
        \inq_ary[13][99] ) );
  LATCHX1_RVT \inq_ary_reg[14][99]  ( .CLK(n3477), .D(n3431), .Q(
        \inq_ary[14][99] ) );
  LATCHX1_RVT \inq_ary_reg[15][99]  ( .CLK(n3476), .D(n3431), .Q(
        \inq_ary[15][99] ) );
  LATCHX1_RVT \dout_reg[99]  ( .CLK(n3492), .D(N361), .Q(dout[99]) );
  LATCHX1_RVT \inq_ary_reg[0][98]  ( .CLK(n3491), .D(n3429), .Q(
        \inq_ary[0][98] ) );
  LATCHX1_RVT \inq_ary_reg[1][98]  ( .CLK(n3490), .D(n3429), .Q(
        \inq_ary[1][98] ) );
  LATCHX1_RVT \inq_ary_reg[2][98]  ( .CLK(n3489), .D(n3429), .Q(
        \inq_ary[2][98] ) );
  LATCHX1_RVT \inq_ary_reg[3][98]  ( .CLK(n3488), .D(n3429), .Q(
        \inq_ary[3][98] ) );
  LATCHX1_RVT \inq_ary_reg[4][98]  ( .CLK(n3487), .D(n3429), .Q(
        \inq_ary[4][98] ) );
  LATCHX1_RVT \inq_ary_reg[5][98]  ( .CLK(n3486), .D(n3429), .Q(
        \inq_ary[5][98] ) );
  LATCHX1_RVT \inq_ary_reg[6][98]  ( .CLK(n3485), .D(n3429), .Q(
        \inq_ary[6][98] ) );
  LATCHX1_RVT \inq_ary_reg[7][98]  ( .CLK(n3484), .D(n3429), .Q(
        \inq_ary[7][98] ) );
  LATCHX1_RVT \inq_ary_reg[8][98]  ( .CLK(n3483), .D(n3429), .Q(
        \inq_ary[8][98] ) );
  LATCHX1_RVT \inq_ary_reg[9][98]  ( .CLK(n3482), .D(n3429), .Q(
        \inq_ary[9][98] ) );
  LATCHX1_RVT \inq_ary_reg[10][98]  ( .CLK(n3481), .D(n3429), .Q(
        \inq_ary[10][98] ) );
  LATCHX1_RVT \inq_ary_reg[11][98]  ( .CLK(n3480), .D(n3429), .Q(
        \inq_ary[11][98] ) );
  LATCHX1_RVT \inq_ary_reg[12][98]  ( .CLK(n3479), .D(n3429), .Q(
        \inq_ary[12][98] ) );
  LATCHX1_RVT \inq_ary_reg[13][98]  ( .CLK(n3478), .D(n3429), .Q(
        \inq_ary[13][98] ) );
  LATCHX1_RVT \inq_ary_reg[14][98]  ( .CLK(n3477), .D(n3429), .Q(
        \inq_ary[14][98] ) );
  LATCHX1_RVT \inq_ary_reg[15][98]  ( .CLK(n3476), .D(n3429), .Q(
        \inq_ary[15][98] ) );
  LATCHX1_RVT \dout_reg[98]  ( .CLK(n3492), .D(N359), .Q(dout[98]) );
  LATCHX1_RVT \inq_ary_reg[0][97]  ( .CLK(n3491), .D(n3427), .Q(
        \inq_ary[0][97] ) );
  LATCHX1_RVT \inq_ary_reg[1][97]  ( .CLK(n3490), .D(n3427), .Q(
        \inq_ary[1][97] ) );
  LATCHX1_RVT \inq_ary_reg[2][97]  ( .CLK(n3489), .D(n3427), .Q(
        \inq_ary[2][97] ) );
  LATCHX1_RVT \inq_ary_reg[3][97]  ( .CLK(n3488), .D(n3427), .Q(
        \inq_ary[3][97] ) );
  LATCHX1_RVT \inq_ary_reg[4][97]  ( .CLK(n3487), .D(n3427), .Q(
        \inq_ary[4][97] ) );
  LATCHX1_RVT \inq_ary_reg[5][97]  ( .CLK(n3486), .D(n3427), .Q(
        \inq_ary[5][97] ) );
  LATCHX1_RVT \inq_ary_reg[6][97]  ( .CLK(n3485), .D(n3427), .Q(
        \inq_ary[6][97] ) );
  LATCHX1_RVT \inq_ary_reg[7][97]  ( .CLK(n3484), .D(n3427), .Q(
        \inq_ary[7][97] ) );
  LATCHX1_RVT \inq_ary_reg[8][97]  ( .CLK(n3483), .D(n3427), .Q(
        \inq_ary[8][97] ) );
  LATCHX1_RVT \inq_ary_reg[9][97]  ( .CLK(n3482), .D(n3427), .Q(
        \inq_ary[9][97] ) );
  LATCHX1_RVT \inq_ary_reg[10][97]  ( .CLK(n3481), .D(n3427), .Q(
        \inq_ary[10][97] ) );
  LATCHX1_RVT \inq_ary_reg[11][97]  ( .CLK(n3480), .D(n3427), .Q(
        \inq_ary[11][97] ) );
  LATCHX1_RVT \inq_ary_reg[12][97]  ( .CLK(n3479), .D(n3427), .Q(
        \inq_ary[12][97] ) );
  LATCHX1_RVT \inq_ary_reg[13][97]  ( .CLK(n3478), .D(n3427), .Q(
        \inq_ary[13][97] ) );
  LATCHX1_RVT \inq_ary_reg[14][97]  ( .CLK(n3477), .D(n3427), .Q(
        \inq_ary[14][97] ) );
  LATCHX1_RVT \inq_ary_reg[15][97]  ( .CLK(n3476), .D(n3427), .Q(
        \inq_ary[15][97] ) );
  LATCHX1_RVT \dout_reg[97]  ( .CLK(n3492), .D(N358), .Q(dout[97]) );
  LATCHX1_RVT \inq_ary_reg[0][96]  ( .CLK(n3491), .D(n3425), .Q(
        \inq_ary[0][96] ) );
  LATCHX1_RVT \inq_ary_reg[1][96]  ( .CLK(n3490), .D(n3425), .Q(
        \inq_ary[1][96] ) );
  LATCHX1_RVT \inq_ary_reg[2][96]  ( .CLK(n3489), .D(n3425), .Q(
        \inq_ary[2][96] ) );
  LATCHX1_RVT \inq_ary_reg[3][96]  ( .CLK(n3488), .D(n3425), .Q(
        \inq_ary[3][96] ) );
  LATCHX1_RVT \inq_ary_reg[4][96]  ( .CLK(n3487), .D(n3425), .Q(
        \inq_ary[4][96] ) );
  LATCHX1_RVT \inq_ary_reg[5][96]  ( .CLK(n3486), .D(n3425), .Q(
        \inq_ary[5][96] ) );
  LATCHX1_RVT \inq_ary_reg[6][96]  ( .CLK(n3485), .D(n3425), .Q(
        \inq_ary[6][96] ) );
  LATCHX1_RVT \inq_ary_reg[7][96]  ( .CLK(n3484), .D(n3425), .Q(
        \inq_ary[7][96] ) );
  LATCHX1_RVT \inq_ary_reg[8][96]  ( .CLK(n3483), .D(n3425), .Q(
        \inq_ary[8][96] ) );
  LATCHX1_RVT \inq_ary_reg[9][96]  ( .CLK(n3482), .D(n3425), .Q(
        \inq_ary[9][96] ) );
  LATCHX1_RVT \inq_ary_reg[10][96]  ( .CLK(n3481), .D(n3425), .Q(
        \inq_ary[10][96] ) );
  LATCHX1_RVT \inq_ary_reg[11][96]  ( .CLK(n3480), .D(n3425), .Q(
        \inq_ary[11][96] ) );
  LATCHX1_RVT \inq_ary_reg[12][96]  ( .CLK(n3479), .D(n3425), .Q(
        \inq_ary[12][96] ) );
  LATCHX1_RVT \inq_ary_reg[13][96]  ( .CLK(n3478), .D(n3425), .Q(
        \inq_ary[13][96] ) );
  LATCHX1_RVT \inq_ary_reg[14][96]  ( .CLK(n3477), .D(n3425), .Q(
        \inq_ary[14][96] ) );
  LATCHX1_RVT \inq_ary_reg[15][96]  ( .CLK(n3476), .D(n3425), .Q(
        \inq_ary[15][96] ) );
  LATCHX1_RVT \dout_reg[96]  ( .CLK(n3492), .D(N357), .Q(dout[96]) );
  LATCHX1_RVT \inq_ary_reg[0][95]  ( .CLK(n3491), .D(n3422), .Q(
        \inq_ary[0][95] ) );
  LATCHX1_RVT \inq_ary_reg[1][95]  ( .CLK(n3490), .D(n3422), .Q(
        \inq_ary[1][95] ) );
  LATCHX1_RVT \inq_ary_reg[2][95]  ( .CLK(n3489), .D(n3422), .Q(
        \inq_ary[2][95] ) );
  LATCHX1_RVT \inq_ary_reg[3][95]  ( .CLK(n3488), .D(n3422), .Q(
        \inq_ary[3][95] ) );
  LATCHX1_RVT \inq_ary_reg[4][95]  ( .CLK(n3487), .D(n3422), .Q(
        \inq_ary[4][95] ) );
  LATCHX1_RVT \inq_ary_reg[5][95]  ( .CLK(n3486), .D(n3422), .Q(
        \inq_ary[5][95] ) );
  LATCHX1_RVT \inq_ary_reg[6][95]  ( .CLK(n3485), .D(n3422), .Q(
        \inq_ary[6][95] ) );
  LATCHX1_RVT \inq_ary_reg[7][95]  ( .CLK(n3484), .D(n3422), .Q(
        \inq_ary[7][95] ) );
  LATCHX1_RVT \inq_ary_reg[8][95]  ( .CLK(n3483), .D(n3422), .Q(
        \inq_ary[8][95] ) );
  LATCHX1_RVT \inq_ary_reg[9][95]  ( .CLK(n3482), .D(n3422), .Q(
        \inq_ary[9][95] ) );
  LATCHX1_RVT \inq_ary_reg[10][95]  ( .CLK(n3481), .D(n3422), .Q(
        \inq_ary[10][95] ) );
  LATCHX1_RVT \inq_ary_reg[11][95]  ( .CLK(n3480), .D(n3422), .Q(
        \inq_ary[11][95] ) );
  LATCHX1_RVT \inq_ary_reg[12][95]  ( .CLK(n3479), .D(n3422), .Q(
        \inq_ary[12][95] ) );
  LATCHX1_RVT \inq_ary_reg[13][95]  ( .CLK(n3478), .D(n3422), .Q(
        \inq_ary[13][95] ) );
  LATCHX1_RVT \inq_ary_reg[14][95]  ( .CLK(n3477), .D(n3422), .Q(
        \inq_ary[14][95] ) );
  LATCHX1_RVT \inq_ary_reg[15][95]  ( .CLK(n3476), .D(n3422), .Q(
        \inq_ary[15][95] ) );
  LATCHX1_RVT \dout_reg[95]  ( .CLK(n3492), .D(N356), .Q(dout[95]) );
  LATCHX1_RVT \inq_ary_reg[0][94]  ( .CLK(n3491), .D(n3420), .Q(
        \inq_ary[0][94] ) );
  LATCHX1_RVT \inq_ary_reg[1][94]  ( .CLK(n3490), .D(n3420), .Q(
        \inq_ary[1][94] ) );
  LATCHX1_RVT \inq_ary_reg[2][94]  ( .CLK(n3489), .D(n3420), .Q(
        \inq_ary[2][94] ) );
  LATCHX1_RVT \inq_ary_reg[3][94]  ( .CLK(n3488), .D(n3420), .Q(
        \inq_ary[3][94] ) );
  LATCHX1_RVT \inq_ary_reg[4][94]  ( .CLK(n3487), .D(n3420), .Q(
        \inq_ary[4][94] ) );
  LATCHX1_RVT \inq_ary_reg[5][94]  ( .CLK(n3486), .D(n3420), .Q(
        \inq_ary[5][94] ) );
  LATCHX1_RVT \inq_ary_reg[6][94]  ( .CLK(n3485), .D(n3420), .Q(
        \inq_ary[6][94] ) );
  LATCHX1_RVT \inq_ary_reg[7][94]  ( .CLK(n3484), .D(n3420), .Q(
        \inq_ary[7][94] ) );
  LATCHX1_RVT \inq_ary_reg[8][94]  ( .CLK(n3483), .D(n3420), .Q(
        \inq_ary[8][94] ) );
  LATCHX1_RVT \inq_ary_reg[9][94]  ( .CLK(n3482), .D(n3420), .Q(
        \inq_ary[9][94] ) );
  LATCHX1_RVT \inq_ary_reg[10][94]  ( .CLK(n3481), .D(n3420), .Q(
        \inq_ary[10][94] ) );
  LATCHX1_RVT \inq_ary_reg[11][94]  ( .CLK(n3480), .D(n3420), .Q(
        \inq_ary[11][94] ) );
  LATCHX1_RVT \inq_ary_reg[12][94]  ( .CLK(n3479), .D(n3420), .Q(
        \inq_ary[12][94] ) );
  LATCHX1_RVT \inq_ary_reg[13][94]  ( .CLK(n3478), .D(n3420), .Q(
        \inq_ary[13][94] ) );
  LATCHX1_RVT \inq_ary_reg[14][94]  ( .CLK(n3477), .D(n3420), .Q(
        \inq_ary[14][94] ) );
  LATCHX1_RVT \inq_ary_reg[15][94]  ( .CLK(n3476), .D(n3420), .Q(
        \inq_ary[15][94] ) );
  LATCHX1_RVT \dout_reg[94]  ( .CLK(n3492), .D(N355), .Q(dout[94]) );
  LATCHX1_RVT \inq_ary_reg[0][93]  ( .CLK(n3491), .D(n3418), .Q(
        \inq_ary[0][93] ) );
  LATCHX1_RVT \inq_ary_reg[1][93]  ( .CLK(n3490), .D(n3418), .Q(
        \inq_ary[1][93] ) );
  LATCHX1_RVT \inq_ary_reg[2][93]  ( .CLK(n3489), .D(n3418), .Q(
        \inq_ary[2][93] ) );
  LATCHX1_RVT \inq_ary_reg[3][93]  ( .CLK(n3488), .D(n3418), .Q(
        \inq_ary[3][93] ) );
  LATCHX1_RVT \inq_ary_reg[4][93]  ( .CLK(n3487), .D(n3418), .Q(
        \inq_ary[4][93] ) );
  LATCHX1_RVT \inq_ary_reg[5][93]  ( .CLK(n3486), .D(n3418), .Q(
        \inq_ary[5][93] ) );
  LATCHX1_RVT \inq_ary_reg[6][93]  ( .CLK(n3485), .D(n3418), .Q(
        \inq_ary[6][93] ) );
  LATCHX1_RVT \inq_ary_reg[7][93]  ( .CLK(n3484), .D(n3418), .Q(
        \inq_ary[7][93] ) );
  LATCHX1_RVT \inq_ary_reg[8][93]  ( .CLK(n3483), .D(n3418), .Q(
        \inq_ary[8][93] ) );
  LATCHX1_RVT \inq_ary_reg[9][93]  ( .CLK(n3482), .D(n3418), .Q(
        \inq_ary[9][93] ) );
  LATCHX1_RVT \inq_ary_reg[10][93]  ( .CLK(n3481), .D(n3418), .Q(
        \inq_ary[10][93] ) );
  LATCHX1_RVT \inq_ary_reg[11][93]  ( .CLK(n3480), .D(n3418), .Q(
        \inq_ary[11][93] ) );
  LATCHX1_RVT \inq_ary_reg[12][93]  ( .CLK(n3479), .D(n3418), .Q(
        \inq_ary[12][93] ) );
  LATCHX1_RVT \inq_ary_reg[13][93]  ( .CLK(n3478), .D(n3418), .Q(
        \inq_ary[13][93] ) );
  LATCHX1_RVT \inq_ary_reg[14][93]  ( .CLK(n3477), .D(n3418), .Q(
        \inq_ary[14][93] ) );
  LATCHX1_RVT \inq_ary_reg[15][93]  ( .CLK(n3476), .D(n3418), .Q(
        \inq_ary[15][93] ) );
  LATCHX1_RVT \dout_reg[93]  ( .CLK(n3492), .D(N354), .Q(dout[93]) );
  LATCHX1_RVT \inq_ary_reg[0][92]  ( .CLK(n3491), .D(n3416), .Q(
        \inq_ary[0][92] ) );
  LATCHX1_RVT \inq_ary_reg[1][92]  ( .CLK(n3490), .D(n3416), .Q(
        \inq_ary[1][92] ) );
  LATCHX1_RVT \inq_ary_reg[2][92]  ( .CLK(n3489), .D(n3416), .Q(
        \inq_ary[2][92] ) );
  LATCHX1_RVT \inq_ary_reg[3][92]  ( .CLK(n3488), .D(n3416), .Q(
        \inq_ary[3][92] ) );
  LATCHX1_RVT \inq_ary_reg[4][92]  ( .CLK(n3487), .D(n3416), .Q(
        \inq_ary[4][92] ) );
  LATCHX1_RVT \inq_ary_reg[5][92]  ( .CLK(n3486), .D(n3416), .Q(
        \inq_ary[5][92] ) );
  LATCHX1_RVT \inq_ary_reg[6][92]  ( .CLK(n3485), .D(n3416), .Q(
        \inq_ary[6][92] ) );
  LATCHX1_RVT \inq_ary_reg[7][92]  ( .CLK(n3484), .D(n3416), .Q(
        \inq_ary[7][92] ) );
  LATCHX1_RVT \inq_ary_reg[8][92]  ( .CLK(n3483), .D(n3416), .Q(
        \inq_ary[8][92] ) );
  LATCHX1_RVT \inq_ary_reg[9][92]  ( .CLK(n3482), .D(n3416), .Q(
        \inq_ary[9][92] ) );
  LATCHX1_RVT \inq_ary_reg[10][92]  ( .CLK(n3481), .D(n3416), .Q(
        \inq_ary[10][92] ) );
  LATCHX1_RVT \inq_ary_reg[11][92]  ( .CLK(n3480), .D(n3416), .Q(
        \inq_ary[11][92] ) );
  LATCHX1_RVT \inq_ary_reg[12][92]  ( .CLK(n3479), .D(n3416), .Q(
        \inq_ary[12][92] ) );
  LATCHX1_RVT \inq_ary_reg[13][92]  ( .CLK(n3478), .D(n3416), .Q(
        \inq_ary[13][92] ) );
  LATCHX1_RVT \inq_ary_reg[14][92]  ( .CLK(n3477), .D(n3416), .Q(
        \inq_ary[14][92] ) );
  LATCHX1_RVT \inq_ary_reg[15][92]  ( .CLK(n3476), .D(n3416), .Q(
        \inq_ary[15][92] ) );
  LATCHX1_RVT \dout_reg[92]  ( .CLK(n3492), .D(N353), .Q(dout[92]) );
  LATCHX1_RVT \inq_ary_reg[0][91]  ( .CLK(n3491), .D(n3423), .Q(
        \inq_ary[0][91] ) );
  LATCHX1_RVT \inq_ary_reg[1][91]  ( .CLK(n3490), .D(n3423), .Q(
        \inq_ary[1][91] ) );
  LATCHX1_RVT \inq_ary_reg[2][91]  ( .CLK(n3489), .D(n3423), .Q(
        \inq_ary[2][91] ) );
  LATCHX1_RVT \inq_ary_reg[3][91]  ( .CLK(n3488), .D(n3423), .Q(
        \inq_ary[3][91] ) );
  LATCHX1_RVT \inq_ary_reg[4][91]  ( .CLK(n3487), .D(n3423), .Q(
        \inq_ary[4][91] ) );
  LATCHX1_RVT \inq_ary_reg[5][91]  ( .CLK(n3486), .D(n3423), .Q(
        \inq_ary[5][91] ) );
  LATCHX1_RVT \inq_ary_reg[6][91]  ( .CLK(n3485), .D(n3423), .Q(
        \inq_ary[6][91] ) );
  LATCHX1_RVT \inq_ary_reg[7][91]  ( .CLK(n3484), .D(n3423), .Q(
        \inq_ary[7][91] ) );
  LATCHX1_RVT \inq_ary_reg[8][91]  ( .CLK(n3483), .D(n3423), .Q(
        \inq_ary[8][91] ) );
  LATCHX1_RVT \inq_ary_reg[9][91]  ( .CLK(n3482), .D(n3423), .Q(
        \inq_ary[9][91] ) );
  LATCHX1_RVT \inq_ary_reg[10][91]  ( .CLK(n3481), .D(n3423), .Q(
        \inq_ary[10][91] ) );
  LATCHX1_RVT \inq_ary_reg[11][91]  ( .CLK(n3480), .D(n3423), .Q(
        \inq_ary[11][91] ) );
  LATCHX1_RVT \inq_ary_reg[12][91]  ( .CLK(n3479), .D(n3423), .Q(
        \inq_ary[12][91] ) );
  LATCHX1_RVT \inq_ary_reg[13][91]  ( .CLK(n3478), .D(n3423), .Q(
        \inq_ary[13][91] ) );
  LATCHX1_RVT \inq_ary_reg[14][91]  ( .CLK(n3477), .D(n3423), .Q(
        \inq_ary[14][91] ) );
  LATCHX1_RVT \inq_ary_reg[15][91]  ( .CLK(n3476), .D(n3423), .Q(
        \inq_ary[15][91] ) );
  LATCHX1_RVT \dout_reg[91]  ( .CLK(n3492), .D(N352), .Q(dout[91]) );
  LATCHX1_RVT \inq_ary_reg[0][90]  ( .CLK(n3491), .D(n3421), .Q(
        \inq_ary[0][90] ) );
  LATCHX1_RVT \inq_ary_reg[1][90]  ( .CLK(n3490), .D(n3421), .Q(
        \inq_ary[1][90] ) );
  LATCHX1_RVT \inq_ary_reg[2][90]  ( .CLK(n3489), .D(n3421), .Q(
        \inq_ary[2][90] ) );
  LATCHX1_RVT \inq_ary_reg[3][90]  ( .CLK(n3488), .D(n3421), .Q(
        \inq_ary[3][90] ) );
  LATCHX1_RVT \inq_ary_reg[4][90]  ( .CLK(n3487), .D(n3421), .Q(
        \inq_ary[4][90] ) );
  LATCHX1_RVT \inq_ary_reg[5][90]  ( .CLK(n3486), .D(n3421), .Q(
        \inq_ary[5][90] ) );
  LATCHX1_RVT \inq_ary_reg[6][90]  ( .CLK(n3485), .D(n3421), .Q(
        \inq_ary[6][90] ) );
  LATCHX1_RVT \inq_ary_reg[7][90]  ( .CLK(n3484), .D(n3421), .Q(
        \inq_ary[7][90] ) );
  LATCHX1_RVT \inq_ary_reg[8][90]  ( .CLK(n3483), .D(n3421), .Q(
        \inq_ary[8][90] ) );
  LATCHX1_RVT \inq_ary_reg[9][90]  ( .CLK(n3482), .D(n3421), .Q(
        \inq_ary[9][90] ) );
  LATCHX1_RVT \inq_ary_reg[10][90]  ( .CLK(n3481), .D(n3421), .Q(
        \inq_ary[10][90] ) );
  LATCHX1_RVT \inq_ary_reg[11][90]  ( .CLK(n3480), .D(n3421), .Q(
        \inq_ary[11][90] ) );
  LATCHX1_RVT \inq_ary_reg[12][90]  ( .CLK(n3479), .D(n3421), .Q(
        \inq_ary[12][90] ) );
  LATCHX1_RVT \inq_ary_reg[13][90]  ( .CLK(n3478), .D(n3421), .Q(
        \inq_ary[13][90] ) );
  LATCHX1_RVT \inq_ary_reg[14][90]  ( .CLK(n3477), .D(n3421), .Q(
        \inq_ary[14][90] ) );
  LATCHX1_RVT \inq_ary_reg[15][90]  ( .CLK(n3476), .D(n3421), .Q(
        \inq_ary[15][90] ) );
  LATCHX1_RVT \dout_reg[90]  ( .CLK(n3492), .D(N351), .Q(dout[90]) );
  LATCHX1_RVT \inq_ary_reg[0][89]  ( .CLK(n3491), .D(n3419), .Q(
        \inq_ary[0][89] ) );
  LATCHX1_RVT \inq_ary_reg[1][89]  ( .CLK(n3490), .D(n3419), .Q(
        \inq_ary[1][89] ) );
  LATCHX1_RVT \inq_ary_reg[2][89]  ( .CLK(n3489), .D(n3419), .Q(
        \inq_ary[2][89] ) );
  LATCHX1_RVT \inq_ary_reg[3][89]  ( .CLK(n3488), .D(n3419), .Q(
        \inq_ary[3][89] ) );
  LATCHX1_RVT \inq_ary_reg[4][89]  ( .CLK(n3487), .D(n3419), .Q(
        \inq_ary[4][89] ) );
  LATCHX1_RVT \inq_ary_reg[5][89]  ( .CLK(n3486), .D(n3419), .Q(
        \inq_ary[5][89] ) );
  LATCHX1_RVT \inq_ary_reg[6][89]  ( .CLK(n3485), .D(n3419), .Q(
        \inq_ary[6][89] ) );
  LATCHX1_RVT \inq_ary_reg[7][89]  ( .CLK(n3484), .D(n3419), .Q(
        \inq_ary[7][89] ) );
  LATCHX1_RVT \inq_ary_reg[8][89]  ( .CLK(n3483), .D(n3419), .Q(
        \inq_ary[8][89] ) );
  LATCHX1_RVT \inq_ary_reg[9][89]  ( .CLK(n3482), .D(n3419), .Q(
        \inq_ary[9][89] ) );
  LATCHX1_RVT \inq_ary_reg[10][89]  ( .CLK(n3481), .D(n3419), .Q(
        \inq_ary[10][89] ) );
  LATCHX1_RVT \inq_ary_reg[11][89]  ( .CLK(n3480), .D(n3419), .Q(
        \inq_ary[11][89] ) );
  LATCHX1_RVT \inq_ary_reg[12][89]  ( .CLK(n3479), .D(n3419), .Q(
        \inq_ary[12][89] ) );
  LATCHX1_RVT \inq_ary_reg[13][89]  ( .CLK(n3478), .D(n3419), .Q(
        \inq_ary[13][89] ) );
  LATCHX1_RVT \inq_ary_reg[14][89]  ( .CLK(n3477), .D(n3419), .Q(
        \inq_ary[14][89] ) );
  LATCHX1_RVT \inq_ary_reg[15][89]  ( .CLK(n3476), .D(n3419), .Q(
        \inq_ary[15][89] ) );
  LATCHX1_RVT \dout_reg[89]  ( .CLK(n3492), .D(N350), .Q(dout[89]) );
  LATCHX1_RVT \inq_ary_reg[0][88]  ( .CLK(n3491), .D(n3417), .Q(
        \inq_ary[0][88] ) );
  LATCHX1_RVT \inq_ary_reg[1][88]  ( .CLK(n3490), .D(n3417), .Q(
        \inq_ary[1][88] ) );
  LATCHX1_RVT \inq_ary_reg[2][88]  ( .CLK(n3489), .D(n3417), .Q(
        \inq_ary[2][88] ) );
  LATCHX1_RVT \inq_ary_reg[3][88]  ( .CLK(n3488), .D(n3417), .Q(
        \inq_ary[3][88] ) );
  LATCHX1_RVT \inq_ary_reg[4][88]  ( .CLK(n3487), .D(n3417), .Q(
        \inq_ary[4][88] ) );
  LATCHX1_RVT \inq_ary_reg[5][88]  ( .CLK(n3486), .D(n3417), .Q(
        \inq_ary[5][88] ) );
  LATCHX1_RVT \inq_ary_reg[6][88]  ( .CLK(n3485), .D(n3417), .Q(
        \inq_ary[6][88] ) );
  LATCHX1_RVT \inq_ary_reg[7][88]  ( .CLK(n3484), .D(n3417), .Q(
        \inq_ary[7][88] ) );
  LATCHX1_RVT \inq_ary_reg[8][88]  ( .CLK(n3483), .D(n3417), .Q(
        \inq_ary[8][88] ) );
  LATCHX1_RVT \inq_ary_reg[9][88]  ( .CLK(n3482), .D(n3417), .Q(
        \inq_ary[9][88] ) );
  LATCHX1_RVT \inq_ary_reg[10][88]  ( .CLK(n3481), .D(n3417), .Q(
        \inq_ary[10][88] ) );
  LATCHX1_RVT \inq_ary_reg[11][88]  ( .CLK(n3480), .D(n3417), .Q(
        \inq_ary[11][88] ) );
  LATCHX1_RVT \inq_ary_reg[12][88]  ( .CLK(n3479), .D(n3417), .Q(
        \inq_ary[12][88] ) );
  LATCHX1_RVT \inq_ary_reg[13][88]  ( .CLK(n3478), .D(n3417), .Q(
        \inq_ary[13][88] ) );
  LATCHX1_RVT \inq_ary_reg[14][88]  ( .CLK(n3477), .D(n3417), .Q(
        \inq_ary[14][88] ) );
  LATCHX1_RVT \inq_ary_reg[15][88]  ( .CLK(n3476), .D(n3417), .Q(
        \inq_ary[15][88] ) );
  LATCHX1_RVT \dout_reg[88]  ( .CLK(n3492), .D(N349), .Q(dout[88]) );
  LATCHX1_RVT \inq_ary_reg[0][87]  ( .CLK(n3491), .D(n3414), .Q(
        \inq_ary[0][87] ) );
  LATCHX1_RVT \inq_ary_reg[1][87]  ( .CLK(n3490), .D(n3414), .Q(
        \inq_ary[1][87] ) );
  LATCHX1_RVT \inq_ary_reg[2][87]  ( .CLK(n3489), .D(n3414), .Q(
        \inq_ary[2][87] ) );
  LATCHX1_RVT \inq_ary_reg[3][87]  ( .CLK(n3488), .D(n3414), .Q(
        \inq_ary[3][87] ) );
  LATCHX1_RVT \inq_ary_reg[4][87]  ( .CLK(n3487), .D(n3414), .Q(
        \inq_ary[4][87] ) );
  LATCHX1_RVT \inq_ary_reg[5][87]  ( .CLK(n3486), .D(n3414), .Q(
        \inq_ary[5][87] ) );
  LATCHX1_RVT \inq_ary_reg[6][87]  ( .CLK(n3485), .D(n3414), .Q(
        \inq_ary[6][87] ) );
  LATCHX1_RVT \inq_ary_reg[7][87]  ( .CLK(n3484), .D(n3414), .Q(
        \inq_ary[7][87] ) );
  LATCHX1_RVT \inq_ary_reg[8][87]  ( .CLK(n3483), .D(n3414), .Q(
        \inq_ary[8][87] ) );
  LATCHX1_RVT \inq_ary_reg[9][87]  ( .CLK(n3482), .D(n3414), .Q(
        \inq_ary[9][87] ) );
  LATCHX1_RVT \inq_ary_reg[10][87]  ( .CLK(n3481), .D(n3414), .Q(
        \inq_ary[10][87] ) );
  LATCHX1_RVT \inq_ary_reg[11][87]  ( .CLK(n3480), .D(n3414), .Q(
        \inq_ary[11][87] ) );
  LATCHX1_RVT \inq_ary_reg[12][87]  ( .CLK(n3479), .D(n3414), .Q(
        \inq_ary[12][87] ) );
  LATCHX1_RVT \inq_ary_reg[13][87]  ( .CLK(n3478), .D(n3414), .Q(
        \inq_ary[13][87] ) );
  LATCHX1_RVT \inq_ary_reg[14][87]  ( .CLK(n3477), .D(n3414), .Q(
        \inq_ary[14][87] ) );
  LATCHX1_RVT \inq_ary_reg[15][87]  ( .CLK(n3476), .D(n3414), .Q(
        \inq_ary[15][87] ) );
  LATCHX1_RVT \dout_reg[87]  ( .CLK(n3492), .D(N348), .Q(dout[87]) );
  LATCHX1_RVT \inq_ary_reg[0][86]  ( .CLK(n3491), .D(n3412), .Q(
        \inq_ary[0][86] ) );
  LATCHX1_RVT \inq_ary_reg[1][86]  ( .CLK(n3490), .D(n3412), .Q(
        \inq_ary[1][86] ) );
  LATCHX1_RVT \inq_ary_reg[2][86]  ( .CLK(n3489), .D(n3412), .Q(
        \inq_ary[2][86] ) );
  LATCHX1_RVT \inq_ary_reg[3][86]  ( .CLK(n3488), .D(n3412), .Q(
        \inq_ary[3][86] ) );
  LATCHX1_RVT \inq_ary_reg[4][86]  ( .CLK(n3487), .D(n3412), .Q(
        \inq_ary[4][86] ) );
  LATCHX1_RVT \inq_ary_reg[5][86]  ( .CLK(n3486), .D(n3412), .Q(
        \inq_ary[5][86] ) );
  LATCHX1_RVT \inq_ary_reg[6][86]  ( .CLK(n3485), .D(n3412), .Q(
        \inq_ary[6][86] ) );
  LATCHX1_RVT \inq_ary_reg[7][86]  ( .CLK(n3484), .D(n3412), .Q(
        \inq_ary[7][86] ) );
  LATCHX1_RVT \inq_ary_reg[8][86]  ( .CLK(n3483), .D(n3412), .Q(
        \inq_ary[8][86] ) );
  LATCHX1_RVT \inq_ary_reg[9][86]  ( .CLK(n3482), .D(n3412), .Q(
        \inq_ary[9][86] ) );
  LATCHX1_RVT \inq_ary_reg[10][86]  ( .CLK(n3481), .D(n3412), .Q(
        \inq_ary[10][86] ) );
  LATCHX1_RVT \inq_ary_reg[11][86]  ( .CLK(n3480), .D(n3412), .Q(
        \inq_ary[11][86] ) );
  LATCHX1_RVT \inq_ary_reg[12][86]  ( .CLK(n3479), .D(n3412), .Q(
        \inq_ary[12][86] ) );
  LATCHX1_RVT \inq_ary_reg[13][86]  ( .CLK(n3478), .D(n3412), .Q(
        \inq_ary[13][86] ) );
  LATCHX1_RVT \inq_ary_reg[14][86]  ( .CLK(n3477), .D(n3412), .Q(
        \inq_ary[14][86] ) );
  LATCHX1_RVT \inq_ary_reg[15][86]  ( .CLK(n3476), .D(n3412), .Q(
        \inq_ary[15][86] ) );
  LATCHX1_RVT \dout_reg[86]  ( .CLK(n3492), .D(N347), .Q(dout[86]) );
  LATCHX1_RVT \inq_ary_reg[0][85]  ( .CLK(n3491), .D(n3410), .Q(
        \inq_ary[0][85] ) );
  LATCHX1_RVT \inq_ary_reg[1][85]  ( .CLK(n3490), .D(n3410), .Q(
        \inq_ary[1][85] ) );
  LATCHX1_RVT \inq_ary_reg[2][85]  ( .CLK(n3489), .D(n3410), .Q(
        \inq_ary[2][85] ) );
  LATCHX1_RVT \inq_ary_reg[3][85]  ( .CLK(n3488), .D(n3410), .Q(
        \inq_ary[3][85] ) );
  LATCHX1_RVT \inq_ary_reg[4][85]  ( .CLK(n3487), .D(n3410), .Q(
        \inq_ary[4][85] ) );
  LATCHX1_RVT \inq_ary_reg[5][85]  ( .CLK(n3486), .D(n3410), .Q(
        \inq_ary[5][85] ) );
  LATCHX1_RVT \inq_ary_reg[6][85]  ( .CLK(n3485), .D(n3410), .Q(
        \inq_ary[6][85] ) );
  LATCHX1_RVT \inq_ary_reg[7][85]  ( .CLK(n3484), .D(n3410), .Q(
        \inq_ary[7][85] ) );
  LATCHX1_RVT \inq_ary_reg[8][85]  ( .CLK(n3483), .D(n3410), .Q(
        \inq_ary[8][85] ) );
  LATCHX1_RVT \inq_ary_reg[9][85]  ( .CLK(n3482), .D(n3410), .Q(
        \inq_ary[9][85] ) );
  LATCHX1_RVT \inq_ary_reg[10][85]  ( .CLK(n3481), .D(n3410), .Q(
        \inq_ary[10][85] ) );
  LATCHX1_RVT \inq_ary_reg[11][85]  ( .CLK(n3480), .D(n3410), .Q(
        \inq_ary[11][85] ) );
  LATCHX1_RVT \inq_ary_reg[12][85]  ( .CLK(n3479), .D(n3410), .Q(
        \inq_ary[12][85] ) );
  LATCHX1_RVT \inq_ary_reg[13][85]  ( .CLK(n3478), .D(n3410), .Q(
        \inq_ary[13][85] ) );
  LATCHX1_RVT \inq_ary_reg[14][85]  ( .CLK(n3477), .D(n3410), .Q(
        \inq_ary[14][85] ) );
  LATCHX1_RVT \inq_ary_reg[15][85]  ( .CLK(n3476), .D(n3410), .Q(
        \inq_ary[15][85] ) );
  LATCHX1_RVT \dout_reg[85]  ( .CLK(n3492), .D(N346), .Q(dout[85]) );
  LATCHX1_RVT \inq_ary_reg[0][84]  ( .CLK(n3491), .D(n3408), .Q(
        \inq_ary[0][84] ) );
  LATCHX1_RVT \inq_ary_reg[1][84]  ( .CLK(n3490), .D(n3408), .Q(
        \inq_ary[1][84] ) );
  LATCHX1_RVT \inq_ary_reg[2][84]  ( .CLK(n3489), .D(n3408), .Q(
        \inq_ary[2][84] ) );
  LATCHX1_RVT \inq_ary_reg[3][84]  ( .CLK(n3488), .D(n3408), .Q(
        \inq_ary[3][84] ) );
  LATCHX1_RVT \inq_ary_reg[4][84]  ( .CLK(n3487), .D(n3408), .Q(
        \inq_ary[4][84] ) );
  LATCHX1_RVT \inq_ary_reg[5][84]  ( .CLK(n3486), .D(n3408), .Q(
        \inq_ary[5][84] ) );
  LATCHX1_RVT \inq_ary_reg[6][84]  ( .CLK(n3485), .D(n3408), .Q(
        \inq_ary[6][84] ) );
  LATCHX1_RVT \inq_ary_reg[7][84]  ( .CLK(n3484), .D(n3408), .Q(
        \inq_ary[7][84] ) );
  LATCHX1_RVT \inq_ary_reg[8][84]  ( .CLK(n3483), .D(n3408), .Q(
        \inq_ary[8][84] ) );
  LATCHX1_RVT \inq_ary_reg[9][84]  ( .CLK(n3482), .D(n3408), .Q(
        \inq_ary[9][84] ) );
  LATCHX1_RVT \inq_ary_reg[10][84]  ( .CLK(n3481), .D(n3408), .Q(
        \inq_ary[10][84] ) );
  LATCHX1_RVT \inq_ary_reg[11][84]  ( .CLK(n3480), .D(n3408), .Q(
        \inq_ary[11][84] ) );
  LATCHX1_RVT \inq_ary_reg[12][84]  ( .CLK(n3479), .D(n3408), .Q(
        \inq_ary[12][84] ) );
  LATCHX1_RVT \inq_ary_reg[13][84]  ( .CLK(n3478), .D(n3408), .Q(
        \inq_ary[13][84] ) );
  LATCHX1_RVT \inq_ary_reg[14][84]  ( .CLK(n3477), .D(n3408), .Q(
        \inq_ary[14][84] ) );
  LATCHX1_RVT \inq_ary_reg[15][84]  ( .CLK(n3476), .D(n3408), .Q(
        \inq_ary[15][84] ) );
  LATCHX1_RVT \dout_reg[84]  ( .CLK(n3492), .D(N345), .Q(dout[84]) );
  LATCHX1_RVT \inq_ary_reg[0][83]  ( .CLK(n3491), .D(n3415), .Q(
        \inq_ary[0][83] ) );
  LATCHX1_RVT \inq_ary_reg[1][83]  ( .CLK(n3490), .D(n3415), .Q(
        \inq_ary[1][83] ) );
  LATCHX1_RVT \inq_ary_reg[2][83]  ( .CLK(n3489), .D(n3415), .Q(
        \inq_ary[2][83] ) );
  LATCHX1_RVT \inq_ary_reg[3][83]  ( .CLK(n3488), .D(n3415), .Q(
        \inq_ary[3][83] ) );
  LATCHX1_RVT \inq_ary_reg[4][83]  ( .CLK(n3487), .D(n3415), .Q(
        \inq_ary[4][83] ) );
  LATCHX1_RVT \inq_ary_reg[5][83]  ( .CLK(n3486), .D(n3415), .Q(
        \inq_ary[5][83] ) );
  LATCHX1_RVT \inq_ary_reg[6][83]  ( .CLK(n3485), .D(n3415), .Q(
        \inq_ary[6][83] ) );
  LATCHX1_RVT \inq_ary_reg[7][83]  ( .CLK(n3484), .D(n3415), .Q(
        \inq_ary[7][83] ) );
  LATCHX1_RVT \inq_ary_reg[8][83]  ( .CLK(n3483), .D(n3415), .Q(
        \inq_ary[8][83] ) );
  LATCHX1_RVT \inq_ary_reg[9][83]  ( .CLK(n3482), .D(n3415), .Q(
        \inq_ary[9][83] ) );
  LATCHX1_RVT \inq_ary_reg[10][83]  ( .CLK(n3481), .D(n3415), .Q(
        \inq_ary[10][83] ) );
  LATCHX1_RVT \inq_ary_reg[11][83]  ( .CLK(n3480), .D(n3415), .Q(
        \inq_ary[11][83] ) );
  LATCHX1_RVT \inq_ary_reg[12][83]  ( .CLK(n3479), .D(n3415), .Q(
        \inq_ary[12][83] ) );
  LATCHX1_RVT \inq_ary_reg[13][83]  ( .CLK(n3478), .D(n3415), .Q(
        \inq_ary[13][83] ) );
  LATCHX1_RVT \inq_ary_reg[14][83]  ( .CLK(n3477), .D(n3415), .Q(
        \inq_ary[14][83] ) );
  LATCHX1_RVT \inq_ary_reg[15][83]  ( .CLK(n3476), .D(n3415), .Q(
        \inq_ary[15][83] ) );
  LATCHX1_RVT \dout_reg[83]  ( .CLK(n3492), .D(N344), .Q(dout[83]) );
  LATCHX1_RVT \inq_ary_reg[0][82]  ( .CLK(n3491), .D(n3413), .Q(
        \inq_ary[0][82] ) );
  LATCHX1_RVT \inq_ary_reg[1][82]  ( .CLK(n3490), .D(n3413), .Q(
        \inq_ary[1][82] ) );
  LATCHX1_RVT \inq_ary_reg[2][82]  ( .CLK(n3489), .D(n3413), .Q(
        \inq_ary[2][82] ) );
  LATCHX1_RVT \inq_ary_reg[3][82]  ( .CLK(n3488), .D(n3413), .Q(
        \inq_ary[3][82] ) );
  LATCHX1_RVT \inq_ary_reg[4][82]  ( .CLK(n3487), .D(n3413), .Q(
        \inq_ary[4][82] ) );
  LATCHX1_RVT \inq_ary_reg[5][82]  ( .CLK(n3486), .D(n3413), .Q(
        \inq_ary[5][82] ) );
  LATCHX1_RVT \inq_ary_reg[6][82]  ( .CLK(n3485), .D(n3413), .Q(
        \inq_ary[6][82] ) );
  LATCHX1_RVT \inq_ary_reg[7][82]  ( .CLK(n3484), .D(n3413), .Q(
        \inq_ary[7][82] ) );
  LATCHX1_RVT \inq_ary_reg[8][82]  ( .CLK(n3483), .D(n3413), .Q(
        \inq_ary[8][82] ) );
  LATCHX1_RVT \inq_ary_reg[9][82]  ( .CLK(n3482), .D(n3413), .Q(
        \inq_ary[9][82] ) );
  LATCHX1_RVT \inq_ary_reg[10][82]  ( .CLK(n3481), .D(n3413), .Q(
        \inq_ary[10][82] ) );
  LATCHX1_RVT \inq_ary_reg[11][82]  ( .CLK(n3480), .D(n3413), .Q(
        \inq_ary[11][82] ) );
  LATCHX1_RVT \inq_ary_reg[12][82]  ( .CLK(n3479), .D(n3413), .Q(
        \inq_ary[12][82] ) );
  LATCHX1_RVT \inq_ary_reg[13][82]  ( .CLK(n3478), .D(n3413), .Q(
        \inq_ary[13][82] ) );
  LATCHX1_RVT \inq_ary_reg[14][82]  ( .CLK(n3477), .D(n3413), .Q(
        \inq_ary[14][82] ) );
  LATCHX1_RVT \inq_ary_reg[15][82]  ( .CLK(n3476), .D(n3413), .Q(
        \inq_ary[15][82] ) );
  LATCHX1_RVT \dout_reg[82]  ( .CLK(n3492), .D(N343), .Q(dout[82]) );
  LATCHX1_RVT \inq_ary_reg[0][81]  ( .CLK(n3491), .D(n3411), .Q(
        \inq_ary[0][81] ) );
  LATCHX1_RVT \inq_ary_reg[1][81]  ( .CLK(n3490), .D(n3411), .Q(
        \inq_ary[1][81] ) );
  LATCHX1_RVT \inq_ary_reg[2][81]  ( .CLK(n3489), .D(n3411), .Q(
        \inq_ary[2][81] ) );
  LATCHX1_RVT \inq_ary_reg[3][81]  ( .CLK(n3488), .D(n3411), .Q(
        \inq_ary[3][81] ) );
  LATCHX1_RVT \inq_ary_reg[4][81]  ( .CLK(n3487), .D(n3411), .Q(
        \inq_ary[4][81] ) );
  LATCHX1_RVT \inq_ary_reg[5][81]  ( .CLK(n3486), .D(n3411), .Q(
        \inq_ary[5][81] ) );
  LATCHX1_RVT \inq_ary_reg[6][81]  ( .CLK(n3485), .D(n3411), .Q(
        \inq_ary[6][81] ) );
  LATCHX1_RVT \inq_ary_reg[7][81]  ( .CLK(n3484), .D(n3411), .Q(
        \inq_ary[7][81] ) );
  LATCHX1_RVT \inq_ary_reg[8][81]  ( .CLK(n3483), .D(n3411), .Q(
        \inq_ary[8][81] ) );
  LATCHX1_RVT \inq_ary_reg[9][81]  ( .CLK(n3482), .D(n3411), .Q(
        \inq_ary[9][81] ) );
  LATCHX1_RVT \inq_ary_reg[10][81]  ( .CLK(n3481), .D(n3411), .Q(
        \inq_ary[10][81] ) );
  LATCHX1_RVT \inq_ary_reg[11][81]  ( .CLK(n3480), .D(n3411), .Q(
        \inq_ary[11][81] ) );
  LATCHX1_RVT \inq_ary_reg[12][81]  ( .CLK(n3479), .D(n3411), .Q(
        \inq_ary[12][81] ) );
  LATCHX1_RVT \inq_ary_reg[13][81]  ( .CLK(n3478), .D(n3411), .Q(
        \inq_ary[13][81] ) );
  LATCHX1_RVT \inq_ary_reg[14][81]  ( .CLK(n3477), .D(n3411), .Q(
        \inq_ary[14][81] ) );
  LATCHX1_RVT \inq_ary_reg[15][81]  ( .CLK(n3476), .D(n3411), .Q(
        \inq_ary[15][81] ) );
  LATCHX1_RVT \dout_reg[81]  ( .CLK(n3492), .D(N342), .Q(dout[81]) );
  LATCHX1_RVT \inq_ary_reg[0][80]  ( .CLK(n3491), .D(n3409), .Q(
        \inq_ary[0][80] ) );
  LATCHX1_RVT \inq_ary_reg[1][80]  ( .CLK(n3490), .D(n3409), .Q(
        \inq_ary[1][80] ) );
  LATCHX1_RVT \inq_ary_reg[2][80]  ( .CLK(n3489), .D(n3409), .Q(
        \inq_ary[2][80] ) );
  LATCHX1_RVT \inq_ary_reg[3][80]  ( .CLK(n3488), .D(n3409), .Q(
        \inq_ary[3][80] ) );
  LATCHX1_RVT \inq_ary_reg[4][80]  ( .CLK(n3487), .D(n3409), .Q(
        \inq_ary[4][80] ) );
  LATCHX1_RVT \inq_ary_reg[5][80]  ( .CLK(n3486), .D(n3409), .Q(
        \inq_ary[5][80] ) );
  LATCHX1_RVT \inq_ary_reg[6][80]  ( .CLK(n3485), .D(n3409), .Q(
        \inq_ary[6][80] ) );
  LATCHX1_RVT \inq_ary_reg[7][80]  ( .CLK(n3484), .D(n3409), .Q(
        \inq_ary[7][80] ) );
  LATCHX1_RVT \inq_ary_reg[8][80]  ( .CLK(n3483), .D(n3409), .Q(
        \inq_ary[8][80] ) );
  LATCHX1_RVT \inq_ary_reg[9][80]  ( .CLK(n3482), .D(n3409), .Q(
        \inq_ary[9][80] ) );
  LATCHX1_RVT \inq_ary_reg[10][80]  ( .CLK(n3481), .D(n3409), .Q(
        \inq_ary[10][80] ) );
  LATCHX1_RVT \inq_ary_reg[11][80]  ( .CLK(n3480), .D(n3409), .Q(
        \inq_ary[11][80] ) );
  LATCHX1_RVT \inq_ary_reg[12][80]  ( .CLK(n3479), .D(n3409), .Q(
        \inq_ary[12][80] ) );
  LATCHX1_RVT \inq_ary_reg[13][80]  ( .CLK(n3478), .D(n3409), .Q(
        \inq_ary[13][80] ) );
  LATCHX1_RVT \inq_ary_reg[14][80]  ( .CLK(n3477), .D(n3409), .Q(
        \inq_ary[14][80] ) );
  LATCHX1_RVT \inq_ary_reg[15][80]  ( .CLK(n3476), .D(n3409), .Q(
        \inq_ary[15][80] ) );
  LATCHX1_RVT \dout_reg[80]  ( .CLK(n3492), .D(N341), .Q(dout[80]) );
  LATCHX1_RVT \inq_ary_reg[0][79]  ( .CLK(n3491), .D(n3406), .Q(
        \inq_ary[0][79] ) );
  LATCHX1_RVT \inq_ary_reg[1][79]  ( .CLK(n3490), .D(n3406), .Q(
        \inq_ary[1][79] ) );
  LATCHX1_RVT \inq_ary_reg[2][79]  ( .CLK(n3489), .D(n3406), .Q(
        \inq_ary[2][79] ) );
  LATCHX1_RVT \inq_ary_reg[3][79]  ( .CLK(n3488), .D(n3406), .Q(
        \inq_ary[3][79] ) );
  LATCHX1_RVT \inq_ary_reg[4][79]  ( .CLK(n3487), .D(n3406), .Q(
        \inq_ary[4][79] ) );
  LATCHX1_RVT \inq_ary_reg[5][79]  ( .CLK(n3486), .D(n3406), .Q(
        \inq_ary[5][79] ) );
  LATCHX1_RVT \inq_ary_reg[6][79]  ( .CLK(n3485), .D(n3406), .Q(
        \inq_ary[6][79] ) );
  LATCHX1_RVT \inq_ary_reg[7][79]  ( .CLK(n3484), .D(n3406), .Q(
        \inq_ary[7][79] ) );
  LATCHX1_RVT \inq_ary_reg[8][79]  ( .CLK(n3483), .D(n3406), .Q(
        \inq_ary[8][79] ) );
  LATCHX1_RVT \inq_ary_reg[9][79]  ( .CLK(n3482), .D(n3406), .Q(
        \inq_ary[9][79] ) );
  LATCHX1_RVT \inq_ary_reg[10][79]  ( .CLK(n3481), .D(n3406), .Q(
        \inq_ary[10][79] ) );
  LATCHX1_RVT \inq_ary_reg[11][79]  ( .CLK(n3480), .D(n3406), .Q(
        \inq_ary[11][79] ) );
  LATCHX1_RVT \inq_ary_reg[12][79]  ( .CLK(n3479), .D(n3406), .Q(
        \inq_ary[12][79] ) );
  LATCHX1_RVT \inq_ary_reg[13][79]  ( .CLK(n3478), .D(n3406), .Q(
        \inq_ary[13][79] ) );
  LATCHX1_RVT \inq_ary_reg[14][79]  ( .CLK(n3477), .D(n3406), .Q(
        \inq_ary[14][79] ) );
  LATCHX1_RVT \inq_ary_reg[15][79]  ( .CLK(n3476), .D(n3406), .Q(
        \inq_ary[15][79] ) );
  LATCHX1_RVT \dout_reg[79]  ( .CLK(n3492), .D(N340), .Q(dout[79]) );
  LATCHX1_RVT \inq_ary_reg[0][78]  ( .CLK(n3491), .D(n3404), .Q(
        \inq_ary[0][78] ) );
  LATCHX1_RVT \inq_ary_reg[1][78]  ( .CLK(n3490), .D(n3404), .Q(
        \inq_ary[1][78] ) );
  LATCHX1_RVT \inq_ary_reg[2][78]  ( .CLK(n3489), .D(n3404), .Q(
        \inq_ary[2][78] ) );
  LATCHX1_RVT \inq_ary_reg[3][78]  ( .CLK(n3488), .D(n3404), .Q(
        \inq_ary[3][78] ) );
  LATCHX1_RVT \inq_ary_reg[4][78]  ( .CLK(n3487), .D(n3404), .Q(
        \inq_ary[4][78] ) );
  LATCHX1_RVT \inq_ary_reg[5][78]  ( .CLK(n3486), .D(n3404), .Q(
        \inq_ary[5][78] ) );
  LATCHX1_RVT \inq_ary_reg[6][78]  ( .CLK(n3485), .D(n3404), .Q(
        \inq_ary[6][78] ) );
  LATCHX1_RVT \inq_ary_reg[7][78]  ( .CLK(n3484), .D(n3404), .Q(
        \inq_ary[7][78] ) );
  LATCHX1_RVT \inq_ary_reg[8][78]  ( .CLK(n3483), .D(n3404), .Q(
        \inq_ary[8][78] ) );
  LATCHX1_RVT \inq_ary_reg[9][78]  ( .CLK(n3482), .D(n3404), .Q(
        \inq_ary[9][78] ) );
  LATCHX1_RVT \inq_ary_reg[10][78]  ( .CLK(n3481), .D(n3404), .Q(
        \inq_ary[10][78] ) );
  LATCHX1_RVT \inq_ary_reg[11][78]  ( .CLK(n3480), .D(n3404), .Q(
        \inq_ary[11][78] ) );
  LATCHX1_RVT \inq_ary_reg[12][78]  ( .CLK(n3479), .D(n3404), .Q(
        \inq_ary[12][78] ) );
  LATCHX1_RVT \inq_ary_reg[13][78]  ( .CLK(n3478), .D(n3404), .Q(
        \inq_ary[13][78] ) );
  LATCHX1_RVT \inq_ary_reg[14][78]  ( .CLK(n3477), .D(n3404), .Q(
        \inq_ary[14][78] ) );
  LATCHX1_RVT \inq_ary_reg[15][78]  ( .CLK(n3476), .D(n3404), .Q(
        \inq_ary[15][78] ) );
  LATCHX1_RVT \dout_reg[78]  ( .CLK(n3492), .D(N339), .Q(dout[78]) );
  LATCHX1_RVT \inq_ary_reg[0][77]  ( .CLK(n3491), .D(n3402), .Q(
        \inq_ary[0][77] ) );
  LATCHX1_RVT \inq_ary_reg[1][77]  ( .CLK(n3490), .D(n3402), .Q(
        \inq_ary[1][77] ) );
  LATCHX1_RVT \inq_ary_reg[2][77]  ( .CLK(n3489), .D(n3402), .Q(
        \inq_ary[2][77] ) );
  LATCHX1_RVT \inq_ary_reg[3][77]  ( .CLK(n3488), .D(n3402), .Q(
        \inq_ary[3][77] ) );
  LATCHX1_RVT \inq_ary_reg[4][77]  ( .CLK(n3487), .D(n3402), .Q(
        \inq_ary[4][77] ) );
  LATCHX1_RVT \inq_ary_reg[5][77]  ( .CLK(n3486), .D(n3402), .Q(
        \inq_ary[5][77] ) );
  LATCHX1_RVT \inq_ary_reg[6][77]  ( .CLK(n3485), .D(n3402), .Q(
        \inq_ary[6][77] ) );
  LATCHX1_RVT \inq_ary_reg[7][77]  ( .CLK(n3484), .D(n3402), .Q(
        \inq_ary[7][77] ) );
  LATCHX1_RVT \inq_ary_reg[8][77]  ( .CLK(n3483), .D(n3402), .Q(
        \inq_ary[8][77] ) );
  LATCHX1_RVT \inq_ary_reg[9][77]  ( .CLK(n3482), .D(n3402), .Q(
        \inq_ary[9][77] ) );
  LATCHX1_RVT \inq_ary_reg[10][77]  ( .CLK(n3481), .D(n3402), .Q(
        \inq_ary[10][77] ) );
  LATCHX1_RVT \inq_ary_reg[11][77]  ( .CLK(n3480), .D(n3402), .Q(
        \inq_ary[11][77] ) );
  LATCHX1_RVT \inq_ary_reg[12][77]  ( .CLK(n3479), .D(n3402), .Q(
        \inq_ary[12][77] ) );
  LATCHX1_RVT \inq_ary_reg[13][77]  ( .CLK(n3478), .D(n3402), .Q(
        \inq_ary[13][77] ) );
  LATCHX1_RVT \inq_ary_reg[14][77]  ( .CLK(n3477), .D(n3402), .Q(
        \inq_ary[14][77] ) );
  LATCHX1_RVT \inq_ary_reg[15][77]  ( .CLK(n3476), .D(n3402), .Q(
        \inq_ary[15][77] ) );
  LATCHX1_RVT \dout_reg[77]  ( .CLK(n3492), .D(N338), .Q(dout[77]) );
  LATCHX1_RVT \inq_ary_reg[0][76]  ( .CLK(n3491), .D(n3400), .Q(
        \inq_ary[0][76] ) );
  LATCHX1_RVT \inq_ary_reg[1][76]  ( .CLK(n3490), .D(n3400), .Q(
        \inq_ary[1][76] ) );
  LATCHX1_RVT \inq_ary_reg[2][76]  ( .CLK(n3489), .D(n3400), .Q(
        \inq_ary[2][76] ) );
  LATCHX1_RVT \inq_ary_reg[3][76]  ( .CLK(n3488), .D(n3400), .Q(
        \inq_ary[3][76] ) );
  LATCHX1_RVT \inq_ary_reg[4][76]  ( .CLK(n3487), .D(n3400), .Q(
        \inq_ary[4][76] ) );
  LATCHX1_RVT \inq_ary_reg[5][76]  ( .CLK(n3486), .D(n3400), .Q(
        \inq_ary[5][76] ) );
  LATCHX1_RVT \inq_ary_reg[6][76]  ( .CLK(n3485), .D(n3400), .Q(
        \inq_ary[6][76] ) );
  LATCHX1_RVT \inq_ary_reg[7][76]  ( .CLK(n3484), .D(n3400), .Q(
        \inq_ary[7][76] ) );
  LATCHX1_RVT \inq_ary_reg[8][76]  ( .CLK(n3483), .D(n3400), .Q(
        \inq_ary[8][76] ) );
  LATCHX1_RVT \inq_ary_reg[9][76]  ( .CLK(n3482), .D(n3400), .Q(
        \inq_ary[9][76] ) );
  LATCHX1_RVT \inq_ary_reg[10][76]  ( .CLK(n3481), .D(n3400), .Q(
        \inq_ary[10][76] ) );
  LATCHX1_RVT \inq_ary_reg[11][76]  ( .CLK(n3480), .D(n3400), .Q(
        \inq_ary[11][76] ) );
  LATCHX1_RVT \inq_ary_reg[12][76]  ( .CLK(n3479), .D(n3400), .Q(
        \inq_ary[12][76] ) );
  LATCHX1_RVT \inq_ary_reg[13][76]  ( .CLK(n3478), .D(n3400), .Q(
        \inq_ary[13][76] ) );
  LATCHX1_RVT \inq_ary_reg[14][76]  ( .CLK(n3477), .D(n3400), .Q(
        \inq_ary[14][76] ) );
  LATCHX1_RVT \inq_ary_reg[15][76]  ( .CLK(n3476), .D(n3400), .Q(
        \inq_ary[15][76] ) );
  LATCHX1_RVT \dout_reg[76]  ( .CLK(n3492), .D(N337), .Q(dout[76]) );
  LATCHX1_RVT \inq_ary_reg[0][75]  ( .CLK(n3491), .D(n3407), .Q(
        \inq_ary[0][75] ) );
  LATCHX1_RVT \inq_ary_reg[1][75]  ( .CLK(n3490), .D(n3407), .Q(
        \inq_ary[1][75] ) );
  LATCHX1_RVT \inq_ary_reg[2][75]  ( .CLK(n3489), .D(n3407), .Q(
        \inq_ary[2][75] ) );
  LATCHX1_RVT \inq_ary_reg[3][75]  ( .CLK(n3488), .D(n3407), .Q(
        \inq_ary[3][75] ) );
  LATCHX1_RVT \inq_ary_reg[4][75]  ( .CLK(n3487), .D(n3407), .Q(
        \inq_ary[4][75] ) );
  LATCHX1_RVT \inq_ary_reg[5][75]  ( .CLK(n3486), .D(n3407), .Q(
        \inq_ary[5][75] ) );
  LATCHX1_RVT \inq_ary_reg[6][75]  ( .CLK(n3485), .D(n3407), .Q(
        \inq_ary[6][75] ) );
  LATCHX1_RVT \inq_ary_reg[7][75]  ( .CLK(n3484), .D(n3407), .Q(
        \inq_ary[7][75] ) );
  LATCHX1_RVT \inq_ary_reg[8][75]  ( .CLK(n3483), .D(n3407), .Q(
        \inq_ary[8][75] ) );
  LATCHX1_RVT \inq_ary_reg[9][75]  ( .CLK(n3482), .D(n3407), .Q(
        \inq_ary[9][75] ) );
  LATCHX1_RVT \inq_ary_reg[10][75]  ( .CLK(n3481), .D(n3407), .Q(
        \inq_ary[10][75] ) );
  LATCHX1_RVT \inq_ary_reg[11][75]  ( .CLK(n3480), .D(n3407), .Q(
        \inq_ary[11][75] ) );
  LATCHX1_RVT \inq_ary_reg[12][75]  ( .CLK(n3479), .D(n3407), .Q(
        \inq_ary[12][75] ) );
  LATCHX1_RVT \inq_ary_reg[13][75]  ( .CLK(n3478), .D(n3407), .Q(
        \inq_ary[13][75] ) );
  LATCHX1_RVT \inq_ary_reg[14][75]  ( .CLK(n3477), .D(n3407), .Q(
        \inq_ary[14][75] ) );
  LATCHX1_RVT \inq_ary_reg[15][75]  ( .CLK(n3476), .D(n3407), .Q(
        \inq_ary[15][75] ) );
  LATCHX1_RVT \dout_reg[75]  ( .CLK(n3492), .D(N336), .Q(dout[75]) );
  LATCHX1_RVT \inq_ary_reg[0][74]  ( .CLK(n3491), .D(n3405), .Q(
        \inq_ary[0][74] ) );
  LATCHX1_RVT \inq_ary_reg[1][74]  ( .CLK(n3490), .D(n3405), .Q(
        \inq_ary[1][74] ) );
  LATCHX1_RVT \inq_ary_reg[2][74]  ( .CLK(n3489), .D(n3405), .Q(
        \inq_ary[2][74] ) );
  LATCHX1_RVT \inq_ary_reg[3][74]  ( .CLK(n3488), .D(n3405), .Q(
        \inq_ary[3][74] ) );
  LATCHX1_RVT \inq_ary_reg[4][74]  ( .CLK(n3487), .D(n3405), .Q(
        \inq_ary[4][74] ) );
  LATCHX1_RVT \inq_ary_reg[5][74]  ( .CLK(n3486), .D(n3405), .Q(
        \inq_ary[5][74] ) );
  LATCHX1_RVT \inq_ary_reg[6][74]  ( .CLK(n3485), .D(n3405), .Q(
        \inq_ary[6][74] ) );
  LATCHX1_RVT \inq_ary_reg[7][74]  ( .CLK(n3484), .D(n3405), .Q(
        \inq_ary[7][74] ) );
  LATCHX1_RVT \inq_ary_reg[8][74]  ( .CLK(n3483), .D(n3405), .Q(
        \inq_ary[8][74] ) );
  LATCHX1_RVT \inq_ary_reg[9][74]  ( .CLK(n3482), .D(n3405), .Q(
        \inq_ary[9][74] ) );
  LATCHX1_RVT \inq_ary_reg[10][74]  ( .CLK(n3481), .D(n3405), .Q(
        \inq_ary[10][74] ) );
  LATCHX1_RVT \inq_ary_reg[11][74]  ( .CLK(n3480), .D(n3405), .Q(
        \inq_ary[11][74] ) );
  LATCHX1_RVT \inq_ary_reg[12][74]  ( .CLK(n3479), .D(n3405), .Q(
        \inq_ary[12][74] ) );
  LATCHX1_RVT \inq_ary_reg[13][74]  ( .CLK(n3478), .D(n3405), .Q(
        \inq_ary[13][74] ) );
  LATCHX1_RVT \inq_ary_reg[14][74]  ( .CLK(n3477), .D(n3405), .Q(
        \inq_ary[14][74] ) );
  LATCHX1_RVT \inq_ary_reg[15][74]  ( .CLK(n3476), .D(n3405), .Q(
        \inq_ary[15][74] ) );
  LATCHX1_RVT \dout_reg[74]  ( .CLK(n3492), .D(N335), .Q(dout[74]) );
  LATCHX1_RVT \inq_ary_reg[0][73]  ( .CLK(n3491), .D(n3403), .Q(
        \inq_ary[0][73] ) );
  LATCHX1_RVT \inq_ary_reg[1][73]  ( .CLK(n3490), .D(n3403), .Q(
        \inq_ary[1][73] ) );
  LATCHX1_RVT \inq_ary_reg[2][73]  ( .CLK(n3489), .D(n3403), .Q(
        \inq_ary[2][73] ) );
  LATCHX1_RVT \inq_ary_reg[3][73]  ( .CLK(n3488), .D(n3403), .Q(
        \inq_ary[3][73] ) );
  LATCHX1_RVT \inq_ary_reg[4][73]  ( .CLK(n3487), .D(n3403), .Q(
        \inq_ary[4][73] ) );
  LATCHX1_RVT \inq_ary_reg[5][73]  ( .CLK(n3486), .D(n3403), .Q(
        \inq_ary[5][73] ) );
  LATCHX1_RVT \inq_ary_reg[6][73]  ( .CLK(n3485), .D(n3403), .Q(
        \inq_ary[6][73] ) );
  LATCHX1_RVT \inq_ary_reg[7][73]  ( .CLK(n3484), .D(n3403), .Q(
        \inq_ary[7][73] ) );
  LATCHX1_RVT \inq_ary_reg[8][73]  ( .CLK(n3483), .D(n3403), .Q(
        \inq_ary[8][73] ) );
  LATCHX1_RVT \inq_ary_reg[9][73]  ( .CLK(n3482), .D(n3403), .Q(
        \inq_ary[9][73] ) );
  LATCHX1_RVT \inq_ary_reg[10][73]  ( .CLK(n3481), .D(n3403), .Q(
        \inq_ary[10][73] ) );
  LATCHX1_RVT \inq_ary_reg[11][73]  ( .CLK(n3480), .D(n3403), .Q(
        \inq_ary[11][73] ) );
  LATCHX1_RVT \inq_ary_reg[12][73]  ( .CLK(n3479), .D(n3403), .Q(
        \inq_ary[12][73] ) );
  LATCHX1_RVT \inq_ary_reg[13][73]  ( .CLK(n3478), .D(n3403), .Q(
        \inq_ary[13][73] ) );
  LATCHX1_RVT \inq_ary_reg[14][73]  ( .CLK(n3477), .D(n3403), .Q(
        \inq_ary[14][73] ) );
  LATCHX1_RVT \inq_ary_reg[15][73]  ( .CLK(n3476), .D(n3403), .Q(
        \inq_ary[15][73] ) );
  LATCHX1_RVT \dout_reg[73]  ( .CLK(n3492), .D(N334), .Q(dout[73]) );
  LATCHX1_RVT \inq_ary_reg[0][72]  ( .CLK(n3491), .D(n3401), .Q(
        \inq_ary[0][72] ) );
  LATCHX1_RVT \inq_ary_reg[1][72]  ( .CLK(n3490), .D(n3401), .Q(
        \inq_ary[1][72] ) );
  LATCHX1_RVT \inq_ary_reg[2][72]  ( .CLK(n3489), .D(n3401), .Q(
        \inq_ary[2][72] ) );
  LATCHX1_RVT \inq_ary_reg[3][72]  ( .CLK(n3488), .D(n3401), .Q(
        \inq_ary[3][72] ) );
  LATCHX1_RVT \inq_ary_reg[4][72]  ( .CLK(n3487), .D(n3401), .Q(
        \inq_ary[4][72] ) );
  LATCHX1_RVT \inq_ary_reg[5][72]  ( .CLK(n3486), .D(n3401), .Q(
        \inq_ary[5][72] ) );
  LATCHX1_RVT \inq_ary_reg[6][72]  ( .CLK(n3485), .D(n3401), .Q(
        \inq_ary[6][72] ) );
  LATCHX1_RVT \inq_ary_reg[7][72]  ( .CLK(n3484), .D(n3401), .Q(
        \inq_ary[7][72] ) );
  LATCHX1_RVT \inq_ary_reg[8][72]  ( .CLK(n3483), .D(n3401), .Q(
        \inq_ary[8][72] ) );
  LATCHX1_RVT \inq_ary_reg[9][72]  ( .CLK(n3482), .D(n3401), .Q(
        \inq_ary[9][72] ) );
  LATCHX1_RVT \inq_ary_reg[10][72]  ( .CLK(n3481), .D(n3401), .Q(
        \inq_ary[10][72] ) );
  LATCHX1_RVT \inq_ary_reg[11][72]  ( .CLK(n3480), .D(n3401), .Q(
        \inq_ary[11][72] ) );
  LATCHX1_RVT \inq_ary_reg[12][72]  ( .CLK(n3479), .D(n3401), .Q(
        \inq_ary[12][72] ) );
  LATCHX1_RVT \inq_ary_reg[13][72]  ( .CLK(n3478), .D(n3401), .Q(
        \inq_ary[13][72] ) );
  LATCHX1_RVT \inq_ary_reg[14][72]  ( .CLK(n3477), .D(n3401), .Q(
        \inq_ary[14][72] ) );
  LATCHX1_RVT \inq_ary_reg[15][72]  ( .CLK(n3476), .D(n3401), .Q(
        \inq_ary[15][72] ) );
  LATCHX1_RVT \dout_reg[72]  ( .CLK(n3492), .D(N333), .Q(dout[72]) );
  LATCHX1_RVT \inq_ary_reg[0][71]  ( .CLK(n3491), .D(n3398), .Q(
        \inq_ary[0][71] ) );
  LATCHX1_RVT \inq_ary_reg[1][71]  ( .CLK(n3490), .D(n3398), .Q(
        \inq_ary[1][71] ) );
  LATCHX1_RVT \inq_ary_reg[2][71]  ( .CLK(n3489), .D(n3398), .Q(
        \inq_ary[2][71] ) );
  LATCHX1_RVT \inq_ary_reg[3][71]  ( .CLK(n3488), .D(n3398), .Q(
        \inq_ary[3][71] ) );
  LATCHX1_RVT \inq_ary_reg[4][71]  ( .CLK(n3487), .D(n3398), .Q(
        \inq_ary[4][71] ) );
  LATCHX1_RVT \inq_ary_reg[5][71]  ( .CLK(n3486), .D(n3398), .Q(
        \inq_ary[5][71] ) );
  LATCHX1_RVT \inq_ary_reg[6][71]  ( .CLK(n3485), .D(n3398), .Q(
        \inq_ary[6][71] ) );
  LATCHX1_RVT \inq_ary_reg[7][71]  ( .CLK(n3484), .D(n3398), .Q(
        \inq_ary[7][71] ) );
  LATCHX1_RVT \inq_ary_reg[8][71]  ( .CLK(n3483), .D(n3398), .Q(
        \inq_ary[8][71] ) );
  LATCHX1_RVT \inq_ary_reg[9][71]  ( .CLK(n3482), .D(n3398), .Q(
        \inq_ary[9][71] ) );
  LATCHX1_RVT \inq_ary_reg[10][71]  ( .CLK(n3481), .D(n3398), .Q(
        \inq_ary[10][71] ) );
  LATCHX1_RVT \inq_ary_reg[11][71]  ( .CLK(n3480), .D(n3398), .Q(
        \inq_ary[11][71] ) );
  LATCHX1_RVT \inq_ary_reg[12][71]  ( .CLK(n3479), .D(n3398), .Q(
        \inq_ary[12][71] ) );
  LATCHX1_RVT \inq_ary_reg[13][71]  ( .CLK(n3478), .D(n3398), .Q(
        \inq_ary[13][71] ) );
  LATCHX1_RVT \inq_ary_reg[14][71]  ( .CLK(n3477), .D(n3398), .Q(
        \inq_ary[14][71] ) );
  LATCHX1_RVT \inq_ary_reg[15][71]  ( .CLK(n3476), .D(n3398), .Q(
        \inq_ary[15][71] ) );
  LATCHX1_RVT \dout_reg[71]  ( .CLK(n3492), .D(N332), .Q(dout[71]) );
  LATCHX1_RVT \inq_ary_reg[0][70]  ( .CLK(n3491), .D(n3396), .Q(
        \inq_ary[0][70] ) );
  LATCHX1_RVT \inq_ary_reg[1][70]  ( .CLK(n3490), .D(n3396), .Q(
        \inq_ary[1][70] ) );
  LATCHX1_RVT \inq_ary_reg[2][70]  ( .CLK(n3489), .D(n3396), .Q(
        \inq_ary[2][70] ) );
  LATCHX1_RVT \inq_ary_reg[3][70]  ( .CLK(n3488), .D(n3396), .Q(
        \inq_ary[3][70] ) );
  LATCHX1_RVT \inq_ary_reg[4][70]  ( .CLK(n3487), .D(n3396), .Q(
        \inq_ary[4][70] ) );
  LATCHX1_RVT \inq_ary_reg[5][70]  ( .CLK(n3486), .D(n3396), .Q(
        \inq_ary[5][70] ) );
  LATCHX1_RVT \inq_ary_reg[6][70]  ( .CLK(n3485), .D(n3396), .Q(
        \inq_ary[6][70] ) );
  LATCHX1_RVT \inq_ary_reg[7][70]  ( .CLK(n3484), .D(n3396), .Q(
        \inq_ary[7][70] ) );
  LATCHX1_RVT \inq_ary_reg[8][70]  ( .CLK(n3483), .D(n3396), .Q(
        \inq_ary[8][70] ) );
  LATCHX1_RVT \inq_ary_reg[9][70]  ( .CLK(n3482), .D(n3396), .Q(
        \inq_ary[9][70] ) );
  LATCHX1_RVT \inq_ary_reg[10][70]  ( .CLK(n3481), .D(n3396), .Q(
        \inq_ary[10][70] ) );
  LATCHX1_RVT \inq_ary_reg[11][70]  ( .CLK(n3480), .D(n3396), .Q(
        \inq_ary[11][70] ) );
  LATCHX1_RVT \inq_ary_reg[12][70]  ( .CLK(n3479), .D(n3396), .Q(
        \inq_ary[12][70] ) );
  LATCHX1_RVT \inq_ary_reg[13][70]  ( .CLK(n3478), .D(n3396), .Q(
        \inq_ary[13][70] ) );
  LATCHX1_RVT \inq_ary_reg[14][70]  ( .CLK(n3477), .D(n3396), .Q(
        \inq_ary[14][70] ) );
  LATCHX1_RVT \inq_ary_reg[15][70]  ( .CLK(n3476), .D(n3396), .Q(
        \inq_ary[15][70] ) );
  LATCHX1_RVT \dout_reg[70]  ( .CLK(n3492), .D(N331), .Q(dout[70]) );
  LATCHX1_RVT \inq_ary_reg[0][69]  ( .CLK(n3491), .D(n3394), .Q(
        \inq_ary[0][69] ) );
  LATCHX1_RVT \inq_ary_reg[1][69]  ( .CLK(n3490), .D(n3394), .Q(
        \inq_ary[1][69] ) );
  LATCHX1_RVT \inq_ary_reg[2][69]  ( .CLK(n3489), .D(n3394), .Q(
        \inq_ary[2][69] ) );
  LATCHX1_RVT \inq_ary_reg[3][69]  ( .CLK(n3488), .D(n3394), .Q(
        \inq_ary[3][69] ) );
  LATCHX1_RVT \inq_ary_reg[4][69]  ( .CLK(n3487), .D(n3394), .Q(
        \inq_ary[4][69] ) );
  LATCHX1_RVT \inq_ary_reg[5][69]  ( .CLK(n3486), .D(n3394), .Q(
        \inq_ary[5][69] ) );
  LATCHX1_RVT \inq_ary_reg[6][69]  ( .CLK(n3485), .D(n3394), .Q(
        \inq_ary[6][69] ) );
  LATCHX1_RVT \inq_ary_reg[7][69]  ( .CLK(n3484), .D(n3394), .Q(
        \inq_ary[7][69] ) );
  LATCHX1_RVT \inq_ary_reg[8][69]  ( .CLK(n3483), .D(n3394), .Q(
        \inq_ary[8][69] ) );
  LATCHX1_RVT \inq_ary_reg[9][69]  ( .CLK(n3482), .D(n3394), .Q(
        \inq_ary[9][69] ) );
  LATCHX1_RVT \inq_ary_reg[10][69]  ( .CLK(n3481), .D(n3394), .Q(
        \inq_ary[10][69] ) );
  LATCHX1_RVT \inq_ary_reg[11][69]  ( .CLK(n3480), .D(n3394), .Q(
        \inq_ary[11][69] ) );
  LATCHX1_RVT \inq_ary_reg[12][69]  ( .CLK(n3479), .D(n3394), .Q(
        \inq_ary[12][69] ) );
  LATCHX1_RVT \inq_ary_reg[13][69]  ( .CLK(n3478), .D(n3394), .Q(
        \inq_ary[13][69] ) );
  LATCHX1_RVT \inq_ary_reg[14][69]  ( .CLK(n3477), .D(n3394), .Q(
        \inq_ary[14][69] ) );
  LATCHX1_RVT \inq_ary_reg[15][69]  ( .CLK(n3476), .D(n3394), .Q(
        \inq_ary[15][69] ) );
  LATCHX1_RVT \dout_reg[69]  ( .CLK(n3492), .D(N330), .Q(dout[69]) );
  LATCHX1_RVT \inq_ary_reg[0][68]  ( .CLK(n3491), .D(n3392), .Q(
        \inq_ary[0][68] ) );
  LATCHX1_RVT \inq_ary_reg[1][68]  ( .CLK(n3490), .D(n3392), .Q(
        \inq_ary[1][68] ) );
  LATCHX1_RVT \inq_ary_reg[2][68]  ( .CLK(n3489), .D(n3392), .Q(
        \inq_ary[2][68] ) );
  LATCHX1_RVT \inq_ary_reg[3][68]  ( .CLK(n3488), .D(n3392), .Q(
        \inq_ary[3][68] ) );
  LATCHX1_RVT \inq_ary_reg[4][68]  ( .CLK(n3487), .D(n3392), .Q(
        \inq_ary[4][68] ) );
  LATCHX1_RVT \inq_ary_reg[5][68]  ( .CLK(n3486), .D(n3392), .Q(
        \inq_ary[5][68] ) );
  LATCHX1_RVT \inq_ary_reg[6][68]  ( .CLK(n3485), .D(n3392), .Q(
        \inq_ary[6][68] ) );
  LATCHX1_RVT \inq_ary_reg[7][68]  ( .CLK(n3484), .D(n3392), .Q(
        \inq_ary[7][68] ) );
  LATCHX1_RVT \inq_ary_reg[8][68]  ( .CLK(n3483), .D(n3392), .Q(
        \inq_ary[8][68] ) );
  LATCHX1_RVT \inq_ary_reg[9][68]  ( .CLK(n3482), .D(n3392), .Q(
        \inq_ary[9][68] ) );
  LATCHX1_RVT \inq_ary_reg[10][68]  ( .CLK(n3481), .D(n3392), .Q(
        \inq_ary[10][68] ) );
  LATCHX1_RVT \inq_ary_reg[11][68]  ( .CLK(n3480), .D(n3392), .Q(
        \inq_ary[11][68] ) );
  LATCHX1_RVT \inq_ary_reg[12][68]  ( .CLK(n3479), .D(n3392), .Q(
        \inq_ary[12][68] ) );
  LATCHX1_RVT \inq_ary_reg[13][68]  ( .CLK(n3478), .D(n3392), .Q(
        \inq_ary[13][68] ) );
  LATCHX1_RVT \inq_ary_reg[14][68]  ( .CLK(n3477), .D(n3392), .Q(
        \inq_ary[14][68] ) );
  LATCHX1_RVT \inq_ary_reg[15][68]  ( .CLK(n3476), .D(n3392), .Q(
        \inq_ary[15][68] ) );
  LATCHX1_RVT \dout_reg[68]  ( .CLK(n3492), .D(N329), .Q(dout[68]) );
  LATCHX1_RVT \inq_ary_reg[0][67]  ( .CLK(n3491), .D(n3399), .Q(
        \inq_ary[0][67] ) );
  LATCHX1_RVT \inq_ary_reg[1][67]  ( .CLK(n3490), .D(n3399), .Q(
        \inq_ary[1][67] ) );
  LATCHX1_RVT \inq_ary_reg[2][67]  ( .CLK(n3489), .D(n3399), .Q(
        \inq_ary[2][67] ) );
  LATCHX1_RVT \inq_ary_reg[3][67]  ( .CLK(n3488), .D(n3399), .Q(
        \inq_ary[3][67] ) );
  LATCHX1_RVT \inq_ary_reg[4][67]  ( .CLK(n3487), .D(n3399), .Q(
        \inq_ary[4][67] ) );
  LATCHX1_RVT \inq_ary_reg[5][67]  ( .CLK(n3486), .D(n3399), .Q(
        \inq_ary[5][67] ) );
  LATCHX1_RVT \inq_ary_reg[6][67]  ( .CLK(n3485), .D(n3399), .Q(
        \inq_ary[6][67] ) );
  LATCHX1_RVT \inq_ary_reg[7][67]  ( .CLK(n3484), .D(n3399), .Q(
        \inq_ary[7][67] ) );
  LATCHX1_RVT \inq_ary_reg[8][67]  ( .CLK(n3483), .D(n3399), .Q(
        \inq_ary[8][67] ) );
  LATCHX1_RVT \inq_ary_reg[9][67]  ( .CLK(n3482), .D(n3399), .Q(
        \inq_ary[9][67] ) );
  LATCHX1_RVT \inq_ary_reg[10][67]  ( .CLK(n3481), .D(n3399), .Q(
        \inq_ary[10][67] ) );
  LATCHX1_RVT \inq_ary_reg[11][67]  ( .CLK(n3480), .D(n3399), .Q(
        \inq_ary[11][67] ) );
  LATCHX1_RVT \inq_ary_reg[12][67]  ( .CLK(n3479), .D(n3399), .Q(
        \inq_ary[12][67] ) );
  LATCHX1_RVT \inq_ary_reg[13][67]  ( .CLK(n3478), .D(n3399), .Q(
        \inq_ary[13][67] ) );
  LATCHX1_RVT \inq_ary_reg[14][67]  ( .CLK(n3477), .D(n3399), .Q(
        \inq_ary[14][67] ) );
  LATCHX1_RVT \inq_ary_reg[15][67]  ( .CLK(n3476), .D(n3399), .Q(
        \inq_ary[15][67] ) );
  LATCHX1_RVT \dout_reg[67]  ( .CLK(n3492), .D(N328), .Q(dout[67]) );
  LATCHX1_RVT \inq_ary_reg[0][66]  ( .CLK(n3491), .D(n3397), .Q(
        \inq_ary[0][66] ) );
  LATCHX1_RVT \inq_ary_reg[1][66]  ( .CLK(n3490), .D(n3397), .Q(
        \inq_ary[1][66] ) );
  LATCHX1_RVT \inq_ary_reg[2][66]  ( .CLK(n3489), .D(n3397), .Q(
        \inq_ary[2][66] ) );
  LATCHX1_RVT \inq_ary_reg[3][66]  ( .CLK(n3488), .D(n3397), .Q(
        \inq_ary[3][66] ) );
  LATCHX1_RVT \inq_ary_reg[4][66]  ( .CLK(n3487), .D(n3397), .Q(
        \inq_ary[4][66] ) );
  LATCHX1_RVT \inq_ary_reg[5][66]  ( .CLK(n3486), .D(n3397), .Q(
        \inq_ary[5][66] ) );
  LATCHX1_RVT \inq_ary_reg[6][66]  ( .CLK(n3485), .D(n3397), .Q(
        \inq_ary[6][66] ) );
  LATCHX1_RVT \inq_ary_reg[7][66]  ( .CLK(n3484), .D(n3397), .Q(
        \inq_ary[7][66] ) );
  LATCHX1_RVT \inq_ary_reg[8][66]  ( .CLK(n3483), .D(n3397), .Q(
        \inq_ary[8][66] ) );
  LATCHX1_RVT \inq_ary_reg[9][66]  ( .CLK(n3482), .D(n3397), .Q(
        \inq_ary[9][66] ) );
  LATCHX1_RVT \inq_ary_reg[10][66]  ( .CLK(n3481), .D(n3397), .Q(
        \inq_ary[10][66] ) );
  LATCHX1_RVT \inq_ary_reg[11][66]  ( .CLK(n3480), .D(n3397), .Q(
        \inq_ary[11][66] ) );
  LATCHX1_RVT \inq_ary_reg[12][66]  ( .CLK(n3479), .D(n3397), .Q(
        \inq_ary[12][66] ) );
  LATCHX1_RVT \inq_ary_reg[13][66]  ( .CLK(n3478), .D(n3397), .Q(
        \inq_ary[13][66] ) );
  LATCHX1_RVT \inq_ary_reg[14][66]  ( .CLK(n3477), .D(n3397), .Q(
        \inq_ary[14][66] ) );
  LATCHX1_RVT \inq_ary_reg[15][66]  ( .CLK(n3476), .D(n3397), .Q(
        \inq_ary[15][66] ) );
  LATCHX1_RVT \dout_reg[66]  ( .CLK(n3492), .D(N327), .Q(dout[66]) );
  LATCHX1_RVT \inq_ary_reg[0][65]  ( .CLK(n3491), .D(n3395), .Q(
        \inq_ary[0][65] ) );
  LATCHX1_RVT \inq_ary_reg[1][65]  ( .CLK(n3490), .D(n3395), .Q(
        \inq_ary[1][65] ) );
  LATCHX1_RVT \inq_ary_reg[2][65]  ( .CLK(n3489), .D(n3395), .Q(
        \inq_ary[2][65] ) );
  LATCHX1_RVT \inq_ary_reg[3][65]  ( .CLK(n3488), .D(n3395), .Q(
        \inq_ary[3][65] ) );
  LATCHX1_RVT \inq_ary_reg[4][65]  ( .CLK(n3487), .D(n3395), .Q(
        \inq_ary[4][65] ) );
  LATCHX1_RVT \inq_ary_reg[5][65]  ( .CLK(n3486), .D(n3395), .Q(
        \inq_ary[5][65] ) );
  LATCHX1_RVT \inq_ary_reg[6][65]  ( .CLK(n3485), .D(n3395), .Q(
        \inq_ary[6][65] ) );
  LATCHX1_RVT \inq_ary_reg[7][65]  ( .CLK(n3484), .D(n3395), .Q(
        \inq_ary[7][65] ) );
  LATCHX1_RVT \inq_ary_reg[8][65]  ( .CLK(n3483), .D(n3395), .Q(
        \inq_ary[8][65] ) );
  LATCHX1_RVT \inq_ary_reg[9][65]  ( .CLK(n3482), .D(n3395), .Q(
        \inq_ary[9][65] ) );
  LATCHX1_RVT \inq_ary_reg[10][65]  ( .CLK(n3481), .D(n3395), .Q(
        \inq_ary[10][65] ) );
  LATCHX1_RVT \inq_ary_reg[11][65]  ( .CLK(n3480), .D(n3395), .Q(
        \inq_ary[11][65] ) );
  LATCHX1_RVT \inq_ary_reg[12][65]  ( .CLK(n3479), .D(n3395), .Q(
        \inq_ary[12][65] ) );
  LATCHX1_RVT \inq_ary_reg[13][65]  ( .CLK(n3478), .D(n3395), .Q(
        \inq_ary[13][65] ) );
  LATCHX1_RVT \inq_ary_reg[14][65]  ( .CLK(n3477), .D(n3395), .Q(
        \inq_ary[14][65] ) );
  LATCHX1_RVT \inq_ary_reg[15][65]  ( .CLK(n3476), .D(n3395), .Q(
        \inq_ary[15][65] ) );
  LATCHX1_RVT \dout_reg[65]  ( .CLK(n3492), .D(N326), .Q(dout[65]) );
  LATCHX1_RVT \inq_ary_reg[0][64]  ( .CLK(n3491), .D(n3393), .Q(
        \inq_ary[0][64] ) );
  LATCHX1_RVT \inq_ary_reg[1][64]  ( .CLK(n3490), .D(n3393), .Q(
        \inq_ary[1][64] ) );
  LATCHX1_RVT \inq_ary_reg[2][64]  ( .CLK(n3489), .D(n3393), .Q(
        \inq_ary[2][64] ) );
  LATCHX1_RVT \inq_ary_reg[3][64]  ( .CLK(n3488), .D(n3393), .Q(
        \inq_ary[3][64] ) );
  LATCHX1_RVT \inq_ary_reg[4][64]  ( .CLK(n3487), .D(n3393), .Q(
        \inq_ary[4][64] ) );
  LATCHX1_RVT \inq_ary_reg[5][64]  ( .CLK(n3486), .D(n3393), .Q(
        \inq_ary[5][64] ) );
  LATCHX1_RVT \inq_ary_reg[6][64]  ( .CLK(n3485), .D(n3393), .Q(
        \inq_ary[6][64] ) );
  LATCHX1_RVT \inq_ary_reg[7][64]  ( .CLK(n3484), .D(n3393), .Q(
        \inq_ary[7][64] ) );
  LATCHX1_RVT \inq_ary_reg[8][64]  ( .CLK(n3483), .D(n3393), .Q(
        \inq_ary[8][64] ) );
  LATCHX1_RVT \inq_ary_reg[9][64]  ( .CLK(n3482), .D(n3393), .Q(
        \inq_ary[9][64] ) );
  LATCHX1_RVT \inq_ary_reg[10][64]  ( .CLK(n3481), .D(n3393), .Q(
        \inq_ary[10][64] ) );
  LATCHX1_RVT \inq_ary_reg[11][64]  ( .CLK(n3480), .D(n3393), .Q(
        \inq_ary[11][64] ) );
  LATCHX1_RVT \inq_ary_reg[12][64]  ( .CLK(n3479), .D(n3393), .Q(
        \inq_ary[12][64] ) );
  LATCHX1_RVT \inq_ary_reg[13][64]  ( .CLK(n3478), .D(n3393), .Q(
        \inq_ary[13][64] ) );
  LATCHX1_RVT \inq_ary_reg[14][64]  ( .CLK(n3477), .D(n3393), .Q(
        \inq_ary[14][64] ) );
  LATCHX1_RVT \inq_ary_reg[15][64]  ( .CLK(n3476), .D(n3393), .Q(
        \inq_ary[15][64] ) );
  LATCHX1_RVT \dout_reg[64]  ( .CLK(n3492), .D(N325), .Q(dout[64]) );
  LATCHX1_RVT \inq_ary_reg[0][63]  ( .CLK(n3491), .D(n1549), .Q(
        \inq_ary[0][63] ) );
  LATCHX1_RVT \inq_ary_reg[1][63]  ( .CLK(n3490), .D(n1549), .Q(
        \inq_ary[1][63] ) );
  LATCHX1_RVT \inq_ary_reg[2][63]  ( .CLK(n3489), .D(n1549), .Q(
        \inq_ary[2][63] ) );
  LATCHX1_RVT \inq_ary_reg[3][63]  ( .CLK(n3488), .D(n1549), .Q(
        \inq_ary[3][63] ) );
  LATCHX1_RVT \inq_ary_reg[4][63]  ( .CLK(n3487), .D(n1549), .Q(
        \inq_ary[4][63] ) );
  LATCHX1_RVT \inq_ary_reg[5][63]  ( .CLK(n3486), .D(n1549), .Q(
        \inq_ary[5][63] ) );
  LATCHX1_RVT \inq_ary_reg[6][63]  ( .CLK(n3485), .D(n1549), .Q(
        \inq_ary[6][63] ) );
  LATCHX1_RVT \inq_ary_reg[7][63]  ( .CLK(n3484), .D(n1549), .Q(
        \inq_ary[7][63] ) );
  LATCHX1_RVT \inq_ary_reg[8][63]  ( .CLK(n3483), .D(n1549), .Q(
        \inq_ary[8][63] ) );
  LATCHX1_RVT \inq_ary_reg[9][63]  ( .CLK(n3482), .D(n1549), .Q(
        \inq_ary[9][63] ) );
  LATCHX1_RVT \inq_ary_reg[10][63]  ( .CLK(n3481), .D(n1549), .Q(
        \inq_ary[10][63] ) );
  LATCHX1_RVT \inq_ary_reg[11][63]  ( .CLK(n3480), .D(n1549), .Q(
        \inq_ary[11][63] ) );
  LATCHX1_RVT \inq_ary_reg[12][63]  ( .CLK(n3479), .D(n1549), .Q(
        \inq_ary[12][63] ) );
  LATCHX1_RVT \inq_ary_reg[13][63]  ( .CLK(n3478), .D(n1549), .Q(
        \inq_ary[13][63] ) );
  LATCHX1_RVT \inq_ary_reg[14][63]  ( .CLK(n3477), .D(n1549), .Q(
        \inq_ary[14][63] ) );
  LATCHX1_RVT \inq_ary_reg[15][63]  ( .CLK(n3476), .D(n1549), .Q(
        \inq_ary[15][63] ) );
  LATCHX1_RVT \dout_reg[63]  ( .CLK(n3492), .D(N324), .Q(dout[63]) );
  LATCHX1_RVT \inq_ary_reg[0][62]  ( .CLK(n3491), .D(n1536), .Q(
        \inq_ary[0][62] ) );
  LATCHX1_RVT \inq_ary_reg[1][62]  ( .CLK(n3490), .D(n1536), .Q(
        \inq_ary[1][62] ) );
  LATCHX1_RVT \inq_ary_reg[2][62]  ( .CLK(n3489), .D(n1536), .Q(
        \inq_ary[2][62] ) );
  LATCHX1_RVT \inq_ary_reg[3][62]  ( .CLK(n3488), .D(n1536), .Q(
        \inq_ary[3][62] ) );
  LATCHX1_RVT \inq_ary_reg[4][62]  ( .CLK(n3487), .D(n1536), .Q(
        \inq_ary[4][62] ) );
  LATCHX1_RVT \inq_ary_reg[5][62]  ( .CLK(n3486), .D(n1536), .Q(
        \inq_ary[5][62] ) );
  LATCHX1_RVT \inq_ary_reg[6][62]  ( .CLK(n3485), .D(n1536), .Q(
        \inq_ary[6][62] ) );
  LATCHX1_RVT \inq_ary_reg[7][62]  ( .CLK(n3484), .D(n1536), .Q(
        \inq_ary[7][62] ) );
  LATCHX1_RVT \inq_ary_reg[8][62]  ( .CLK(n3483), .D(n1536), .Q(
        \inq_ary[8][62] ) );
  LATCHX1_RVT \inq_ary_reg[9][62]  ( .CLK(n3482), .D(n1536), .Q(
        \inq_ary[9][62] ) );
  LATCHX1_RVT \inq_ary_reg[10][62]  ( .CLK(n3481), .D(n1536), .Q(
        \inq_ary[10][62] ) );
  LATCHX1_RVT \inq_ary_reg[11][62]  ( .CLK(n3480), .D(n1536), .Q(
        \inq_ary[11][62] ) );
  LATCHX1_RVT \inq_ary_reg[12][62]  ( .CLK(n3479), .D(n1536), .Q(
        \inq_ary[12][62] ) );
  LATCHX1_RVT \inq_ary_reg[13][62]  ( .CLK(n3478), .D(n1536), .Q(
        \inq_ary[13][62] ) );
  LATCHX1_RVT \inq_ary_reg[14][62]  ( .CLK(n3477), .D(n1536), .Q(
        \inq_ary[14][62] ) );
  LATCHX1_RVT \inq_ary_reg[15][62]  ( .CLK(n3476), .D(n1536), .Q(
        \inq_ary[15][62] ) );
  LATCHX1_RVT \dout_reg[62]  ( .CLK(n3492), .D(N323), .Q(dout[62]) );
  LATCHX1_RVT \inq_ary_reg[0][61]  ( .CLK(n3491), .D(n3391), .Q(
        \inq_ary[0][61] ) );
  LATCHX1_RVT \inq_ary_reg[1][61]  ( .CLK(n3490), .D(n3391), .Q(
        \inq_ary[1][61] ) );
  LATCHX1_RVT \inq_ary_reg[2][61]  ( .CLK(n3489), .D(n3391), .Q(
        \inq_ary[2][61] ) );
  LATCHX1_RVT \inq_ary_reg[3][61]  ( .CLK(n3488), .D(n3391), .Q(
        \inq_ary[3][61] ) );
  LATCHX1_RVT \inq_ary_reg[4][61]  ( .CLK(n3487), .D(n3391), .Q(
        \inq_ary[4][61] ) );
  LATCHX1_RVT \inq_ary_reg[5][61]  ( .CLK(n3486), .D(n3391), .Q(
        \inq_ary[5][61] ) );
  LATCHX1_RVT \inq_ary_reg[6][61]  ( .CLK(n3485), .D(n3391), .Q(
        \inq_ary[6][61] ) );
  LATCHX1_RVT \inq_ary_reg[7][61]  ( .CLK(n3484), .D(n3391), .Q(
        \inq_ary[7][61] ) );
  LATCHX1_RVT \inq_ary_reg[8][61]  ( .CLK(n3483), .D(n3391), .Q(
        \inq_ary[8][61] ) );
  LATCHX1_RVT \inq_ary_reg[9][61]  ( .CLK(n3482), .D(n3391), .Q(
        \inq_ary[9][61] ) );
  LATCHX1_RVT \inq_ary_reg[10][61]  ( .CLK(n3481), .D(n3391), .Q(
        \inq_ary[10][61] ) );
  LATCHX1_RVT \inq_ary_reg[11][61]  ( .CLK(n3480), .D(n3391), .Q(
        \inq_ary[11][61] ) );
  LATCHX1_RVT \inq_ary_reg[12][61]  ( .CLK(n3479), .D(n3391), .Q(
        \inq_ary[12][61] ) );
  LATCHX1_RVT \inq_ary_reg[13][61]  ( .CLK(n3478), .D(n3391), .Q(
        \inq_ary[13][61] ) );
  LATCHX1_RVT \inq_ary_reg[14][61]  ( .CLK(n3477), .D(n3391), .Q(
        \inq_ary[14][61] ) );
  LATCHX1_RVT \inq_ary_reg[15][61]  ( .CLK(n3476), .D(n3391), .Q(
        \inq_ary[15][61] ) );
  LATCHX1_RVT \dout_reg[61]  ( .CLK(n3492), .D(N322), .Q(dout[61]) );
  LATCHX1_RVT \inq_ary_reg[0][60]  ( .CLK(n3491), .D(n3390), .Q(
        \inq_ary[0][60] ) );
  LATCHX1_RVT \inq_ary_reg[1][60]  ( .CLK(n3490), .D(n3390), .Q(
        \inq_ary[1][60] ) );
  LATCHX1_RVT \inq_ary_reg[2][60]  ( .CLK(n3489), .D(n3390), .Q(
        \inq_ary[2][60] ) );
  LATCHX1_RVT \inq_ary_reg[3][60]  ( .CLK(n3488), .D(n3390), .Q(
        \inq_ary[3][60] ) );
  LATCHX1_RVT \inq_ary_reg[4][60]  ( .CLK(n3487), .D(n3390), .Q(
        \inq_ary[4][60] ) );
  LATCHX1_RVT \inq_ary_reg[5][60]  ( .CLK(n3486), .D(n3390), .Q(
        \inq_ary[5][60] ) );
  LATCHX1_RVT \inq_ary_reg[6][60]  ( .CLK(n3485), .D(n3390), .Q(
        \inq_ary[6][60] ) );
  LATCHX1_RVT \inq_ary_reg[7][60]  ( .CLK(n3484), .D(n3390), .Q(
        \inq_ary[7][60] ) );
  LATCHX1_RVT \inq_ary_reg[8][60]  ( .CLK(n3483), .D(n3390), .Q(
        \inq_ary[8][60] ) );
  LATCHX1_RVT \inq_ary_reg[9][60]  ( .CLK(n3482), .D(n3390), .Q(
        \inq_ary[9][60] ) );
  LATCHX1_RVT \inq_ary_reg[10][60]  ( .CLK(n3481), .D(n3390), .Q(
        \inq_ary[10][60] ) );
  LATCHX1_RVT \inq_ary_reg[11][60]  ( .CLK(n3480), .D(n3390), .Q(
        \inq_ary[11][60] ) );
  LATCHX1_RVT \inq_ary_reg[12][60]  ( .CLK(n3479), .D(n3390), .Q(
        \inq_ary[12][60] ) );
  LATCHX1_RVT \inq_ary_reg[13][60]  ( .CLK(n3478), .D(n3390), .Q(
        \inq_ary[13][60] ) );
  LATCHX1_RVT \inq_ary_reg[14][60]  ( .CLK(n3477), .D(n3390), .Q(
        \inq_ary[14][60] ) );
  LATCHX1_RVT \inq_ary_reg[15][60]  ( .CLK(n3476), .D(n3390), .Q(
        \inq_ary[15][60] ) );
  LATCHX1_RVT \dout_reg[60]  ( .CLK(n3492), .D(N321), .Q(dout[60]) );
  LATCHX1_RVT \inq_ary_reg[0][59]  ( .CLK(n3491), .D(n1524), .Q(
        \inq_ary[0][59] ) );
  LATCHX1_RVT \inq_ary_reg[1][59]  ( .CLK(n3490), .D(n1524), .Q(
        \inq_ary[1][59] ) );
  LATCHX1_RVT \inq_ary_reg[2][59]  ( .CLK(n3489), .D(n1524), .Q(
        \inq_ary[2][59] ) );
  LATCHX1_RVT \inq_ary_reg[3][59]  ( .CLK(n3488), .D(n1524), .Q(
        \inq_ary[3][59] ) );
  LATCHX1_RVT \inq_ary_reg[4][59]  ( .CLK(n3487), .D(n1524), .Q(
        \inq_ary[4][59] ) );
  LATCHX1_RVT \inq_ary_reg[5][59]  ( .CLK(n3486), .D(n1524), .Q(
        \inq_ary[5][59] ) );
  LATCHX1_RVT \inq_ary_reg[6][59]  ( .CLK(n3485), .D(n1524), .Q(
        \inq_ary[6][59] ) );
  LATCHX1_RVT \inq_ary_reg[7][59]  ( .CLK(n3484), .D(n1524), .Q(
        \inq_ary[7][59] ) );
  LATCHX1_RVT \inq_ary_reg[8][59]  ( .CLK(n3483), .D(n1524), .Q(
        \inq_ary[8][59] ) );
  LATCHX1_RVT \inq_ary_reg[9][59]  ( .CLK(n3482), .D(n1524), .Q(
        \inq_ary[9][59] ) );
  LATCHX1_RVT \inq_ary_reg[10][59]  ( .CLK(n3481), .D(n1524), .Q(
        \inq_ary[10][59] ) );
  LATCHX1_RVT \inq_ary_reg[11][59]  ( .CLK(n3480), .D(n1524), .Q(
        \inq_ary[11][59] ) );
  LATCHX1_RVT \inq_ary_reg[12][59]  ( .CLK(n3479), .D(n1524), .Q(
        \inq_ary[12][59] ) );
  LATCHX1_RVT \inq_ary_reg[13][59]  ( .CLK(n3478), .D(n1524), .Q(
        \inq_ary[13][59] ) );
  LATCHX1_RVT \inq_ary_reg[14][59]  ( .CLK(n3477), .D(n1524), .Q(
        \inq_ary[14][59] ) );
  LATCHX1_RVT \inq_ary_reg[15][59]  ( .CLK(n3476), .D(n1524), .Q(
        \inq_ary[15][59] ) );
  LATCHX1_RVT \dout_reg[59]  ( .CLK(n3492), .D(N320), .Q(dout[59]) );
  LATCHX1_RVT \inq_ary_reg[0][58]  ( .CLK(n3491), .D(n1562), .Q(
        \inq_ary[0][58] ) );
  LATCHX1_RVT \inq_ary_reg[1][58]  ( .CLK(n3490), .D(n1562), .Q(
        \inq_ary[1][58] ) );
  LATCHX1_RVT \inq_ary_reg[2][58]  ( .CLK(n3489), .D(n1562), .Q(
        \inq_ary[2][58] ) );
  LATCHX1_RVT \inq_ary_reg[3][58]  ( .CLK(n3488), .D(n1562), .Q(
        \inq_ary[3][58] ) );
  LATCHX1_RVT \inq_ary_reg[4][58]  ( .CLK(n3487), .D(n1562), .Q(
        \inq_ary[4][58] ) );
  LATCHX1_RVT \inq_ary_reg[5][58]  ( .CLK(n3486), .D(n1562), .Q(
        \inq_ary[5][58] ) );
  LATCHX1_RVT \inq_ary_reg[6][58]  ( .CLK(n3485), .D(n1562), .Q(
        \inq_ary[6][58] ) );
  LATCHX1_RVT \inq_ary_reg[7][58]  ( .CLK(n3484), .D(n1562), .Q(
        \inq_ary[7][58] ) );
  LATCHX1_RVT \inq_ary_reg[8][58]  ( .CLK(n3483), .D(n1562), .Q(
        \inq_ary[8][58] ) );
  LATCHX1_RVT \inq_ary_reg[9][58]  ( .CLK(n3482), .D(n1562), .Q(
        \inq_ary[9][58] ) );
  LATCHX1_RVT \inq_ary_reg[10][58]  ( .CLK(n3481), .D(n1562), .Q(
        \inq_ary[10][58] ) );
  LATCHX1_RVT \inq_ary_reg[11][58]  ( .CLK(n3480), .D(n1562), .Q(
        \inq_ary[11][58] ) );
  LATCHX1_RVT \inq_ary_reg[12][58]  ( .CLK(n3479), .D(n1562), .Q(
        \inq_ary[12][58] ) );
  LATCHX1_RVT \inq_ary_reg[13][58]  ( .CLK(n3478), .D(n1562), .Q(
        \inq_ary[13][58] ) );
  LATCHX1_RVT \inq_ary_reg[14][58]  ( .CLK(n3477), .D(n1562), .Q(
        \inq_ary[14][58] ) );
  LATCHX1_RVT \inq_ary_reg[15][58]  ( .CLK(n3476), .D(n1562), .Q(
        \inq_ary[15][58] ) );
  LATCHX1_RVT \dout_reg[58]  ( .CLK(n3492), .D(N319), .Q(dout[58]) );
  LATCHX1_RVT \inq_ary_reg[0][57]  ( .CLK(n3491), .D(n1574), .Q(
        \inq_ary[0][57] ) );
  LATCHX1_RVT \inq_ary_reg[1][57]  ( .CLK(n3490), .D(n1574), .Q(
        \inq_ary[1][57] ) );
  LATCHX1_RVT \inq_ary_reg[2][57]  ( .CLK(n3489), .D(n1574), .Q(
        \inq_ary[2][57] ) );
  LATCHX1_RVT \inq_ary_reg[3][57]  ( .CLK(n3488), .D(n1574), .Q(
        \inq_ary[3][57] ) );
  LATCHX1_RVT \inq_ary_reg[4][57]  ( .CLK(n3487), .D(n1574), .Q(
        \inq_ary[4][57] ) );
  LATCHX1_RVT \inq_ary_reg[5][57]  ( .CLK(n3486), .D(n1574), .Q(
        \inq_ary[5][57] ) );
  LATCHX1_RVT \inq_ary_reg[6][57]  ( .CLK(n3485), .D(n1574), .Q(
        \inq_ary[6][57] ) );
  LATCHX1_RVT \inq_ary_reg[7][57]  ( .CLK(n3484), .D(n1574), .Q(
        \inq_ary[7][57] ) );
  LATCHX1_RVT \inq_ary_reg[8][57]  ( .CLK(n3483), .D(n1574), .Q(
        \inq_ary[8][57] ) );
  LATCHX1_RVT \inq_ary_reg[9][57]  ( .CLK(n3482), .D(n1574), .Q(
        \inq_ary[9][57] ) );
  LATCHX1_RVT \inq_ary_reg[10][57]  ( .CLK(n3481), .D(n1574), .Q(
        \inq_ary[10][57] ) );
  LATCHX1_RVT \inq_ary_reg[11][57]  ( .CLK(n3480), .D(n1574), .Q(
        \inq_ary[11][57] ) );
  LATCHX1_RVT \inq_ary_reg[12][57]  ( .CLK(n3479), .D(n1574), .Q(
        \inq_ary[12][57] ) );
  LATCHX1_RVT \inq_ary_reg[13][57]  ( .CLK(n3478), .D(n1574), .Q(
        \inq_ary[13][57] ) );
  LATCHX1_RVT \inq_ary_reg[14][57]  ( .CLK(n3477), .D(n1574), .Q(
        \inq_ary[14][57] ) );
  LATCHX1_RVT \inq_ary_reg[15][57]  ( .CLK(n3476), .D(n1574), .Q(
        \inq_ary[15][57] ) );
  LATCHX1_RVT \dout_reg[57]  ( .CLK(n3492), .D(N318), .Q(dout[57]) );
  LATCHX1_RVT \inq_ary_reg[0][56]  ( .CLK(n3491), .D(n1586), .Q(
        \inq_ary[0][56] ) );
  LATCHX1_RVT \inq_ary_reg[1][56]  ( .CLK(n3490), .D(n1586), .Q(
        \inq_ary[1][56] ) );
  LATCHX1_RVT \inq_ary_reg[2][56]  ( .CLK(n3489), .D(n1586), .Q(
        \inq_ary[2][56] ) );
  LATCHX1_RVT \inq_ary_reg[3][56]  ( .CLK(n3488), .D(n1586), .Q(
        \inq_ary[3][56] ) );
  LATCHX1_RVT \inq_ary_reg[4][56]  ( .CLK(n3487), .D(n1586), .Q(
        \inq_ary[4][56] ) );
  LATCHX1_RVT \inq_ary_reg[5][56]  ( .CLK(n3486), .D(n1586), .Q(
        \inq_ary[5][56] ) );
  LATCHX1_RVT \inq_ary_reg[6][56]  ( .CLK(n3485), .D(n1586), .Q(
        \inq_ary[6][56] ) );
  LATCHX1_RVT \inq_ary_reg[7][56]  ( .CLK(n3484), .D(n1586), .Q(
        \inq_ary[7][56] ) );
  LATCHX1_RVT \inq_ary_reg[8][56]  ( .CLK(n3483), .D(n1586), .Q(
        \inq_ary[8][56] ) );
  LATCHX1_RVT \inq_ary_reg[9][56]  ( .CLK(n3482), .D(n1586), .Q(
        \inq_ary[9][56] ) );
  LATCHX1_RVT \inq_ary_reg[10][56]  ( .CLK(n3481), .D(n1586), .Q(
        \inq_ary[10][56] ) );
  LATCHX1_RVT \inq_ary_reg[11][56]  ( .CLK(n3480), .D(n1586), .Q(
        \inq_ary[11][56] ) );
  LATCHX1_RVT \inq_ary_reg[12][56]  ( .CLK(n3479), .D(n1586), .Q(
        \inq_ary[12][56] ) );
  LATCHX1_RVT \inq_ary_reg[13][56]  ( .CLK(n3478), .D(n1586), .Q(
        \inq_ary[13][56] ) );
  LATCHX1_RVT \inq_ary_reg[14][56]  ( .CLK(n3477), .D(n1586), .Q(
        \inq_ary[14][56] ) );
  LATCHX1_RVT \inq_ary_reg[15][56]  ( .CLK(n3476), .D(n1586), .Q(
        \inq_ary[15][56] ) );
  LATCHX1_RVT \dout_reg[56]  ( .CLK(n3492), .D(N317), .Q(dout[56]) );
  LATCHX1_RVT \inq_ary_reg[0][55]  ( .CLK(n3491), .D(n3388), .Q(
        \inq_ary[0][55] ) );
  LATCHX1_RVT \inq_ary_reg[1][55]  ( .CLK(n3490), .D(n3388), .Q(
        \inq_ary[1][55] ) );
  LATCHX1_RVT \inq_ary_reg[2][55]  ( .CLK(n3489), .D(n3388), .Q(
        \inq_ary[2][55] ) );
  LATCHX1_RVT \inq_ary_reg[3][55]  ( .CLK(n3488), .D(n3388), .Q(
        \inq_ary[3][55] ) );
  LATCHX1_RVT \inq_ary_reg[4][55]  ( .CLK(n3487), .D(n3388), .Q(
        \inq_ary[4][55] ) );
  LATCHX1_RVT \inq_ary_reg[5][55]  ( .CLK(n3486), .D(n3388), .Q(
        \inq_ary[5][55] ) );
  LATCHX1_RVT \inq_ary_reg[6][55]  ( .CLK(n3485), .D(n3388), .Q(
        \inq_ary[6][55] ) );
  LATCHX1_RVT \inq_ary_reg[7][55]  ( .CLK(n3484), .D(n3388), .Q(
        \inq_ary[7][55] ) );
  LATCHX1_RVT \inq_ary_reg[8][55]  ( .CLK(n3483), .D(n3388), .Q(
        \inq_ary[8][55] ) );
  LATCHX1_RVT \inq_ary_reg[9][55]  ( .CLK(n3482), .D(n3388), .Q(
        \inq_ary[9][55] ) );
  LATCHX1_RVT \inq_ary_reg[10][55]  ( .CLK(n3481), .D(n3388), .Q(
        \inq_ary[10][55] ) );
  LATCHX1_RVT \inq_ary_reg[11][55]  ( .CLK(n3480), .D(n3388), .Q(
        \inq_ary[11][55] ) );
  LATCHX1_RVT \inq_ary_reg[12][55]  ( .CLK(n3479), .D(n3388), .Q(
        \inq_ary[12][55] ) );
  LATCHX1_RVT \inq_ary_reg[13][55]  ( .CLK(n3478), .D(n3388), .Q(
        \inq_ary[13][55] ) );
  LATCHX1_RVT \inq_ary_reg[14][55]  ( .CLK(n3477), .D(n3388), .Q(
        \inq_ary[14][55] ) );
  LATCHX1_RVT \inq_ary_reg[15][55]  ( .CLK(n3476), .D(n3388), .Q(
        \inq_ary[15][55] ) );
  LATCHX1_RVT \dout_reg[55]  ( .CLK(n3492), .D(N316), .Q(dout[55]) );
  LATCHX1_RVT \inq_ary_reg[0][54]  ( .CLK(n3491), .D(n3386), .Q(
        \inq_ary[0][54] ) );
  LATCHX1_RVT \inq_ary_reg[1][54]  ( .CLK(n3490), .D(n3386), .Q(
        \inq_ary[1][54] ) );
  LATCHX1_RVT \inq_ary_reg[2][54]  ( .CLK(n3489), .D(n3386), .Q(
        \inq_ary[2][54] ) );
  LATCHX1_RVT \inq_ary_reg[3][54]  ( .CLK(n3488), .D(n3386), .Q(
        \inq_ary[3][54] ) );
  LATCHX1_RVT \inq_ary_reg[4][54]  ( .CLK(n3487), .D(n3386), .Q(
        \inq_ary[4][54] ) );
  LATCHX1_RVT \inq_ary_reg[5][54]  ( .CLK(n3486), .D(n3386), .Q(
        \inq_ary[5][54] ) );
  LATCHX1_RVT \inq_ary_reg[6][54]  ( .CLK(n3485), .D(n3386), .Q(
        \inq_ary[6][54] ) );
  LATCHX1_RVT \inq_ary_reg[7][54]  ( .CLK(n3484), .D(n3386), .Q(
        \inq_ary[7][54] ) );
  LATCHX1_RVT \inq_ary_reg[8][54]  ( .CLK(n3483), .D(n3386), .Q(
        \inq_ary[8][54] ) );
  LATCHX1_RVT \inq_ary_reg[9][54]  ( .CLK(n3482), .D(n3386), .Q(
        \inq_ary[9][54] ) );
  LATCHX1_RVT \inq_ary_reg[10][54]  ( .CLK(n3481), .D(n3386), .Q(
        \inq_ary[10][54] ) );
  LATCHX1_RVT \inq_ary_reg[11][54]  ( .CLK(n3480), .D(n3386), .Q(
        \inq_ary[11][54] ) );
  LATCHX1_RVT \inq_ary_reg[12][54]  ( .CLK(n3479), .D(n3386), .Q(
        \inq_ary[12][54] ) );
  LATCHX1_RVT \inq_ary_reg[13][54]  ( .CLK(n3478), .D(n3386), .Q(
        \inq_ary[13][54] ) );
  LATCHX1_RVT \inq_ary_reg[14][54]  ( .CLK(n3477), .D(n3386), .Q(
        \inq_ary[14][54] ) );
  LATCHX1_RVT \inq_ary_reg[15][54]  ( .CLK(n3476), .D(n3386), .Q(
        \inq_ary[15][54] ) );
  LATCHX1_RVT \dout_reg[54]  ( .CLK(n3492), .D(N315), .Q(dout[54]) );
  LATCHX1_RVT \inq_ary_reg[0][53]  ( .CLK(n3491), .D(n3384), .Q(
        \inq_ary[0][53] ) );
  LATCHX1_RVT \inq_ary_reg[1][53]  ( .CLK(n3490), .D(n3384), .Q(
        \inq_ary[1][53] ) );
  LATCHX1_RVT \inq_ary_reg[2][53]  ( .CLK(n3489), .D(n3384), .Q(
        \inq_ary[2][53] ) );
  LATCHX1_RVT \inq_ary_reg[3][53]  ( .CLK(n3488), .D(n3384), .Q(
        \inq_ary[3][53] ) );
  LATCHX1_RVT \inq_ary_reg[4][53]  ( .CLK(n3487), .D(n3384), .Q(
        \inq_ary[4][53] ) );
  LATCHX1_RVT \inq_ary_reg[5][53]  ( .CLK(n3486), .D(n3384), .Q(
        \inq_ary[5][53] ) );
  LATCHX1_RVT \inq_ary_reg[6][53]  ( .CLK(n3485), .D(n3384), .Q(
        \inq_ary[6][53] ) );
  LATCHX1_RVT \inq_ary_reg[7][53]  ( .CLK(n3484), .D(n3384), .Q(
        \inq_ary[7][53] ) );
  LATCHX1_RVT \inq_ary_reg[8][53]  ( .CLK(n3483), .D(n3384), .Q(
        \inq_ary[8][53] ) );
  LATCHX1_RVT \inq_ary_reg[9][53]  ( .CLK(n3482), .D(n3384), .Q(
        \inq_ary[9][53] ) );
  LATCHX1_RVT \inq_ary_reg[10][53]  ( .CLK(n3481), .D(n3384), .Q(
        \inq_ary[10][53] ) );
  LATCHX1_RVT \inq_ary_reg[11][53]  ( .CLK(n3480), .D(n3384), .Q(
        \inq_ary[11][53] ) );
  LATCHX1_RVT \inq_ary_reg[12][53]  ( .CLK(n3479), .D(n3384), .Q(
        \inq_ary[12][53] ) );
  LATCHX1_RVT \inq_ary_reg[13][53]  ( .CLK(n3478), .D(n3384), .Q(
        \inq_ary[13][53] ) );
  LATCHX1_RVT \inq_ary_reg[14][53]  ( .CLK(n3477), .D(n3384), .Q(
        \inq_ary[14][53] ) );
  LATCHX1_RVT \inq_ary_reg[15][53]  ( .CLK(n3476), .D(n3384), .Q(
        \inq_ary[15][53] ) );
  LATCHX1_RVT \dout_reg[53]  ( .CLK(n3492), .D(N314), .Q(dout[53]) );
  LATCHX1_RVT \inq_ary_reg[0][52]  ( .CLK(n3491), .D(n1599), .Q(
        \inq_ary[0][52] ) );
  LATCHX1_RVT \inq_ary_reg[1][52]  ( .CLK(n3490), .D(n1599), .Q(
        \inq_ary[1][52] ) );
  LATCHX1_RVT \inq_ary_reg[2][52]  ( .CLK(n3489), .D(n1599), .Q(
        \inq_ary[2][52] ) );
  LATCHX1_RVT \inq_ary_reg[3][52]  ( .CLK(n3488), .D(n1599), .Q(
        \inq_ary[3][52] ) );
  LATCHX1_RVT \inq_ary_reg[4][52]  ( .CLK(n3487), .D(n1599), .Q(
        \inq_ary[4][52] ) );
  LATCHX1_RVT \inq_ary_reg[5][52]  ( .CLK(n3486), .D(n1599), .Q(
        \inq_ary[5][52] ) );
  LATCHX1_RVT \inq_ary_reg[6][52]  ( .CLK(n3485), .D(n1599), .Q(
        \inq_ary[6][52] ) );
  LATCHX1_RVT \inq_ary_reg[7][52]  ( .CLK(n3484), .D(n1599), .Q(
        \inq_ary[7][52] ) );
  LATCHX1_RVT \inq_ary_reg[8][52]  ( .CLK(n3483), .D(n1599), .Q(
        \inq_ary[8][52] ) );
  LATCHX1_RVT \inq_ary_reg[9][52]  ( .CLK(n3482), .D(n1599), .Q(
        \inq_ary[9][52] ) );
  LATCHX1_RVT \inq_ary_reg[10][52]  ( .CLK(n3481), .D(n1599), .Q(
        \inq_ary[10][52] ) );
  LATCHX1_RVT \inq_ary_reg[11][52]  ( .CLK(n3480), .D(n1599), .Q(
        \inq_ary[11][52] ) );
  LATCHX1_RVT \inq_ary_reg[12][52]  ( .CLK(n3479), .D(n1599), .Q(
        \inq_ary[12][52] ) );
  LATCHX1_RVT \inq_ary_reg[13][52]  ( .CLK(n3478), .D(n1599), .Q(
        \inq_ary[13][52] ) );
  LATCHX1_RVT \inq_ary_reg[14][52]  ( .CLK(n3477), .D(n1599), .Q(
        \inq_ary[14][52] ) );
  LATCHX1_RVT \inq_ary_reg[15][52]  ( .CLK(n3476), .D(n1599), .Q(
        \inq_ary[15][52] ) );
  LATCHX1_RVT \dout_reg[52]  ( .CLK(n3492), .D(N313), .Q(dout[52]) );
  LATCHX1_RVT \inq_ary_reg[0][51]  ( .CLK(n3491), .D(n3389), .Q(
        \inq_ary[0][51] ) );
  LATCHX1_RVT \inq_ary_reg[1][51]  ( .CLK(n3490), .D(n3389), .Q(
        \inq_ary[1][51] ) );
  LATCHX1_RVT \inq_ary_reg[2][51]  ( .CLK(n3489), .D(n3389), .Q(
        \inq_ary[2][51] ) );
  LATCHX1_RVT \inq_ary_reg[3][51]  ( .CLK(n3488), .D(n3389), .Q(
        \inq_ary[3][51] ) );
  LATCHX1_RVT \inq_ary_reg[4][51]  ( .CLK(n3487), .D(n3389), .Q(
        \inq_ary[4][51] ) );
  LATCHX1_RVT \inq_ary_reg[5][51]  ( .CLK(n3486), .D(n3389), .Q(
        \inq_ary[5][51] ) );
  LATCHX1_RVT \inq_ary_reg[6][51]  ( .CLK(n3485), .D(n3389), .Q(
        \inq_ary[6][51] ) );
  LATCHX1_RVT \inq_ary_reg[7][51]  ( .CLK(n3484), .D(n3389), .Q(
        \inq_ary[7][51] ) );
  LATCHX1_RVT \inq_ary_reg[8][51]  ( .CLK(n3483), .D(n3389), .Q(
        \inq_ary[8][51] ) );
  LATCHX1_RVT \inq_ary_reg[9][51]  ( .CLK(n3482), .D(n3389), .Q(
        \inq_ary[9][51] ) );
  LATCHX1_RVT \inq_ary_reg[10][51]  ( .CLK(n3481), .D(n3389), .Q(
        \inq_ary[10][51] ) );
  LATCHX1_RVT \inq_ary_reg[11][51]  ( .CLK(n3480), .D(n3389), .Q(
        \inq_ary[11][51] ) );
  LATCHX1_RVT \inq_ary_reg[12][51]  ( .CLK(n3479), .D(n3389), .Q(
        \inq_ary[12][51] ) );
  LATCHX1_RVT \inq_ary_reg[13][51]  ( .CLK(n3478), .D(n3389), .Q(
        \inq_ary[13][51] ) );
  LATCHX1_RVT \inq_ary_reg[14][51]  ( .CLK(n3477), .D(n3389), .Q(
        \inq_ary[14][51] ) );
  LATCHX1_RVT \inq_ary_reg[15][51]  ( .CLK(n3476), .D(n3389), .Q(
        \inq_ary[15][51] ) );
  LATCHX1_RVT \dout_reg[51]  ( .CLK(n3492), .D(N312), .Q(dout[51]) );
  LATCHX1_RVT \inq_ary_reg[0][50]  ( .CLK(n3491), .D(n3387), .Q(
        \inq_ary[0][50] ) );
  LATCHX1_RVT \inq_ary_reg[1][50]  ( .CLK(n3490), .D(n3387), .Q(
        \inq_ary[1][50] ) );
  LATCHX1_RVT \inq_ary_reg[2][50]  ( .CLK(n3489), .D(n3387), .Q(
        \inq_ary[2][50] ) );
  LATCHX1_RVT \inq_ary_reg[3][50]  ( .CLK(n3488), .D(n3387), .Q(
        \inq_ary[3][50] ) );
  LATCHX1_RVT \inq_ary_reg[4][50]  ( .CLK(n3487), .D(n3387), .Q(
        \inq_ary[4][50] ) );
  LATCHX1_RVT \inq_ary_reg[5][50]  ( .CLK(n3486), .D(n3387), .Q(
        \inq_ary[5][50] ) );
  LATCHX1_RVT \inq_ary_reg[6][50]  ( .CLK(n3485), .D(n3387), .Q(
        \inq_ary[6][50] ) );
  LATCHX1_RVT \inq_ary_reg[7][50]  ( .CLK(n3484), .D(n3387), .Q(
        \inq_ary[7][50] ) );
  LATCHX1_RVT \inq_ary_reg[8][50]  ( .CLK(n3483), .D(n3387), .Q(
        \inq_ary[8][50] ) );
  LATCHX1_RVT \inq_ary_reg[9][50]  ( .CLK(n3482), .D(n3387), .Q(
        \inq_ary[9][50] ) );
  LATCHX1_RVT \inq_ary_reg[10][50]  ( .CLK(n3481), .D(n3387), .Q(
        \inq_ary[10][50] ) );
  LATCHX1_RVT \inq_ary_reg[11][50]  ( .CLK(n3480), .D(n3387), .Q(
        \inq_ary[11][50] ) );
  LATCHX1_RVT \inq_ary_reg[12][50]  ( .CLK(n3479), .D(n3387), .Q(
        \inq_ary[12][50] ) );
  LATCHX1_RVT \inq_ary_reg[13][50]  ( .CLK(n3478), .D(n3387), .Q(
        \inq_ary[13][50] ) );
  LATCHX1_RVT \inq_ary_reg[14][50]  ( .CLK(n3477), .D(n3387), .Q(
        \inq_ary[14][50] ) );
  LATCHX1_RVT \inq_ary_reg[15][50]  ( .CLK(n3476), .D(n3387), .Q(
        \inq_ary[15][50] ) );
  LATCHX1_RVT \dout_reg[50]  ( .CLK(n3492), .D(N311), .Q(dout[50]) );
  LATCHX1_RVT \inq_ary_reg[0][49]  ( .CLK(n3491), .D(n3385), .Q(
        \inq_ary[0][49] ) );
  LATCHX1_RVT \inq_ary_reg[1][49]  ( .CLK(n3490), .D(n3385), .Q(
        \inq_ary[1][49] ) );
  LATCHX1_RVT \inq_ary_reg[2][49]  ( .CLK(n3489), .D(n3385), .Q(
        \inq_ary[2][49] ) );
  LATCHX1_RVT \inq_ary_reg[3][49]  ( .CLK(n3488), .D(n3385), .Q(
        \inq_ary[3][49] ) );
  LATCHX1_RVT \inq_ary_reg[4][49]  ( .CLK(n3487), .D(n3385), .Q(
        \inq_ary[4][49] ) );
  LATCHX1_RVT \inq_ary_reg[5][49]  ( .CLK(n3486), .D(n3385), .Q(
        \inq_ary[5][49] ) );
  LATCHX1_RVT \inq_ary_reg[6][49]  ( .CLK(n3485), .D(n3385), .Q(
        \inq_ary[6][49] ) );
  LATCHX1_RVT \inq_ary_reg[7][49]  ( .CLK(n3484), .D(n3385), .Q(
        \inq_ary[7][49] ) );
  LATCHX1_RVT \inq_ary_reg[8][49]  ( .CLK(n3483), .D(n3385), .Q(
        \inq_ary[8][49] ) );
  LATCHX1_RVT \inq_ary_reg[9][49]  ( .CLK(n3482), .D(n3385), .Q(
        \inq_ary[9][49] ) );
  LATCHX1_RVT \inq_ary_reg[10][49]  ( .CLK(n3481), .D(n3385), .Q(
        \inq_ary[10][49] ) );
  LATCHX1_RVT \inq_ary_reg[11][49]  ( .CLK(n3480), .D(n3385), .Q(
        \inq_ary[11][49] ) );
  LATCHX1_RVT \inq_ary_reg[12][49]  ( .CLK(n3479), .D(n3385), .Q(
        \inq_ary[12][49] ) );
  LATCHX1_RVT \inq_ary_reg[13][49]  ( .CLK(n3478), .D(n3385), .Q(
        \inq_ary[13][49] ) );
  LATCHX1_RVT \inq_ary_reg[14][49]  ( .CLK(n3477), .D(n3385), .Q(
        \inq_ary[14][49] ) );
  LATCHX1_RVT \inq_ary_reg[15][49]  ( .CLK(n3476), .D(n3385), .Q(
        \inq_ary[15][49] ) );
  LATCHX1_RVT \dout_reg[49]  ( .CLK(n3492), .D(N310), .Q(dout[49]) );
  LATCHX1_RVT \inq_ary_reg[0][48]  ( .CLK(n3491), .D(n3383), .Q(
        \inq_ary[0][48] ) );
  LATCHX1_RVT \inq_ary_reg[1][48]  ( .CLK(n3490), .D(n3383), .Q(
        \inq_ary[1][48] ) );
  LATCHX1_RVT \inq_ary_reg[2][48]  ( .CLK(n3489), .D(n3383), .Q(
        \inq_ary[2][48] ) );
  LATCHX1_RVT \inq_ary_reg[3][48]  ( .CLK(n3488), .D(n3383), .Q(
        \inq_ary[3][48] ) );
  LATCHX1_RVT \inq_ary_reg[4][48]  ( .CLK(n3487), .D(n3383), .Q(
        \inq_ary[4][48] ) );
  LATCHX1_RVT \inq_ary_reg[5][48]  ( .CLK(n3486), .D(n3383), .Q(
        \inq_ary[5][48] ) );
  LATCHX1_RVT \inq_ary_reg[6][48]  ( .CLK(n3485), .D(n3383), .Q(
        \inq_ary[6][48] ) );
  LATCHX1_RVT \inq_ary_reg[7][48]  ( .CLK(n3484), .D(n3383), .Q(
        \inq_ary[7][48] ) );
  LATCHX1_RVT \inq_ary_reg[8][48]  ( .CLK(n3483), .D(n3383), .Q(
        \inq_ary[8][48] ) );
  LATCHX1_RVT \inq_ary_reg[9][48]  ( .CLK(n3482), .D(n3383), .Q(
        \inq_ary[9][48] ) );
  LATCHX1_RVT \inq_ary_reg[10][48]  ( .CLK(n3481), .D(n3383), .Q(
        \inq_ary[10][48] ) );
  LATCHX1_RVT \inq_ary_reg[11][48]  ( .CLK(n3480), .D(n3383), .Q(
        \inq_ary[11][48] ) );
  LATCHX1_RVT \inq_ary_reg[12][48]  ( .CLK(n3479), .D(n3383), .Q(
        \inq_ary[12][48] ) );
  LATCHX1_RVT \inq_ary_reg[13][48]  ( .CLK(n3478), .D(n3383), .Q(
        \inq_ary[13][48] ) );
  LATCHX1_RVT \inq_ary_reg[14][48]  ( .CLK(n3477), .D(n3383), .Q(
        \inq_ary[14][48] ) );
  LATCHX1_RVT \inq_ary_reg[15][48]  ( .CLK(n3476), .D(n3383), .Q(
        \inq_ary[15][48] ) );
  LATCHX1_RVT \dout_reg[48]  ( .CLK(n3492), .D(N309), .Q(dout[48]) );
  LATCHX1_RVT \inq_ary_reg[0][47]  ( .CLK(n3491), .D(n3381), .Q(
        \inq_ary[0][47] ) );
  LATCHX1_RVT \inq_ary_reg[1][47]  ( .CLK(n3490), .D(n3381), .Q(
        \inq_ary[1][47] ) );
  LATCHX1_RVT \inq_ary_reg[2][47]  ( .CLK(n3489), .D(n3381), .Q(
        \inq_ary[2][47] ) );
  LATCHX1_RVT \inq_ary_reg[3][47]  ( .CLK(n3488), .D(n3381), .Q(
        \inq_ary[3][47] ) );
  LATCHX1_RVT \inq_ary_reg[4][47]  ( .CLK(n3487), .D(n3381), .Q(
        \inq_ary[4][47] ) );
  LATCHX1_RVT \inq_ary_reg[5][47]  ( .CLK(n3486), .D(n3381), .Q(
        \inq_ary[5][47] ) );
  LATCHX1_RVT \inq_ary_reg[6][47]  ( .CLK(n3485), .D(n3381), .Q(
        \inq_ary[6][47] ) );
  LATCHX1_RVT \inq_ary_reg[7][47]  ( .CLK(n3484), .D(n3381), .Q(
        \inq_ary[7][47] ) );
  LATCHX1_RVT \inq_ary_reg[8][47]  ( .CLK(n3483), .D(n3381), .Q(
        \inq_ary[8][47] ) );
  LATCHX1_RVT \inq_ary_reg[9][47]  ( .CLK(n3482), .D(n3381), .Q(
        \inq_ary[9][47] ) );
  LATCHX1_RVT \inq_ary_reg[10][47]  ( .CLK(n3481), .D(n3381), .Q(
        \inq_ary[10][47] ) );
  LATCHX1_RVT \inq_ary_reg[11][47]  ( .CLK(n3480), .D(n3381), .Q(
        \inq_ary[11][47] ) );
  LATCHX1_RVT \inq_ary_reg[12][47]  ( .CLK(n3479), .D(n3381), .Q(
        \inq_ary[12][47] ) );
  LATCHX1_RVT \inq_ary_reg[13][47]  ( .CLK(n3478), .D(n3381), .Q(
        \inq_ary[13][47] ) );
  LATCHX1_RVT \inq_ary_reg[14][47]  ( .CLK(n3477), .D(n3381), .Q(
        \inq_ary[14][47] ) );
  LATCHX1_RVT \inq_ary_reg[15][47]  ( .CLK(n3476), .D(n3381), .Q(
        \inq_ary[15][47] ) );
  LATCHX1_RVT \dout_reg[47]  ( .CLK(n3492), .D(N308), .Q(dout[47]) );
  LATCHX1_RVT \inq_ary_reg[0][46]  ( .CLK(n3491), .D(n3379), .Q(
        \inq_ary[0][46] ) );
  LATCHX1_RVT \inq_ary_reg[1][46]  ( .CLK(n3490), .D(n3379), .Q(
        \inq_ary[1][46] ) );
  LATCHX1_RVT \inq_ary_reg[2][46]  ( .CLK(n3489), .D(n3379), .Q(
        \inq_ary[2][46] ) );
  LATCHX1_RVT \inq_ary_reg[3][46]  ( .CLK(n3488), .D(n3379), .Q(
        \inq_ary[3][46] ) );
  LATCHX1_RVT \inq_ary_reg[4][46]  ( .CLK(n3487), .D(n3379), .Q(
        \inq_ary[4][46] ) );
  LATCHX1_RVT \inq_ary_reg[5][46]  ( .CLK(n3486), .D(n3379), .Q(
        \inq_ary[5][46] ) );
  LATCHX1_RVT \inq_ary_reg[6][46]  ( .CLK(n3485), .D(n3379), .Q(
        \inq_ary[6][46] ) );
  LATCHX1_RVT \inq_ary_reg[7][46]  ( .CLK(n3484), .D(n3379), .Q(
        \inq_ary[7][46] ) );
  LATCHX1_RVT \inq_ary_reg[8][46]  ( .CLK(n3483), .D(n3379), .Q(
        \inq_ary[8][46] ) );
  LATCHX1_RVT \inq_ary_reg[9][46]  ( .CLK(n3482), .D(n3379), .Q(
        \inq_ary[9][46] ) );
  LATCHX1_RVT \inq_ary_reg[10][46]  ( .CLK(n3481), .D(n3379), .Q(
        \inq_ary[10][46] ) );
  LATCHX1_RVT \inq_ary_reg[11][46]  ( .CLK(n3480), .D(n3379), .Q(
        \inq_ary[11][46] ) );
  LATCHX1_RVT \inq_ary_reg[12][46]  ( .CLK(n3479), .D(n3379), .Q(
        \inq_ary[12][46] ) );
  LATCHX1_RVT \inq_ary_reg[13][46]  ( .CLK(n3478), .D(n3379), .Q(
        \inq_ary[13][46] ) );
  LATCHX1_RVT \inq_ary_reg[14][46]  ( .CLK(n3477), .D(n3379), .Q(
        \inq_ary[14][46] ) );
  LATCHX1_RVT \inq_ary_reg[15][46]  ( .CLK(n3476), .D(n3379), .Q(
        \inq_ary[15][46] ) );
  LATCHX1_RVT \dout_reg[46]  ( .CLK(n3492), .D(N307), .Q(dout[46]) );
  LATCHX1_RVT \inq_ary_reg[0][45]  ( .CLK(n3491), .D(n3377), .Q(
        \inq_ary[0][45] ) );
  LATCHX1_RVT \inq_ary_reg[1][45]  ( .CLK(n3490), .D(n3377), .Q(
        \inq_ary[1][45] ) );
  LATCHX1_RVT \inq_ary_reg[2][45]  ( .CLK(n3489), .D(n3377), .Q(
        \inq_ary[2][45] ) );
  LATCHX1_RVT \inq_ary_reg[3][45]  ( .CLK(n3488), .D(n3377), .Q(
        \inq_ary[3][45] ) );
  LATCHX1_RVT \inq_ary_reg[4][45]  ( .CLK(n3487), .D(n3377), .Q(
        \inq_ary[4][45] ) );
  LATCHX1_RVT \inq_ary_reg[5][45]  ( .CLK(n3486), .D(n3377), .Q(
        \inq_ary[5][45] ) );
  LATCHX1_RVT \inq_ary_reg[6][45]  ( .CLK(n3485), .D(n3377), .Q(
        \inq_ary[6][45] ) );
  LATCHX1_RVT \inq_ary_reg[7][45]  ( .CLK(n3484), .D(n3377), .Q(
        \inq_ary[7][45] ) );
  LATCHX1_RVT \inq_ary_reg[8][45]  ( .CLK(n3483), .D(n3377), .Q(
        \inq_ary[8][45] ) );
  LATCHX1_RVT \inq_ary_reg[9][45]  ( .CLK(n3482), .D(n3377), .Q(
        \inq_ary[9][45] ) );
  LATCHX1_RVT \inq_ary_reg[10][45]  ( .CLK(n3481), .D(n3377), .Q(
        \inq_ary[10][45] ) );
  LATCHX1_RVT \inq_ary_reg[11][45]  ( .CLK(n3480), .D(n3377), .Q(
        \inq_ary[11][45] ) );
  LATCHX1_RVT \inq_ary_reg[12][45]  ( .CLK(n3479), .D(n3377), .Q(
        \inq_ary[12][45] ) );
  LATCHX1_RVT \inq_ary_reg[13][45]  ( .CLK(n3478), .D(n3377), .Q(
        \inq_ary[13][45] ) );
  LATCHX1_RVT \inq_ary_reg[14][45]  ( .CLK(n3477), .D(n3377), .Q(
        \inq_ary[14][45] ) );
  LATCHX1_RVT \inq_ary_reg[15][45]  ( .CLK(n3476), .D(n3377), .Q(
        \inq_ary[15][45] ) );
  LATCHX1_RVT \dout_reg[45]  ( .CLK(n3492), .D(N306), .Q(dout[45]) );
  LATCHX1_RVT \inq_ary_reg[0][44]  ( .CLK(n3491), .D(n3375), .Q(
        \inq_ary[0][44] ) );
  LATCHX1_RVT \inq_ary_reg[1][44]  ( .CLK(n3490), .D(n3375), .Q(
        \inq_ary[1][44] ) );
  LATCHX1_RVT \inq_ary_reg[2][44]  ( .CLK(n3489), .D(n3375), .Q(
        \inq_ary[2][44] ) );
  LATCHX1_RVT \inq_ary_reg[3][44]  ( .CLK(n3488), .D(n3375), .Q(
        \inq_ary[3][44] ) );
  LATCHX1_RVT \inq_ary_reg[4][44]  ( .CLK(n3487), .D(n3375), .Q(
        \inq_ary[4][44] ) );
  LATCHX1_RVT \inq_ary_reg[5][44]  ( .CLK(n3486), .D(n3375), .Q(
        \inq_ary[5][44] ) );
  LATCHX1_RVT \inq_ary_reg[6][44]  ( .CLK(n3485), .D(n3375), .Q(
        \inq_ary[6][44] ) );
  LATCHX1_RVT \inq_ary_reg[7][44]  ( .CLK(n3484), .D(n3375), .Q(
        \inq_ary[7][44] ) );
  LATCHX1_RVT \inq_ary_reg[8][44]  ( .CLK(n3483), .D(n3375), .Q(
        \inq_ary[8][44] ) );
  LATCHX1_RVT \inq_ary_reg[9][44]  ( .CLK(n3482), .D(n3375), .Q(
        \inq_ary[9][44] ) );
  LATCHX1_RVT \inq_ary_reg[10][44]  ( .CLK(n3481), .D(n3375), .Q(
        \inq_ary[10][44] ) );
  LATCHX1_RVT \inq_ary_reg[11][44]  ( .CLK(n3480), .D(n3375), .Q(
        \inq_ary[11][44] ) );
  LATCHX1_RVT \inq_ary_reg[12][44]  ( .CLK(n3479), .D(n3375), .Q(
        \inq_ary[12][44] ) );
  LATCHX1_RVT \inq_ary_reg[13][44]  ( .CLK(n3478), .D(n3375), .Q(
        \inq_ary[13][44] ) );
  LATCHX1_RVT \inq_ary_reg[14][44]  ( .CLK(n3477), .D(n3375), .Q(
        \inq_ary[14][44] ) );
  LATCHX1_RVT \inq_ary_reg[15][44]  ( .CLK(n3476), .D(n3375), .Q(
        \inq_ary[15][44] ) );
  LATCHX1_RVT \dout_reg[44]  ( .CLK(n3492), .D(N305), .Q(dout[44]) );
  LATCHX1_RVT \inq_ary_reg[0][43]  ( .CLK(n3491), .D(n3382), .Q(
        \inq_ary[0][43] ) );
  LATCHX1_RVT \inq_ary_reg[1][43]  ( .CLK(n3490), .D(n3382), .Q(
        \inq_ary[1][43] ) );
  LATCHX1_RVT \inq_ary_reg[2][43]  ( .CLK(n3489), .D(n3382), .Q(
        \inq_ary[2][43] ) );
  LATCHX1_RVT \inq_ary_reg[3][43]  ( .CLK(n3488), .D(n3382), .Q(
        \inq_ary[3][43] ) );
  LATCHX1_RVT \inq_ary_reg[4][43]  ( .CLK(n3487), .D(n3382), .Q(
        \inq_ary[4][43] ) );
  LATCHX1_RVT \inq_ary_reg[5][43]  ( .CLK(n3486), .D(n3382), .Q(
        \inq_ary[5][43] ) );
  LATCHX1_RVT \inq_ary_reg[6][43]  ( .CLK(n3485), .D(n3382), .Q(
        \inq_ary[6][43] ) );
  LATCHX1_RVT \inq_ary_reg[7][43]  ( .CLK(n3484), .D(n3382), .Q(
        \inq_ary[7][43] ) );
  LATCHX1_RVT \inq_ary_reg[8][43]  ( .CLK(n3483), .D(n3382), .Q(
        \inq_ary[8][43] ) );
  LATCHX1_RVT \inq_ary_reg[9][43]  ( .CLK(n3482), .D(n3382), .Q(
        \inq_ary[9][43] ) );
  LATCHX1_RVT \inq_ary_reg[10][43]  ( .CLK(n3481), .D(n3382), .Q(
        \inq_ary[10][43] ) );
  LATCHX1_RVT \inq_ary_reg[11][43]  ( .CLK(n3480), .D(n3382), .Q(
        \inq_ary[11][43] ) );
  LATCHX1_RVT \inq_ary_reg[12][43]  ( .CLK(n3479), .D(n3382), .Q(
        \inq_ary[12][43] ) );
  LATCHX1_RVT \inq_ary_reg[13][43]  ( .CLK(n3478), .D(n3382), .Q(
        \inq_ary[13][43] ) );
  LATCHX1_RVT \inq_ary_reg[14][43]  ( .CLK(n3477), .D(n3382), .Q(
        \inq_ary[14][43] ) );
  LATCHX1_RVT \inq_ary_reg[15][43]  ( .CLK(n3476), .D(n3382), .Q(
        \inq_ary[15][43] ) );
  LATCHX1_RVT \dout_reg[43]  ( .CLK(n3492), .D(N304), .Q(dout[43]) );
  LATCHX1_RVT \inq_ary_reg[0][42]  ( .CLK(n3491), .D(n3380), .Q(
        \inq_ary[0][42] ) );
  LATCHX1_RVT \inq_ary_reg[1][42]  ( .CLK(n3490), .D(n3380), .Q(
        \inq_ary[1][42] ) );
  LATCHX1_RVT \inq_ary_reg[2][42]  ( .CLK(n3489), .D(n3380), .Q(
        \inq_ary[2][42] ) );
  LATCHX1_RVT \inq_ary_reg[3][42]  ( .CLK(n3488), .D(n3380), .Q(
        \inq_ary[3][42] ) );
  LATCHX1_RVT \inq_ary_reg[4][42]  ( .CLK(n3487), .D(n3380), .Q(
        \inq_ary[4][42] ) );
  LATCHX1_RVT \inq_ary_reg[5][42]  ( .CLK(n3486), .D(n3380), .Q(
        \inq_ary[5][42] ) );
  LATCHX1_RVT \inq_ary_reg[6][42]  ( .CLK(n3485), .D(n3380), .Q(
        \inq_ary[6][42] ) );
  LATCHX1_RVT \inq_ary_reg[7][42]  ( .CLK(n3484), .D(n3380), .Q(
        \inq_ary[7][42] ) );
  LATCHX1_RVT \inq_ary_reg[8][42]  ( .CLK(n3483), .D(n3380), .Q(
        \inq_ary[8][42] ) );
  LATCHX1_RVT \inq_ary_reg[9][42]  ( .CLK(n3482), .D(n3380), .Q(
        \inq_ary[9][42] ) );
  LATCHX1_RVT \inq_ary_reg[10][42]  ( .CLK(n3481), .D(n3380), .Q(
        \inq_ary[10][42] ) );
  LATCHX1_RVT \inq_ary_reg[11][42]  ( .CLK(n3480), .D(n3380), .Q(
        \inq_ary[11][42] ) );
  LATCHX1_RVT \inq_ary_reg[12][42]  ( .CLK(n3479), .D(n3380), .Q(
        \inq_ary[12][42] ) );
  LATCHX1_RVT \inq_ary_reg[13][42]  ( .CLK(n3478), .D(n3380), .Q(
        \inq_ary[13][42] ) );
  LATCHX1_RVT \inq_ary_reg[14][42]  ( .CLK(n3477), .D(n3380), .Q(
        \inq_ary[14][42] ) );
  LATCHX1_RVT \inq_ary_reg[15][42]  ( .CLK(n3476), .D(n3380), .Q(
        \inq_ary[15][42] ) );
  LATCHX1_RVT \dout_reg[42]  ( .CLK(n3492), .D(N303), .Q(dout[42]) );
  LATCHX1_RVT \inq_ary_reg[0][41]  ( .CLK(n3491), .D(n3378), .Q(
        \inq_ary[0][41] ) );
  LATCHX1_RVT \inq_ary_reg[1][41]  ( .CLK(n3490), .D(n3378), .Q(
        \inq_ary[1][41] ) );
  LATCHX1_RVT \inq_ary_reg[2][41]  ( .CLK(n3489), .D(n3378), .Q(
        \inq_ary[2][41] ) );
  LATCHX1_RVT \inq_ary_reg[3][41]  ( .CLK(n3488), .D(n3378), .Q(
        \inq_ary[3][41] ) );
  LATCHX1_RVT \inq_ary_reg[4][41]  ( .CLK(n3487), .D(n3378), .Q(
        \inq_ary[4][41] ) );
  LATCHX1_RVT \inq_ary_reg[5][41]  ( .CLK(n3486), .D(n3378), .Q(
        \inq_ary[5][41] ) );
  LATCHX1_RVT \inq_ary_reg[6][41]  ( .CLK(n3485), .D(n3378), .Q(
        \inq_ary[6][41] ) );
  LATCHX1_RVT \inq_ary_reg[7][41]  ( .CLK(n3484), .D(n3378), .Q(
        \inq_ary[7][41] ) );
  LATCHX1_RVT \inq_ary_reg[8][41]  ( .CLK(n3483), .D(n3378), .Q(
        \inq_ary[8][41] ) );
  LATCHX1_RVT \inq_ary_reg[9][41]  ( .CLK(n3482), .D(n3378), .Q(
        \inq_ary[9][41] ) );
  LATCHX1_RVT \inq_ary_reg[10][41]  ( .CLK(n3481), .D(n3378), .Q(
        \inq_ary[10][41] ) );
  LATCHX1_RVT \inq_ary_reg[11][41]  ( .CLK(n3480), .D(n3378), .Q(
        \inq_ary[11][41] ) );
  LATCHX1_RVT \inq_ary_reg[12][41]  ( .CLK(n3479), .D(n3378), .Q(
        \inq_ary[12][41] ) );
  LATCHX1_RVT \inq_ary_reg[13][41]  ( .CLK(n3478), .D(n3378), .Q(
        \inq_ary[13][41] ) );
  LATCHX1_RVT \inq_ary_reg[14][41]  ( .CLK(n3477), .D(n3378), .Q(
        \inq_ary[14][41] ) );
  LATCHX1_RVT \inq_ary_reg[15][41]  ( .CLK(n3476), .D(n3378), .Q(
        \inq_ary[15][41] ) );
  LATCHX1_RVT \dout_reg[41]  ( .CLK(n3492), .D(N302), .Q(dout[41]) );
  LATCHX1_RVT \inq_ary_reg[0][40]  ( .CLK(n3491), .D(n3376), .Q(
        \inq_ary[0][40] ) );
  LATCHX1_RVT \inq_ary_reg[1][40]  ( .CLK(n3490), .D(n3376), .Q(
        \inq_ary[1][40] ) );
  LATCHX1_RVT \inq_ary_reg[2][40]  ( .CLK(n3489), .D(n3376), .Q(
        \inq_ary[2][40] ) );
  LATCHX1_RVT \inq_ary_reg[3][40]  ( .CLK(n3488), .D(n3376), .Q(
        \inq_ary[3][40] ) );
  LATCHX1_RVT \inq_ary_reg[4][40]  ( .CLK(n3487), .D(n3376), .Q(
        \inq_ary[4][40] ) );
  LATCHX1_RVT \inq_ary_reg[5][40]  ( .CLK(n3486), .D(n3376), .Q(
        \inq_ary[5][40] ) );
  LATCHX1_RVT \inq_ary_reg[6][40]  ( .CLK(n3485), .D(n3376), .Q(
        \inq_ary[6][40] ) );
  LATCHX1_RVT \inq_ary_reg[7][40]  ( .CLK(n3484), .D(n3376), .Q(
        \inq_ary[7][40] ) );
  LATCHX1_RVT \inq_ary_reg[8][40]  ( .CLK(n3483), .D(n3376), .Q(
        \inq_ary[8][40] ) );
  LATCHX1_RVT \inq_ary_reg[9][40]  ( .CLK(n3482), .D(n3376), .Q(
        \inq_ary[9][40] ) );
  LATCHX1_RVT \inq_ary_reg[10][40]  ( .CLK(n3481), .D(n3376), .Q(
        \inq_ary[10][40] ) );
  LATCHX1_RVT \inq_ary_reg[11][40]  ( .CLK(n3480), .D(n3376), .Q(
        \inq_ary[11][40] ) );
  LATCHX1_RVT \inq_ary_reg[12][40]  ( .CLK(n3479), .D(n3376), .Q(
        \inq_ary[12][40] ) );
  LATCHX1_RVT \inq_ary_reg[13][40]  ( .CLK(n3478), .D(n3376), .Q(
        \inq_ary[13][40] ) );
  LATCHX1_RVT \inq_ary_reg[14][40]  ( .CLK(n3477), .D(n3376), .Q(
        \inq_ary[14][40] ) );
  LATCHX1_RVT \inq_ary_reg[15][40]  ( .CLK(n3476), .D(n3376), .Q(
        \inq_ary[15][40] ) );
  LATCHX1_RVT \dout_reg[40]  ( .CLK(n3492), .D(N301), .Q(dout[40]) );
  LATCHX1_RVT \inq_ary_reg[0][39]  ( .CLK(n3491), .D(n3373), .Q(
        \inq_ary[0][39] ) );
  LATCHX1_RVT \inq_ary_reg[1][39]  ( .CLK(n3490), .D(n3373), .Q(
        \inq_ary[1][39] ) );
  LATCHX1_RVT \inq_ary_reg[2][39]  ( .CLK(n3489), .D(n3373), .Q(
        \inq_ary[2][39] ) );
  LATCHX1_RVT \inq_ary_reg[3][39]  ( .CLK(n3488), .D(n3373), .Q(
        \inq_ary[3][39] ) );
  LATCHX1_RVT \inq_ary_reg[4][39]  ( .CLK(n3487), .D(n3373), .Q(
        \inq_ary[4][39] ) );
  LATCHX1_RVT \inq_ary_reg[5][39]  ( .CLK(n3486), .D(n3373), .Q(
        \inq_ary[5][39] ) );
  LATCHX1_RVT \inq_ary_reg[6][39]  ( .CLK(n3485), .D(n3373), .Q(
        \inq_ary[6][39] ) );
  LATCHX1_RVT \inq_ary_reg[7][39]  ( .CLK(n3484), .D(n3373), .Q(
        \inq_ary[7][39] ) );
  LATCHX1_RVT \inq_ary_reg[8][39]  ( .CLK(n3483), .D(n3373), .Q(
        \inq_ary[8][39] ) );
  LATCHX1_RVT \inq_ary_reg[9][39]  ( .CLK(n3482), .D(n3373), .Q(
        \inq_ary[9][39] ) );
  LATCHX1_RVT \inq_ary_reg[10][39]  ( .CLK(n3481), .D(n3373), .Q(
        \inq_ary[10][39] ) );
  LATCHX1_RVT \inq_ary_reg[11][39]  ( .CLK(n3480), .D(n3373), .Q(
        \inq_ary[11][39] ) );
  LATCHX1_RVT \inq_ary_reg[12][39]  ( .CLK(n3479), .D(n3373), .Q(
        \inq_ary[12][39] ) );
  LATCHX1_RVT \inq_ary_reg[13][39]  ( .CLK(n3478), .D(n3373), .Q(
        \inq_ary[13][39] ) );
  LATCHX1_RVT \inq_ary_reg[14][39]  ( .CLK(n3477), .D(n3373), .Q(
        \inq_ary[14][39] ) );
  LATCHX1_RVT \inq_ary_reg[15][39]  ( .CLK(n3476), .D(n3373), .Q(
        \inq_ary[15][39] ) );
  LATCHX1_RVT \dout_reg[39]  ( .CLK(n3492), .D(N300), .Q(dout[39]) );
  LATCHX1_RVT \inq_ary_reg[0][38]  ( .CLK(n3491), .D(n3371), .Q(
        \inq_ary[0][38] ) );
  LATCHX1_RVT \inq_ary_reg[1][38]  ( .CLK(n3490), .D(n3371), .Q(
        \inq_ary[1][38] ) );
  LATCHX1_RVT \inq_ary_reg[2][38]  ( .CLK(n3489), .D(n3371), .Q(
        \inq_ary[2][38] ) );
  LATCHX1_RVT \inq_ary_reg[3][38]  ( .CLK(n3488), .D(n3371), .Q(
        \inq_ary[3][38] ) );
  LATCHX1_RVT \inq_ary_reg[4][38]  ( .CLK(n3487), .D(n3371), .Q(
        \inq_ary[4][38] ) );
  LATCHX1_RVT \inq_ary_reg[5][38]  ( .CLK(n3486), .D(n3371), .Q(
        \inq_ary[5][38] ) );
  LATCHX1_RVT \inq_ary_reg[6][38]  ( .CLK(n3485), .D(n3371), .Q(
        \inq_ary[6][38] ) );
  LATCHX1_RVT \inq_ary_reg[7][38]  ( .CLK(n3484), .D(n3371), .Q(
        \inq_ary[7][38] ) );
  LATCHX1_RVT \inq_ary_reg[8][38]  ( .CLK(n3483), .D(n3371), .Q(
        \inq_ary[8][38] ) );
  LATCHX1_RVT \inq_ary_reg[9][38]  ( .CLK(n3482), .D(n3371), .Q(
        \inq_ary[9][38] ) );
  LATCHX1_RVT \inq_ary_reg[10][38]  ( .CLK(n3481), .D(n3371), .Q(
        \inq_ary[10][38] ) );
  LATCHX1_RVT \inq_ary_reg[11][38]  ( .CLK(n3480), .D(n3371), .Q(
        \inq_ary[11][38] ) );
  LATCHX1_RVT \inq_ary_reg[12][38]  ( .CLK(n3479), .D(n3371), .Q(
        \inq_ary[12][38] ) );
  LATCHX1_RVT \inq_ary_reg[13][38]  ( .CLK(n3478), .D(n3371), .Q(
        \inq_ary[13][38] ) );
  LATCHX1_RVT \inq_ary_reg[14][38]  ( .CLK(n3477), .D(n3371), .Q(
        \inq_ary[14][38] ) );
  LATCHX1_RVT \inq_ary_reg[15][38]  ( .CLK(n3476), .D(n3371), .Q(
        \inq_ary[15][38] ) );
  LATCHX1_RVT \dout_reg[38]  ( .CLK(n3492), .D(N299), .Q(dout[38]) );
  LATCHX1_RVT \inq_ary_reg[0][37]  ( .CLK(n3491), .D(n3369), .Q(
        \inq_ary[0][37] ) );
  LATCHX1_RVT \inq_ary_reg[1][37]  ( .CLK(n3490), .D(n3369), .Q(
        \inq_ary[1][37] ) );
  LATCHX1_RVT \inq_ary_reg[2][37]  ( .CLK(n3489), .D(n3369), .Q(
        \inq_ary[2][37] ) );
  LATCHX1_RVT \inq_ary_reg[3][37]  ( .CLK(n3488), .D(n3369), .Q(
        \inq_ary[3][37] ) );
  LATCHX1_RVT \inq_ary_reg[4][37]  ( .CLK(n3487), .D(n3369), .Q(
        \inq_ary[4][37] ) );
  LATCHX1_RVT \inq_ary_reg[5][37]  ( .CLK(n3486), .D(n3369), .Q(
        \inq_ary[5][37] ) );
  LATCHX1_RVT \inq_ary_reg[6][37]  ( .CLK(n3485), .D(n3369), .Q(
        \inq_ary[6][37] ) );
  LATCHX1_RVT \inq_ary_reg[7][37]  ( .CLK(n3484), .D(n3369), .Q(
        \inq_ary[7][37] ) );
  LATCHX1_RVT \inq_ary_reg[8][37]  ( .CLK(n3483), .D(n3369), .Q(
        \inq_ary[8][37] ) );
  LATCHX1_RVT \inq_ary_reg[9][37]  ( .CLK(n3482), .D(n3369), .Q(
        \inq_ary[9][37] ) );
  LATCHX1_RVT \inq_ary_reg[10][37]  ( .CLK(n3481), .D(n3369), .Q(
        \inq_ary[10][37] ) );
  LATCHX1_RVT \inq_ary_reg[11][37]  ( .CLK(n3480), .D(n3369), .Q(
        \inq_ary[11][37] ) );
  LATCHX1_RVT \inq_ary_reg[12][37]  ( .CLK(n3479), .D(n3369), .Q(
        \inq_ary[12][37] ) );
  LATCHX1_RVT \inq_ary_reg[13][37]  ( .CLK(n3478), .D(n3369), .Q(
        \inq_ary[13][37] ) );
  LATCHX1_RVT \inq_ary_reg[14][37]  ( .CLK(n3477), .D(n3369), .Q(
        \inq_ary[14][37] ) );
  LATCHX1_RVT \inq_ary_reg[15][37]  ( .CLK(n3476), .D(n3369), .Q(
        \inq_ary[15][37] ) );
  LATCHX1_RVT \dout_reg[37]  ( .CLK(n3492), .D(N298), .Q(dout[37]) );
  LATCHX1_RVT \inq_ary_reg[0][36]  ( .CLK(n3491), .D(n3367), .Q(
        \inq_ary[0][36] ) );
  LATCHX1_RVT \inq_ary_reg[1][36]  ( .CLK(n3490), .D(n3367), .Q(
        \inq_ary[1][36] ) );
  LATCHX1_RVT \inq_ary_reg[2][36]  ( .CLK(n3489), .D(n3367), .Q(
        \inq_ary[2][36] ) );
  LATCHX1_RVT \inq_ary_reg[3][36]  ( .CLK(n3488), .D(n3367), .Q(
        \inq_ary[3][36] ) );
  LATCHX1_RVT \inq_ary_reg[4][36]  ( .CLK(n3487), .D(n3367), .Q(
        \inq_ary[4][36] ) );
  LATCHX1_RVT \inq_ary_reg[5][36]  ( .CLK(n3486), .D(n3367), .Q(
        \inq_ary[5][36] ) );
  LATCHX1_RVT \inq_ary_reg[6][36]  ( .CLK(n3485), .D(n3367), .Q(
        \inq_ary[6][36] ) );
  LATCHX1_RVT \inq_ary_reg[7][36]  ( .CLK(n3484), .D(n3367), .Q(
        \inq_ary[7][36] ) );
  LATCHX1_RVT \inq_ary_reg[8][36]  ( .CLK(n3483), .D(n3367), .Q(
        \inq_ary[8][36] ) );
  LATCHX1_RVT \inq_ary_reg[9][36]  ( .CLK(n3482), .D(n3367), .Q(
        \inq_ary[9][36] ) );
  LATCHX1_RVT \inq_ary_reg[10][36]  ( .CLK(n3481), .D(n3367), .Q(
        \inq_ary[10][36] ) );
  LATCHX1_RVT \inq_ary_reg[11][36]  ( .CLK(n3480), .D(n3367), .Q(
        \inq_ary[11][36] ) );
  LATCHX1_RVT \inq_ary_reg[12][36]  ( .CLK(n3479), .D(n3367), .Q(
        \inq_ary[12][36] ) );
  LATCHX1_RVT \inq_ary_reg[13][36]  ( .CLK(n3478), .D(n3367), .Q(
        \inq_ary[13][36] ) );
  LATCHX1_RVT \inq_ary_reg[14][36]  ( .CLK(n3477), .D(n3367), .Q(
        \inq_ary[14][36] ) );
  LATCHX1_RVT \inq_ary_reg[15][36]  ( .CLK(n3476), .D(n3367), .Q(
        \inq_ary[15][36] ) );
  LATCHX1_RVT \dout_reg[36]  ( .CLK(n3492), .D(N297), .Q(dout[36]) );
  LATCHX1_RVT \inq_ary_reg[0][35]  ( .CLK(n3491), .D(n3374), .Q(
        \inq_ary[0][35] ) );
  LATCHX1_RVT \inq_ary_reg[1][35]  ( .CLK(n3490), .D(n3374), .Q(
        \inq_ary[1][35] ) );
  LATCHX1_RVT \inq_ary_reg[2][35]  ( .CLK(n3489), .D(n3374), .Q(
        \inq_ary[2][35] ) );
  LATCHX1_RVT \inq_ary_reg[3][35]  ( .CLK(n3488), .D(n3374), .Q(
        \inq_ary[3][35] ) );
  LATCHX1_RVT \inq_ary_reg[4][35]  ( .CLK(n3487), .D(n3374), .Q(
        \inq_ary[4][35] ) );
  LATCHX1_RVT \inq_ary_reg[5][35]  ( .CLK(n3486), .D(n3374), .Q(
        \inq_ary[5][35] ) );
  LATCHX1_RVT \inq_ary_reg[6][35]  ( .CLK(n3485), .D(n3374), .Q(
        \inq_ary[6][35] ) );
  LATCHX1_RVT \inq_ary_reg[7][35]  ( .CLK(n3484), .D(n3374), .Q(
        \inq_ary[7][35] ) );
  LATCHX1_RVT \inq_ary_reg[8][35]  ( .CLK(n3483), .D(n3374), .Q(
        \inq_ary[8][35] ) );
  LATCHX1_RVT \inq_ary_reg[9][35]  ( .CLK(n3482), .D(n3374), .Q(
        \inq_ary[9][35] ) );
  LATCHX1_RVT \inq_ary_reg[10][35]  ( .CLK(n3481), .D(n3374), .Q(
        \inq_ary[10][35] ) );
  LATCHX1_RVT \inq_ary_reg[11][35]  ( .CLK(n3480), .D(n3374), .Q(
        \inq_ary[11][35] ) );
  LATCHX1_RVT \inq_ary_reg[12][35]  ( .CLK(n3479), .D(n3374), .Q(
        \inq_ary[12][35] ) );
  LATCHX1_RVT \inq_ary_reg[13][35]  ( .CLK(n3478), .D(n3374), .Q(
        \inq_ary[13][35] ) );
  LATCHX1_RVT \inq_ary_reg[14][35]  ( .CLK(n3477), .D(n3374), .Q(
        \inq_ary[14][35] ) );
  LATCHX1_RVT \inq_ary_reg[15][35]  ( .CLK(n3476), .D(n3374), .Q(
        \inq_ary[15][35] ) );
  LATCHX1_RVT \dout_reg[35]  ( .CLK(n3492), .D(N296), .Q(dout[35]) );
  LATCHX1_RVT \inq_ary_reg[0][34]  ( .CLK(n3491), .D(n3372), .Q(
        \inq_ary[0][34] ) );
  LATCHX1_RVT \inq_ary_reg[1][34]  ( .CLK(n3490), .D(n3372), .Q(
        \inq_ary[1][34] ) );
  LATCHX1_RVT \inq_ary_reg[2][34]  ( .CLK(n3489), .D(n3372), .Q(
        \inq_ary[2][34] ) );
  LATCHX1_RVT \inq_ary_reg[3][34]  ( .CLK(n3488), .D(n3372), .Q(
        \inq_ary[3][34] ) );
  LATCHX1_RVT \inq_ary_reg[4][34]  ( .CLK(n3487), .D(n3372), .Q(
        \inq_ary[4][34] ) );
  LATCHX1_RVT \inq_ary_reg[5][34]  ( .CLK(n3486), .D(n3372), .Q(
        \inq_ary[5][34] ) );
  LATCHX1_RVT \inq_ary_reg[6][34]  ( .CLK(n3485), .D(n3372), .Q(
        \inq_ary[6][34] ) );
  LATCHX1_RVT \inq_ary_reg[7][34]  ( .CLK(n3484), .D(n3372), .Q(
        \inq_ary[7][34] ) );
  LATCHX1_RVT \inq_ary_reg[8][34]  ( .CLK(n3483), .D(n3372), .Q(
        \inq_ary[8][34] ) );
  LATCHX1_RVT \inq_ary_reg[9][34]  ( .CLK(n3482), .D(n3372), .Q(
        \inq_ary[9][34] ) );
  LATCHX1_RVT \inq_ary_reg[10][34]  ( .CLK(n3481), .D(n3372), .Q(
        \inq_ary[10][34] ) );
  LATCHX1_RVT \inq_ary_reg[11][34]  ( .CLK(n3480), .D(n3372), .Q(
        \inq_ary[11][34] ) );
  LATCHX1_RVT \inq_ary_reg[12][34]  ( .CLK(n3479), .D(n3372), .Q(
        \inq_ary[12][34] ) );
  LATCHX1_RVT \inq_ary_reg[13][34]  ( .CLK(n3478), .D(n3372), .Q(
        \inq_ary[13][34] ) );
  LATCHX1_RVT \inq_ary_reg[14][34]  ( .CLK(n3477), .D(n3372), .Q(
        \inq_ary[14][34] ) );
  LATCHX1_RVT \inq_ary_reg[15][34]  ( .CLK(n3476), .D(n3372), .Q(
        \inq_ary[15][34] ) );
  LATCHX1_RVT \dout_reg[34]  ( .CLK(n3492), .D(N295), .Q(dout[34]) );
  LATCHX1_RVT \inq_ary_reg[0][33]  ( .CLK(n3491), .D(n3370), .Q(
        \inq_ary[0][33] ) );
  LATCHX1_RVT \inq_ary_reg[1][33]  ( .CLK(n3490), .D(n3370), .Q(
        \inq_ary[1][33] ) );
  LATCHX1_RVT \inq_ary_reg[2][33]  ( .CLK(n3489), .D(n3370), .Q(
        \inq_ary[2][33] ) );
  LATCHX1_RVT \inq_ary_reg[3][33]  ( .CLK(n3488), .D(n3370), .Q(
        \inq_ary[3][33] ) );
  LATCHX1_RVT \inq_ary_reg[4][33]  ( .CLK(n3487), .D(n3370), .Q(
        \inq_ary[4][33] ) );
  LATCHX1_RVT \inq_ary_reg[5][33]  ( .CLK(n3486), .D(n3370), .Q(
        \inq_ary[5][33] ) );
  LATCHX1_RVT \inq_ary_reg[6][33]  ( .CLK(n3485), .D(n3370), .Q(
        \inq_ary[6][33] ) );
  LATCHX1_RVT \inq_ary_reg[7][33]  ( .CLK(n3484), .D(n3370), .Q(
        \inq_ary[7][33] ) );
  LATCHX1_RVT \inq_ary_reg[8][33]  ( .CLK(n3483), .D(n3370), .Q(
        \inq_ary[8][33] ) );
  LATCHX1_RVT \inq_ary_reg[9][33]  ( .CLK(n3482), .D(n3370), .Q(
        \inq_ary[9][33] ) );
  LATCHX1_RVT \inq_ary_reg[10][33]  ( .CLK(n3481), .D(n3370), .Q(
        \inq_ary[10][33] ) );
  LATCHX1_RVT \inq_ary_reg[11][33]  ( .CLK(n3480), .D(n3370), .Q(
        \inq_ary[11][33] ) );
  LATCHX1_RVT \inq_ary_reg[12][33]  ( .CLK(n3479), .D(n3370), .Q(
        \inq_ary[12][33] ) );
  LATCHX1_RVT \inq_ary_reg[13][33]  ( .CLK(n3478), .D(n3370), .Q(
        \inq_ary[13][33] ) );
  LATCHX1_RVT \inq_ary_reg[14][33]  ( .CLK(n3477), .D(n3370), .Q(
        \inq_ary[14][33] ) );
  LATCHX1_RVT \inq_ary_reg[15][33]  ( .CLK(n3476), .D(n3370), .Q(
        \inq_ary[15][33] ) );
  LATCHX1_RVT \dout_reg[33]  ( .CLK(n3492), .D(N294), .Q(dout[33]) );
  LATCHX1_RVT \inq_ary_reg[0][32]  ( .CLK(n3491), .D(n3368), .Q(
        \inq_ary[0][32] ) );
  LATCHX1_RVT \inq_ary_reg[1][32]  ( .CLK(n3490), .D(n3368), .Q(
        \inq_ary[1][32] ) );
  LATCHX1_RVT \inq_ary_reg[2][32]  ( .CLK(n3489), .D(n3368), .Q(
        \inq_ary[2][32] ) );
  LATCHX1_RVT \inq_ary_reg[3][32]  ( .CLK(n3488), .D(n3368), .Q(
        \inq_ary[3][32] ) );
  LATCHX1_RVT \inq_ary_reg[4][32]  ( .CLK(n3487), .D(n3368), .Q(
        \inq_ary[4][32] ) );
  LATCHX1_RVT \inq_ary_reg[5][32]  ( .CLK(n3486), .D(n3368), .Q(
        \inq_ary[5][32] ) );
  LATCHX1_RVT \inq_ary_reg[6][32]  ( .CLK(n3485), .D(n3368), .Q(
        \inq_ary[6][32] ) );
  LATCHX1_RVT \inq_ary_reg[7][32]  ( .CLK(n3484), .D(n3368), .Q(
        \inq_ary[7][32] ) );
  LATCHX1_RVT \inq_ary_reg[8][32]  ( .CLK(n3483), .D(n3368), .Q(
        \inq_ary[8][32] ) );
  LATCHX1_RVT \inq_ary_reg[9][32]  ( .CLK(n3482), .D(n3368), .Q(
        \inq_ary[9][32] ) );
  LATCHX1_RVT \inq_ary_reg[10][32]  ( .CLK(n3481), .D(n3368), .Q(
        \inq_ary[10][32] ) );
  LATCHX1_RVT \inq_ary_reg[11][32]  ( .CLK(n3480), .D(n3368), .Q(
        \inq_ary[11][32] ) );
  LATCHX1_RVT \inq_ary_reg[12][32]  ( .CLK(n3479), .D(n3368), .Q(
        \inq_ary[12][32] ) );
  LATCHX1_RVT \inq_ary_reg[13][32]  ( .CLK(n3478), .D(n3368), .Q(
        \inq_ary[13][32] ) );
  LATCHX1_RVT \inq_ary_reg[14][32]  ( .CLK(n3477), .D(n3368), .Q(
        \inq_ary[14][32] ) );
  LATCHX1_RVT \inq_ary_reg[15][32]  ( .CLK(n3476), .D(n3368), .Q(
        \inq_ary[15][32] ) );
  LATCHX1_RVT \dout_reg[32]  ( .CLK(n3492), .D(N293), .Q(dout[32]) );
  LATCHX1_RVT \inq_ary_reg[0][31]  ( .CLK(n3491), .D(n3365), .Q(
        \inq_ary[0][31] ) );
  LATCHX1_RVT \inq_ary_reg[1][31]  ( .CLK(n3490), .D(n3365), .Q(
        \inq_ary[1][31] ) );
  LATCHX1_RVT \inq_ary_reg[2][31]  ( .CLK(n3489), .D(n3365), .Q(
        \inq_ary[2][31] ) );
  LATCHX1_RVT \inq_ary_reg[3][31]  ( .CLK(n3488), .D(n3365), .Q(
        \inq_ary[3][31] ) );
  LATCHX1_RVT \inq_ary_reg[4][31]  ( .CLK(n3487), .D(n3365), .Q(
        \inq_ary[4][31] ) );
  LATCHX1_RVT \inq_ary_reg[5][31]  ( .CLK(n3486), .D(n3365), .Q(
        \inq_ary[5][31] ) );
  LATCHX1_RVT \inq_ary_reg[6][31]  ( .CLK(n3485), .D(n3365), .Q(
        \inq_ary[6][31] ) );
  LATCHX1_RVT \inq_ary_reg[7][31]  ( .CLK(n3484), .D(n3365), .Q(
        \inq_ary[7][31] ) );
  LATCHX1_RVT \inq_ary_reg[8][31]  ( .CLK(n3483), .D(n3365), .Q(
        \inq_ary[8][31] ) );
  LATCHX1_RVT \inq_ary_reg[9][31]  ( .CLK(n3482), .D(n3365), .Q(
        \inq_ary[9][31] ) );
  LATCHX1_RVT \inq_ary_reg[10][31]  ( .CLK(n3481), .D(n3365), .Q(
        \inq_ary[10][31] ) );
  LATCHX1_RVT \inq_ary_reg[11][31]  ( .CLK(n3480), .D(n3365), .Q(
        \inq_ary[11][31] ) );
  LATCHX1_RVT \inq_ary_reg[12][31]  ( .CLK(n3479), .D(n3365), .Q(
        \inq_ary[12][31] ) );
  LATCHX1_RVT \inq_ary_reg[13][31]  ( .CLK(n3478), .D(n3365), .Q(
        \inq_ary[13][31] ) );
  LATCHX1_RVT \inq_ary_reg[14][31]  ( .CLK(n3477), .D(n3365), .Q(
        \inq_ary[14][31] ) );
  LATCHX1_RVT \inq_ary_reg[15][31]  ( .CLK(n3476), .D(n3365), .Q(
        \inq_ary[15][31] ) );
  LATCHX1_RVT \dout_reg[31]  ( .CLK(n3492), .D(N292), .Q(dout[31]) );
  LATCHX1_RVT \inq_ary_reg[0][30]  ( .CLK(n3491), .D(n3363), .Q(
        \inq_ary[0][30] ) );
  LATCHX1_RVT \inq_ary_reg[1][30]  ( .CLK(n3490), .D(n3363), .Q(
        \inq_ary[1][30] ) );
  LATCHX1_RVT \inq_ary_reg[2][30]  ( .CLK(n3489), .D(n3363), .Q(
        \inq_ary[2][30] ) );
  LATCHX1_RVT \inq_ary_reg[3][30]  ( .CLK(n3488), .D(n3363), .Q(
        \inq_ary[3][30] ) );
  LATCHX1_RVT \inq_ary_reg[4][30]  ( .CLK(n3487), .D(n3363), .Q(
        \inq_ary[4][30] ) );
  LATCHX1_RVT \inq_ary_reg[5][30]  ( .CLK(n3486), .D(n3363), .Q(
        \inq_ary[5][30] ) );
  LATCHX1_RVT \inq_ary_reg[6][30]  ( .CLK(n3485), .D(n3363), .Q(
        \inq_ary[6][30] ) );
  LATCHX1_RVT \inq_ary_reg[7][30]  ( .CLK(n3484), .D(n3363), .Q(
        \inq_ary[7][30] ) );
  LATCHX1_RVT \inq_ary_reg[8][30]  ( .CLK(n3483), .D(n3363), .Q(
        \inq_ary[8][30] ) );
  LATCHX1_RVT \inq_ary_reg[9][30]  ( .CLK(n3482), .D(n3363), .Q(
        \inq_ary[9][30] ) );
  LATCHX1_RVT \inq_ary_reg[10][30]  ( .CLK(n3481), .D(n3363), .Q(
        \inq_ary[10][30] ) );
  LATCHX1_RVT \inq_ary_reg[11][30]  ( .CLK(n3480), .D(n3363), .Q(
        \inq_ary[11][30] ) );
  LATCHX1_RVT \inq_ary_reg[12][30]  ( .CLK(n3479), .D(n3363), .Q(
        \inq_ary[12][30] ) );
  LATCHX1_RVT \inq_ary_reg[13][30]  ( .CLK(n3478), .D(n3363), .Q(
        \inq_ary[13][30] ) );
  LATCHX1_RVT \inq_ary_reg[14][30]  ( .CLK(n3477), .D(n3363), .Q(
        \inq_ary[14][30] ) );
  LATCHX1_RVT \inq_ary_reg[15][30]  ( .CLK(n3476), .D(n3363), .Q(
        \inq_ary[15][30] ) );
  LATCHX1_RVT \dout_reg[30]  ( .CLK(n3492), .D(N291), .Q(dout[30]) );
  LATCHX1_RVT \inq_ary_reg[0][29]  ( .CLK(n3491), .D(n3361), .Q(
        \inq_ary[0][29] ) );
  LATCHX1_RVT \inq_ary_reg[1][29]  ( .CLK(n3490), .D(n3361), .Q(
        \inq_ary[1][29] ) );
  LATCHX1_RVT \inq_ary_reg[2][29]  ( .CLK(n3489), .D(n3361), .Q(
        \inq_ary[2][29] ) );
  LATCHX1_RVT \inq_ary_reg[3][29]  ( .CLK(n3488), .D(n3361), .Q(
        \inq_ary[3][29] ) );
  LATCHX1_RVT \inq_ary_reg[4][29]  ( .CLK(n3487), .D(n3361), .Q(
        \inq_ary[4][29] ) );
  LATCHX1_RVT \inq_ary_reg[5][29]  ( .CLK(n3486), .D(n3361), .Q(
        \inq_ary[5][29] ) );
  LATCHX1_RVT \inq_ary_reg[6][29]  ( .CLK(n3485), .D(n3361), .Q(
        \inq_ary[6][29] ) );
  LATCHX1_RVT \inq_ary_reg[7][29]  ( .CLK(n3484), .D(n3361), .Q(
        \inq_ary[7][29] ) );
  LATCHX1_RVT \inq_ary_reg[8][29]  ( .CLK(n3483), .D(n3361), .Q(
        \inq_ary[8][29] ) );
  LATCHX1_RVT \inq_ary_reg[9][29]  ( .CLK(n3482), .D(n3361), .Q(
        \inq_ary[9][29] ) );
  LATCHX1_RVT \inq_ary_reg[10][29]  ( .CLK(n3481), .D(n3361), .Q(
        \inq_ary[10][29] ) );
  LATCHX1_RVT \inq_ary_reg[11][29]  ( .CLK(n3480), .D(n3361), .Q(
        \inq_ary[11][29] ) );
  LATCHX1_RVT \inq_ary_reg[12][29]  ( .CLK(n3479), .D(n3361), .Q(
        \inq_ary[12][29] ) );
  LATCHX1_RVT \inq_ary_reg[13][29]  ( .CLK(n3478), .D(n3361), .Q(
        \inq_ary[13][29] ) );
  LATCHX1_RVT \inq_ary_reg[14][29]  ( .CLK(n3477), .D(n3361), .Q(
        \inq_ary[14][29] ) );
  LATCHX1_RVT \inq_ary_reg[15][29]  ( .CLK(n3476), .D(n3361), .Q(
        \inq_ary[15][29] ) );
  LATCHX1_RVT \dout_reg[29]  ( .CLK(n3492), .D(N290), .Q(dout[29]) );
  LATCHX1_RVT \inq_ary_reg[0][28]  ( .CLK(n3491), .D(n3359), .Q(
        \inq_ary[0][28] ) );
  LATCHX1_RVT \inq_ary_reg[1][28]  ( .CLK(n3490), .D(n3359), .Q(
        \inq_ary[1][28] ) );
  LATCHX1_RVT \inq_ary_reg[2][28]  ( .CLK(n3489), .D(n3359), .Q(
        \inq_ary[2][28] ) );
  LATCHX1_RVT \inq_ary_reg[3][28]  ( .CLK(n3488), .D(n3359), .Q(
        \inq_ary[3][28] ) );
  LATCHX1_RVT \inq_ary_reg[4][28]  ( .CLK(n3487), .D(n3359), .Q(
        \inq_ary[4][28] ) );
  LATCHX1_RVT \inq_ary_reg[5][28]  ( .CLK(n3486), .D(n3359), .Q(
        \inq_ary[5][28] ) );
  LATCHX1_RVT \inq_ary_reg[6][28]  ( .CLK(n3485), .D(n3359), .Q(
        \inq_ary[6][28] ) );
  LATCHX1_RVT \inq_ary_reg[7][28]  ( .CLK(n3484), .D(n3359), .Q(
        \inq_ary[7][28] ) );
  LATCHX1_RVT \inq_ary_reg[8][28]  ( .CLK(n3483), .D(n3359), .Q(
        \inq_ary[8][28] ) );
  LATCHX1_RVT \inq_ary_reg[9][28]  ( .CLK(n3482), .D(n3359), .Q(
        \inq_ary[9][28] ) );
  LATCHX1_RVT \inq_ary_reg[10][28]  ( .CLK(n3481), .D(n3359), .Q(
        \inq_ary[10][28] ) );
  LATCHX1_RVT \inq_ary_reg[11][28]  ( .CLK(n3480), .D(n3359), .Q(
        \inq_ary[11][28] ) );
  LATCHX1_RVT \inq_ary_reg[12][28]  ( .CLK(n3479), .D(n3359), .Q(
        \inq_ary[12][28] ) );
  LATCHX1_RVT \inq_ary_reg[13][28]  ( .CLK(n3478), .D(n3359), .Q(
        \inq_ary[13][28] ) );
  LATCHX1_RVT \inq_ary_reg[14][28]  ( .CLK(n3477), .D(n3359), .Q(
        \inq_ary[14][28] ) );
  LATCHX1_RVT \inq_ary_reg[15][28]  ( .CLK(n3476), .D(n3359), .Q(
        \inq_ary[15][28] ) );
  LATCHX1_RVT \dout_reg[28]  ( .CLK(n3492), .D(N289), .Q(dout[28]) );
  LATCHX1_RVT \inq_ary_reg[0][27]  ( .CLK(n3491), .D(n3366), .Q(
        \inq_ary[0][27] ) );
  LATCHX1_RVT \inq_ary_reg[1][27]  ( .CLK(n3490), .D(n3366), .Q(
        \inq_ary[1][27] ) );
  LATCHX1_RVT \inq_ary_reg[2][27]  ( .CLK(n3489), .D(n3366), .Q(
        \inq_ary[2][27] ) );
  LATCHX1_RVT \inq_ary_reg[3][27]  ( .CLK(n3488), .D(n3366), .Q(
        \inq_ary[3][27] ) );
  LATCHX1_RVT \inq_ary_reg[4][27]  ( .CLK(n3487), .D(n3366), .Q(
        \inq_ary[4][27] ) );
  LATCHX1_RVT \inq_ary_reg[5][27]  ( .CLK(n3486), .D(n3366), .Q(
        \inq_ary[5][27] ) );
  LATCHX1_RVT \inq_ary_reg[6][27]  ( .CLK(n3485), .D(n3366), .Q(
        \inq_ary[6][27] ) );
  LATCHX1_RVT \inq_ary_reg[7][27]  ( .CLK(n3484), .D(n3366), .Q(
        \inq_ary[7][27] ) );
  LATCHX1_RVT \inq_ary_reg[8][27]  ( .CLK(n3483), .D(n3366), .Q(
        \inq_ary[8][27] ) );
  LATCHX1_RVT \inq_ary_reg[9][27]  ( .CLK(n3482), .D(n3366), .Q(
        \inq_ary[9][27] ) );
  LATCHX1_RVT \inq_ary_reg[10][27]  ( .CLK(n3481), .D(n3366), .Q(
        \inq_ary[10][27] ) );
  LATCHX1_RVT \inq_ary_reg[11][27]  ( .CLK(n3480), .D(n3366), .Q(
        \inq_ary[11][27] ) );
  LATCHX1_RVT \inq_ary_reg[12][27]  ( .CLK(n3479), .D(n3366), .Q(
        \inq_ary[12][27] ) );
  LATCHX1_RVT \inq_ary_reg[13][27]  ( .CLK(n3478), .D(n3366), .Q(
        \inq_ary[13][27] ) );
  LATCHX1_RVT \inq_ary_reg[14][27]  ( .CLK(n3477), .D(n3366), .Q(
        \inq_ary[14][27] ) );
  LATCHX1_RVT \inq_ary_reg[15][27]  ( .CLK(n3476), .D(n3366), .Q(
        \inq_ary[15][27] ) );
  LATCHX1_RVT \dout_reg[27]  ( .CLK(n3492), .D(N288), .Q(dout[27]) );
  LATCHX1_RVT \inq_ary_reg[0][26]  ( .CLK(n3491), .D(n3364), .Q(
        \inq_ary[0][26] ) );
  LATCHX1_RVT \inq_ary_reg[1][26]  ( .CLK(n3490), .D(n3364), .Q(
        \inq_ary[1][26] ) );
  LATCHX1_RVT \inq_ary_reg[2][26]  ( .CLK(n3489), .D(n3364), .Q(
        \inq_ary[2][26] ) );
  LATCHX1_RVT \inq_ary_reg[3][26]  ( .CLK(n3488), .D(n3364), .Q(
        \inq_ary[3][26] ) );
  LATCHX1_RVT \inq_ary_reg[4][26]  ( .CLK(n3487), .D(n3364), .Q(
        \inq_ary[4][26] ) );
  LATCHX1_RVT \inq_ary_reg[5][26]  ( .CLK(n3486), .D(n3364), .Q(
        \inq_ary[5][26] ) );
  LATCHX1_RVT \inq_ary_reg[6][26]  ( .CLK(n3485), .D(n3364), .Q(
        \inq_ary[6][26] ) );
  LATCHX1_RVT \inq_ary_reg[7][26]  ( .CLK(n3484), .D(n3364), .Q(
        \inq_ary[7][26] ) );
  LATCHX1_RVT \inq_ary_reg[8][26]  ( .CLK(n3483), .D(n3364), .Q(
        \inq_ary[8][26] ) );
  LATCHX1_RVT \inq_ary_reg[9][26]  ( .CLK(n3482), .D(n3364), .Q(
        \inq_ary[9][26] ) );
  LATCHX1_RVT \inq_ary_reg[10][26]  ( .CLK(n3481), .D(n3364), .Q(
        \inq_ary[10][26] ) );
  LATCHX1_RVT \inq_ary_reg[11][26]  ( .CLK(n3480), .D(n3364), .Q(
        \inq_ary[11][26] ) );
  LATCHX1_RVT \inq_ary_reg[12][26]  ( .CLK(n3479), .D(n3364), .Q(
        \inq_ary[12][26] ) );
  LATCHX1_RVT \inq_ary_reg[13][26]  ( .CLK(n3478), .D(n3364), .Q(
        \inq_ary[13][26] ) );
  LATCHX1_RVT \inq_ary_reg[14][26]  ( .CLK(n3477), .D(n3364), .Q(
        \inq_ary[14][26] ) );
  LATCHX1_RVT \inq_ary_reg[15][26]  ( .CLK(n3476), .D(n3364), .Q(
        \inq_ary[15][26] ) );
  LATCHX1_RVT \dout_reg[26]  ( .CLK(n3492), .D(N287), .Q(dout[26]) );
  LATCHX1_RVT \inq_ary_reg[0][25]  ( .CLK(n3491), .D(n3362), .Q(
        \inq_ary[0][25] ) );
  LATCHX1_RVT \inq_ary_reg[1][25]  ( .CLK(n3490), .D(n3362), .Q(
        \inq_ary[1][25] ) );
  LATCHX1_RVT \inq_ary_reg[2][25]  ( .CLK(n3489), .D(n3362), .Q(
        \inq_ary[2][25] ) );
  LATCHX1_RVT \inq_ary_reg[3][25]  ( .CLK(n3488), .D(n3362), .Q(
        \inq_ary[3][25] ) );
  LATCHX1_RVT \inq_ary_reg[4][25]  ( .CLK(n3487), .D(n3362), .Q(
        \inq_ary[4][25] ) );
  LATCHX1_RVT \inq_ary_reg[5][25]  ( .CLK(n3486), .D(n3362), .Q(
        \inq_ary[5][25] ) );
  LATCHX1_RVT \inq_ary_reg[6][25]  ( .CLK(n3485), .D(n3362), .Q(
        \inq_ary[6][25] ) );
  LATCHX1_RVT \inq_ary_reg[7][25]  ( .CLK(n3484), .D(n3362), .Q(
        \inq_ary[7][25] ) );
  LATCHX1_RVT \inq_ary_reg[8][25]  ( .CLK(n3483), .D(n3362), .Q(
        \inq_ary[8][25] ) );
  LATCHX1_RVT \inq_ary_reg[9][25]  ( .CLK(n3482), .D(n3362), .Q(
        \inq_ary[9][25] ) );
  LATCHX1_RVT \inq_ary_reg[10][25]  ( .CLK(n3481), .D(n3362), .Q(
        \inq_ary[10][25] ) );
  LATCHX1_RVT \inq_ary_reg[11][25]  ( .CLK(n3480), .D(n3362), .Q(
        \inq_ary[11][25] ) );
  LATCHX1_RVT \inq_ary_reg[12][25]  ( .CLK(n3479), .D(n3362), .Q(
        \inq_ary[12][25] ) );
  LATCHX1_RVT \inq_ary_reg[13][25]  ( .CLK(n3478), .D(n3362), .Q(
        \inq_ary[13][25] ) );
  LATCHX1_RVT \inq_ary_reg[14][25]  ( .CLK(n3477), .D(n3362), .Q(
        \inq_ary[14][25] ) );
  LATCHX1_RVT \inq_ary_reg[15][25]  ( .CLK(n3476), .D(n3362), .Q(
        \inq_ary[15][25] ) );
  LATCHX1_RVT \dout_reg[25]  ( .CLK(n3492), .D(N286), .Q(dout[25]) );
  LATCHX1_RVT \inq_ary_reg[0][24]  ( .CLK(n3491), .D(n3360), .Q(
        \inq_ary[0][24] ) );
  LATCHX1_RVT \inq_ary_reg[1][24]  ( .CLK(n3490), .D(n3360), .Q(
        \inq_ary[1][24] ) );
  LATCHX1_RVT \inq_ary_reg[2][24]  ( .CLK(n3489), .D(n3360), .Q(
        \inq_ary[2][24] ) );
  LATCHX1_RVT \inq_ary_reg[3][24]  ( .CLK(n3488), .D(n3360), .Q(
        \inq_ary[3][24] ) );
  LATCHX1_RVT \inq_ary_reg[4][24]  ( .CLK(n3487), .D(n3360), .Q(
        \inq_ary[4][24] ) );
  LATCHX1_RVT \inq_ary_reg[5][24]  ( .CLK(n3486), .D(n3360), .Q(
        \inq_ary[5][24] ) );
  LATCHX1_RVT \inq_ary_reg[6][24]  ( .CLK(n3485), .D(n3360), .Q(
        \inq_ary[6][24] ) );
  LATCHX1_RVT \inq_ary_reg[7][24]  ( .CLK(n3484), .D(n3360), .Q(
        \inq_ary[7][24] ) );
  LATCHX1_RVT \inq_ary_reg[8][24]  ( .CLK(n3483), .D(n3360), .Q(
        \inq_ary[8][24] ) );
  LATCHX1_RVT \inq_ary_reg[9][24]  ( .CLK(n3482), .D(n3360), .Q(
        \inq_ary[9][24] ) );
  LATCHX1_RVT \inq_ary_reg[10][24]  ( .CLK(n3481), .D(n3360), .Q(
        \inq_ary[10][24] ) );
  LATCHX1_RVT \inq_ary_reg[11][24]  ( .CLK(n3480), .D(n3360), .Q(
        \inq_ary[11][24] ) );
  LATCHX1_RVT \inq_ary_reg[12][24]  ( .CLK(n3479), .D(n3360), .Q(
        \inq_ary[12][24] ) );
  LATCHX1_RVT \inq_ary_reg[13][24]  ( .CLK(n3478), .D(n3360), .Q(
        \inq_ary[13][24] ) );
  LATCHX1_RVT \inq_ary_reg[14][24]  ( .CLK(n3477), .D(n3360), .Q(
        \inq_ary[14][24] ) );
  LATCHX1_RVT \inq_ary_reg[15][24]  ( .CLK(n3476), .D(n3360), .Q(
        \inq_ary[15][24] ) );
  LATCHX1_RVT \dout_reg[24]  ( .CLK(n3492), .D(N285), .Q(dout[24]) );
  LATCHX1_RVT \inq_ary_reg[0][23]  ( .CLK(n3491), .D(n3357), .Q(
        \inq_ary[0][23] ) );
  LATCHX1_RVT \inq_ary_reg[1][23]  ( .CLK(n3490), .D(n3357), .Q(
        \inq_ary[1][23] ) );
  LATCHX1_RVT \inq_ary_reg[2][23]  ( .CLK(n3489), .D(n3357), .Q(
        \inq_ary[2][23] ) );
  LATCHX1_RVT \inq_ary_reg[3][23]  ( .CLK(n3488), .D(n3357), .Q(
        \inq_ary[3][23] ) );
  LATCHX1_RVT \inq_ary_reg[4][23]  ( .CLK(n3487), .D(n3357), .Q(
        \inq_ary[4][23] ) );
  LATCHX1_RVT \inq_ary_reg[5][23]  ( .CLK(n3486), .D(n3357), .Q(
        \inq_ary[5][23] ) );
  LATCHX1_RVT \inq_ary_reg[6][23]  ( .CLK(n3485), .D(n3357), .Q(
        \inq_ary[6][23] ) );
  LATCHX1_RVT \inq_ary_reg[7][23]  ( .CLK(n3484), .D(n3357), .Q(
        \inq_ary[7][23] ) );
  LATCHX1_RVT \inq_ary_reg[8][23]  ( .CLK(n3483), .D(n3357), .Q(
        \inq_ary[8][23] ) );
  LATCHX1_RVT \inq_ary_reg[9][23]  ( .CLK(n3482), .D(n3357), .Q(
        \inq_ary[9][23] ) );
  LATCHX1_RVT \inq_ary_reg[10][23]  ( .CLK(n3481), .D(n3357), .Q(
        \inq_ary[10][23] ) );
  LATCHX1_RVT \inq_ary_reg[11][23]  ( .CLK(n3480), .D(n3357), .Q(
        \inq_ary[11][23] ) );
  LATCHX1_RVT \inq_ary_reg[12][23]  ( .CLK(n3479), .D(n3357), .Q(
        \inq_ary[12][23] ) );
  LATCHX1_RVT \inq_ary_reg[13][23]  ( .CLK(n3478), .D(n3357), .Q(
        \inq_ary[13][23] ) );
  LATCHX1_RVT \inq_ary_reg[14][23]  ( .CLK(n3477), .D(n3357), .Q(
        \inq_ary[14][23] ) );
  LATCHX1_RVT \inq_ary_reg[15][23]  ( .CLK(n3476), .D(n3357), .Q(
        \inq_ary[15][23] ) );
  LATCHX1_RVT \dout_reg[23]  ( .CLK(n3492), .D(N284), .Q(dout[23]) );
  LATCHX1_RVT \inq_ary_reg[0][22]  ( .CLK(n3491), .D(n3355), .Q(
        \inq_ary[0][22] ) );
  LATCHX1_RVT \inq_ary_reg[1][22]  ( .CLK(n3490), .D(n3355), .Q(
        \inq_ary[1][22] ) );
  LATCHX1_RVT \inq_ary_reg[2][22]  ( .CLK(n3489), .D(n3355), .Q(
        \inq_ary[2][22] ) );
  LATCHX1_RVT \inq_ary_reg[3][22]  ( .CLK(n3488), .D(n3355), .Q(
        \inq_ary[3][22] ) );
  LATCHX1_RVT \inq_ary_reg[4][22]  ( .CLK(n3487), .D(n3355), .Q(
        \inq_ary[4][22] ) );
  LATCHX1_RVT \inq_ary_reg[5][22]  ( .CLK(n3486), .D(n3355), .Q(
        \inq_ary[5][22] ) );
  LATCHX1_RVT \inq_ary_reg[6][22]  ( .CLK(n3485), .D(n3355), .Q(
        \inq_ary[6][22] ) );
  LATCHX1_RVT \inq_ary_reg[7][22]  ( .CLK(n3484), .D(n3355), .Q(
        \inq_ary[7][22] ) );
  LATCHX1_RVT \inq_ary_reg[8][22]  ( .CLK(n3483), .D(n3355), .Q(
        \inq_ary[8][22] ) );
  LATCHX1_RVT \inq_ary_reg[9][22]  ( .CLK(n3482), .D(n3355), .Q(
        \inq_ary[9][22] ) );
  LATCHX1_RVT \inq_ary_reg[10][22]  ( .CLK(n3481), .D(n3355), .Q(
        \inq_ary[10][22] ) );
  LATCHX1_RVT \inq_ary_reg[11][22]  ( .CLK(n3480), .D(n3355), .Q(
        \inq_ary[11][22] ) );
  LATCHX1_RVT \inq_ary_reg[12][22]  ( .CLK(n3479), .D(n3355), .Q(
        \inq_ary[12][22] ) );
  LATCHX1_RVT \inq_ary_reg[13][22]  ( .CLK(n3478), .D(n3355), .Q(
        \inq_ary[13][22] ) );
  LATCHX1_RVT \inq_ary_reg[14][22]  ( .CLK(n3477), .D(n3355), .Q(
        \inq_ary[14][22] ) );
  LATCHX1_RVT \inq_ary_reg[15][22]  ( .CLK(n3476), .D(n3355), .Q(
        \inq_ary[15][22] ) );
  LATCHX1_RVT \dout_reg[22]  ( .CLK(n3492), .D(N283), .Q(dout[22]) );
  LATCHX1_RVT \inq_ary_reg[0][21]  ( .CLK(n3491), .D(n3353), .Q(
        \inq_ary[0][21] ) );
  LATCHX1_RVT \inq_ary_reg[1][21]  ( .CLK(n3490), .D(n3353), .Q(
        \inq_ary[1][21] ) );
  LATCHX1_RVT \inq_ary_reg[2][21]  ( .CLK(n3489), .D(n3353), .Q(
        \inq_ary[2][21] ) );
  LATCHX1_RVT \inq_ary_reg[3][21]  ( .CLK(n3488), .D(n3353), .Q(
        \inq_ary[3][21] ) );
  LATCHX1_RVT \inq_ary_reg[4][21]  ( .CLK(n3487), .D(n3353), .Q(
        \inq_ary[4][21] ) );
  LATCHX1_RVT \inq_ary_reg[5][21]  ( .CLK(n3486), .D(n3353), .Q(
        \inq_ary[5][21] ) );
  LATCHX1_RVT \inq_ary_reg[6][21]  ( .CLK(n3485), .D(n3353), .Q(
        \inq_ary[6][21] ) );
  LATCHX1_RVT \inq_ary_reg[7][21]  ( .CLK(n3484), .D(n3353), .Q(
        \inq_ary[7][21] ) );
  LATCHX1_RVT \inq_ary_reg[8][21]  ( .CLK(n3483), .D(n3353), .Q(
        \inq_ary[8][21] ) );
  LATCHX1_RVT \inq_ary_reg[9][21]  ( .CLK(n3482), .D(n3353), .Q(
        \inq_ary[9][21] ) );
  LATCHX1_RVT \inq_ary_reg[10][21]  ( .CLK(n3481), .D(n3353), .Q(
        \inq_ary[10][21] ) );
  LATCHX1_RVT \inq_ary_reg[11][21]  ( .CLK(n3480), .D(n3353), .Q(
        \inq_ary[11][21] ) );
  LATCHX1_RVT \inq_ary_reg[12][21]  ( .CLK(n3479), .D(n3353), .Q(
        \inq_ary[12][21] ) );
  LATCHX1_RVT \inq_ary_reg[13][21]  ( .CLK(n3478), .D(n3353), .Q(
        \inq_ary[13][21] ) );
  LATCHX1_RVT \inq_ary_reg[14][21]  ( .CLK(n3477), .D(n3353), .Q(
        \inq_ary[14][21] ) );
  LATCHX1_RVT \inq_ary_reg[15][21]  ( .CLK(n3476), .D(n3353), .Q(
        \inq_ary[15][21] ) );
  LATCHX1_RVT \dout_reg[21]  ( .CLK(n3492), .D(N282), .Q(dout[21]) );
  LATCHX1_RVT \inq_ary_reg[0][20]  ( .CLK(n3491), .D(n3351), .Q(
        \inq_ary[0][20] ) );
  LATCHX1_RVT \inq_ary_reg[1][20]  ( .CLK(n3490), .D(n3351), .Q(
        \inq_ary[1][20] ) );
  LATCHX1_RVT \inq_ary_reg[2][20]  ( .CLK(n3489), .D(n3351), .Q(
        \inq_ary[2][20] ) );
  LATCHX1_RVT \inq_ary_reg[3][20]  ( .CLK(n3488), .D(n3351), .Q(
        \inq_ary[3][20] ) );
  LATCHX1_RVT \inq_ary_reg[4][20]  ( .CLK(n3487), .D(n3351), .Q(
        \inq_ary[4][20] ) );
  LATCHX1_RVT \inq_ary_reg[5][20]  ( .CLK(n3486), .D(n3351), .Q(
        \inq_ary[5][20] ) );
  LATCHX1_RVT \inq_ary_reg[6][20]  ( .CLK(n3485), .D(n3351), .Q(
        \inq_ary[6][20] ) );
  LATCHX1_RVT \inq_ary_reg[7][20]  ( .CLK(n3484), .D(n3351), .Q(
        \inq_ary[7][20] ) );
  LATCHX1_RVT \inq_ary_reg[8][20]  ( .CLK(n3483), .D(n3351), .Q(
        \inq_ary[8][20] ) );
  LATCHX1_RVT \inq_ary_reg[9][20]  ( .CLK(n3482), .D(n3351), .Q(
        \inq_ary[9][20] ) );
  LATCHX1_RVT \inq_ary_reg[10][20]  ( .CLK(n3481), .D(n3351), .Q(
        \inq_ary[10][20] ) );
  LATCHX1_RVT \inq_ary_reg[11][20]  ( .CLK(n3480), .D(n3351), .Q(
        \inq_ary[11][20] ) );
  LATCHX1_RVT \inq_ary_reg[12][20]  ( .CLK(n3479), .D(n3351), .Q(
        \inq_ary[12][20] ) );
  LATCHX1_RVT \inq_ary_reg[13][20]  ( .CLK(n3478), .D(n3351), .Q(
        \inq_ary[13][20] ) );
  LATCHX1_RVT \inq_ary_reg[14][20]  ( .CLK(n3477), .D(n3351), .Q(
        \inq_ary[14][20] ) );
  LATCHX1_RVT \inq_ary_reg[15][20]  ( .CLK(n3476), .D(n3351), .Q(
        \inq_ary[15][20] ) );
  LATCHX1_RVT \dout_reg[20]  ( .CLK(n3492), .D(N281), .Q(dout[20]) );
  LATCHX1_RVT \inq_ary_reg[0][19]  ( .CLK(n3491), .D(n3358), .Q(
        \inq_ary[0][19] ) );
  LATCHX1_RVT \inq_ary_reg[1][19]  ( .CLK(n3490), .D(n3358), .Q(
        \inq_ary[1][19] ) );
  LATCHX1_RVT \inq_ary_reg[2][19]  ( .CLK(n3489), .D(n3358), .Q(
        \inq_ary[2][19] ) );
  LATCHX1_RVT \inq_ary_reg[3][19]  ( .CLK(n3488), .D(n3358), .Q(
        \inq_ary[3][19] ) );
  LATCHX1_RVT \inq_ary_reg[4][19]  ( .CLK(n3487), .D(n3358), .Q(
        \inq_ary[4][19] ) );
  LATCHX1_RVT \inq_ary_reg[5][19]  ( .CLK(n3486), .D(n3358), .Q(
        \inq_ary[5][19] ) );
  LATCHX1_RVT \inq_ary_reg[6][19]  ( .CLK(n3485), .D(n3358), .Q(
        \inq_ary[6][19] ) );
  LATCHX1_RVT \inq_ary_reg[7][19]  ( .CLK(n3484), .D(n3358), .Q(
        \inq_ary[7][19] ) );
  LATCHX1_RVT \inq_ary_reg[8][19]  ( .CLK(n3483), .D(n3358), .Q(
        \inq_ary[8][19] ) );
  LATCHX1_RVT \inq_ary_reg[9][19]  ( .CLK(n3482), .D(n3358), .Q(
        \inq_ary[9][19] ) );
  LATCHX1_RVT \inq_ary_reg[10][19]  ( .CLK(n3481), .D(n3358), .Q(
        \inq_ary[10][19] ) );
  LATCHX1_RVT \inq_ary_reg[11][19]  ( .CLK(n3480), .D(n3358), .Q(
        \inq_ary[11][19] ) );
  LATCHX1_RVT \inq_ary_reg[12][19]  ( .CLK(n3479), .D(n3358), .Q(
        \inq_ary[12][19] ) );
  LATCHX1_RVT \inq_ary_reg[13][19]  ( .CLK(n3478), .D(n3358), .Q(
        \inq_ary[13][19] ) );
  LATCHX1_RVT \inq_ary_reg[14][19]  ( .CLK(n3477), .D(n3358), .Q(
        \inq_ary[14][19] ) );
  LATCHX1_RVT \inq_ary_reg[15][19]  ( .CLK(n3476), .D(n3358), .Q(
        \inq_ary[15][19] ) );
  LATCHX1_RVT \dout_reg[19]  ( .CLK(n3492), .D(N280), .Q(dout[19]) );
  LATCHX1_RVT \inq_ary_reg[0][18]  ( .CLK(n3491), .D(n3356), .Q(
        \inq_ary[0][18] ) );
  LATCHX1_RVT \inq_ary_reg[1][18]  ( .CLK(n3490), .D(n3356), .Q(
        \inq_ary[1][18] ) );
  LATCHX1_RVT \inq_ary_reg[2][18]  ( .CLK(n3489), .D(n3356), .Q(
        \inq_ary[2][18] ) );
  LATCHX1_RVT \inq_ary_reg[3][18]  ( .CLK(n3488), .D(n3356), .Q(
        \inq_ary[3][18] ) );
  LATCHX1_RVT \inq_ary_reg[4][18]  ( .CLK(n3487), .D(n3356), .Q(
        \inq_ary[4][18] ) );
  LATCHX1_RVT \inq_ary_reg[5][18]  ( .CLK(n3486), .D(n3356), .Q(
        \inq_ary[5][18] ) );
  LATCHX1_RVT \inq_ary_reg[6][18]  ( .CLK(n3485), .D(n3356), .Q(
        \inq_ary[6][18] ) );
  LATCHX1_RVT \inq_ary_reg[7][18]  ( .CLK(n3484), .D(n3356), .Q(
        \inq_ary[7][18] ) );
  LATCHX1_RVT \inq_ary_reg[8][18]  ( .CLK(n3483), .D(n3356), .Q(
        \inq_ary[8][18] ) );
  LATCHX1_RVT \inq_ary_reg[9][18]  ( .CLK(n3482), .D(n3356), .Q(
        \inq_ary[9][18] ) );
  LATCHX1_RVT \inq_ary_reg[10][18]  ( .CLK(n3481), .D(n3356), .Q(
        \inq_ary[10][18] ) );
  LATCHX1_RVT \inq_ary_reg[11][18]  ( .CLK(n3480), .D(n3356), .Q(
        \inq_ary[11][18] ) );
  LATCHX1_RVT \inq_ary_reg[12][18]  ( .CLK(n3479), .D(n3356), .Q(
        \inq_ary[12][18] ) );
  LATCHX1_RVT \inq_ary_reg[13][18]  ( .CLK(n3478), .D(n3356), .Q(
        \inq_ary[13][18] ) );
  LATCHX1_RVT \inq_ary_reg[14][18]  ( .CLK(n3477), .D(n3356), .Q(
        \inq_ary[14][18] ) );
  LATCHX1_RVT \inq_ary_reg[15][18]  ( .CLK(n3476), .D(n3356), .Q(
        \inq_ary[15][18] ) );
  LATCHX1_RVT \dout_reg[18]  ( .CLK(n3492), .D(N279), .Q(dout[18]) );
  LATCHX1_RVT \inq_ary_reg[0][17]  ( .CLK(n3491), .D(n3354), .Q(
        \inq_ary[0][17] ) );
  LATCHX1_RVT \inq_ary_reg[1][17]  ( .CLK(n3490), .D(n3354), .Q(
        \inq_ary[1][17] ) );
  LATCHX1_RVT \inq_ary_reg[2][17]  ( .CLK(n3489), .D(n3354), .Q(
        \inq_ary[2][17] ) );
  LATCHX1_RVT \inq_ary_reg[3][17]  ( .CLK(n3488), .D(n3354), .Q(
        \inq_ary[3][17] ) );
  LATCHX1_RVT \inq_ary_reg[4][17]  ( .CLK(n3487), .D(n3354), .Q(
        \inq_ary[4][17] ) );
  LATCHX1_RVT \inq_ary_reg[5][17]  ( .CLK(n3486), .D(n3354), .Q(
        \inq_ary[5][17] ) );
  LATCHX1_RVT \inq_ary_reg[6][17]  ( .CLK(n3485), .D(n3354), .Q(
        \inq_ary[6][17] ) );
  LATCHX1_RVT \inq_ary_reg[7][17]  ( .CLK(n3484), .D(n3354), .Q(
        \inq_ary[7][17] ) );
  LATCHX1_RVT \inq_ary_reg[8][17]  ( .CLK(n3483), .D(n3354), .Q(
        \inq_ary[8][17] ) );
  LATCHX1_RVT \inq_ary_reg[9][17]  ( .CLK(n3482), .D(n3354), .Q(
        \inq_ary[9][17] ) );
  LATCHX1_RVT \inq_ary_reg[10][17]  ( .CLK(n3481), .D(n3354), .Q(
        \inq_ary[10][17] ) );
  LATCHX1_RVT \inq_ary_reg[11][17]  ( .CLK(n3480), .D(n3354), .Q(
        \inq_ary[11][17] ) );
  LATCHX1_RVT \inq_ary_reg[12][17]  ( .CLK(n3479), .D(n3354), .Q(
        \inq_ary[12][17] ) );
  LATCHX1_RVT \inq_ary_reg[13][17]  ( .CLK(n3478), .D(n3354), .Q(
        \inq_ary[13][17] ) );
  LATCHX1_RVT \inq_ary_reg[14][17]  ( .CLK(n3477), .D(n3354), .Q(
        \inq_ary[14][17] ) );
  LATCHX1_RVT \inq_ary_reg[15][17]  ( .CLK(n3476), .D(n3354), .Q(
        \inq_ary[15][17] ) );
  LATCHX1_RVT \dout_reg[17]  ( .CLK(n3492), .D(N278), .Q(dout[17]) );
  LATCHX1_RVT \inq_ary_reg[0][16]  ( .CLK(n3491), .D(n3352), .Q(
        \inq_ary[0][16] ) );
  LATCHX1_RVT \inq_ary_reg[1][16]  ( .CLK(n3490), .D(n3352), .Q(
        \inq_ary[1][16] ) );
  LATCHX1_RVT \inq_ary_reg[2][16]  ( .CLK(n3489), .D(n3352), .Q(
        \inq_ary[2][16] ) );
  LATCHX1_RVT \inq_ary_reg[3][16]  ( .CLK(n3488), .D(n3352), .Q(
        \inq_ary[3][16] ) );
  LATCHX1_RVT \inq_ary_reg[4][16]  ( .CLK(n3487), .D(n3352), .Q(
        \inq_ary[4][16] ) );
  LATCHX1_RVT \inq_ary_reg[5][16]  ( .CLK(n3486), .D(n3352), .Q(
        \inq_ary[5][16] ) );
  LATCHX1_RVT \inq_ary_reg[6][16]  ( .CLK(n3485), .D(n3352), .Q(
        \inq_ary[6][16] ) );
  LATCHX1_RVT \inq_ary_reg[7][16]  ( .CLK(n3484), .D(n3352), .Q(
        \inq_ary[7][16] ) );
  LATCHX1_RVT \inq_ary_reg[8][16]  ( .CLK(n3483), .D(n3352), .Q(
        \inq_ary[8][16] ) );
  LATCHX1_RVT \inq_ary_reg[9][16]  ( .CLK(n3482), .D(n3352), .Q(
        \inq_ary[9][16] ) );
  LATCHX1_RVT \inq_ary_reg[10][16]  ( .CLK(n3481), .D(n3352), .Q(
        \inq_ary[10][16] ) );
  LATCHX1_RVT \inq_ary_reg[11][16]  ( .CLK(n3480), .D(n3352), .Q(
        \inq_ary[11][16] ) );
  LATCHX1_RVT \inq_ary_reg[12][16]  ( .CLK(n3479), .D(n3352), .Q(
        \inq_ary[12][16] ) );
  LATCHX1_RVT \inq_ary_reg[13][16]  ( .CLK(n3478), .D(n3352), .Q(
        \inq_ary[13][16] ) );
  LATCHX1_RVT \inq_ary_reg[14][16]  ( .CLK(n3477), .D(n3352), .Q(
        \inq_ary[14][16] ) );
  LATCHX1_RVT \inq_ary_reg[15][16]  ( .CLK(n3476), .D(n3352), .Q(
        \inq_ary[15][16] ) );
  LATCHX1_RVT \dout_reg[16]  ( .CLK(n3492), .D(N277), .Q(dout[16]) );
  LATCHX1_RVT \inq_ary_reg[0][15]  ( .CLK(n3491), .D(n3349), .Q(
        \inq_ary[0][15] ) );
  LATCHX1_RVT \inq_ary_reg[1][15]  ( .CLK(n3490), .D(n3349), .Q(
        \inq_ary[1][15] ) );
  LATCHX1_RVT \inq_ary_reg[2][15]  ( .CLK(n3489), .D(n3349), .Q(
        \inq_ary[2][15] ) );
  LATCHX1_RVT \inq_ary_reg[3][15]  ( .CLK(n3488), .D(n3349), .Q(
        \inq_ary[3][15] ) );
  LATCHX1_RVT \inq_ary_reg[4][15]  ( .CLK(n3487), .D(n3349), .Q(
        \inq_ary[4][15] ) );
  LATCHX1_RVT \inq_ary_reg[5][15]  ( .CLK(n3486), .D(n3349), .Q(
        \inq_ary[5][15] ) );
  LATCHX1_RVT \inq_ary_reg[6][15]  ( .CLK(n3485), .D(n3349), .Q(
        \inq_ary[6][15] ) );
  LATCHX1_RVT \inq_ary_reg[7][15]  ( .CLK(n3484), .D(n3349), .Q(
        \inq_ary[7][15] ) );
  LATCHX1_RVT \inq_ary_reg[8][15]  ( .CLK(n3483), .D(n3349), .Q(
        \inq_ary[8][15] ) );
  LATCHX1_RVT \inq_ary_reg[9][15]  ( .CLK(n3482), .D(n3349), .Q(
        \inq_ary[9][15] ) );
  LATCHX1_RVT \inq_ary_reg[10][15]  ( .CLK(n3481), .D(n3349), .Q(
        \inq_ary[10][15] ) );
  LATCHX1_RVT \inq_ary_reg[11][15]  ( .CLK(n3480), .D(n3349), .Q(
        \inq_ary[11][15] ) );
  LATCHX1_RVT \inq_ary_reg[12][15]  ( .CLK(n3479), .D(n3349), .Q(
        \inq_ary[12][15] ) );
  LATCHX1_RVT \inq_ary_reg[13][15]  ( .CLK(n3478), .D(n3349), .Q(
        \inq_ary[13][15] ) );
  LATCHX1_RVT \inq_ary_reg[14][15]  ( .CLK(n3477), .D(n3349), .Q(
        \inq_ary[14][15] ) );
  LATCHX1_RVT \inq_ary_reg[15][15]  ( .CLK(n3476), .D(n3349), .Q(
        \inq_ary[15][15] ) );
  LATCHX1_RVT \dout_reg[15]  ( .CLK(n3492), .D(N276), .Q(dout[15]) );
  LATCHX1_RVT \inq_ary_reg[0][14]  ( .CLK(n3491), .D(n3347), .Q(
        \inq_ary[0][14] ) );
  LATCHX1_RVT \inq_ary_reg[1][14]  ( .CLK(n3490), .D(n3347), .Q(
        \inq_ary[1][14] ) );
  LATCHX1_RVT \inq_ary_reg[2][14]  ( .CLK(n3489), .D(n3347), .Q(
        \inq_ary[2][14] ) );
  LATCHX1_RVT \inq_ary_reg[3][14]  ( .CLK(n3488), .D(n3347), .Q(
        \inq_ary[3][14] ) );
  LATCHX1_RVT \inq_ary_reg[4][14]  ( .CLK(n3487), .D(n3347), .Q(
        \inq_ary[4][14] ) );
  LATCHX1_RVT \inq_ary_reg[5][14]  ( .CLK(n3486), .D(n3347), .Q(
        \inq_ary[5][14] ) );
  LATCHX1_RVT \inq_ary_reg[6][14]  ( .CLK(n3485), .D(n3347), .Q(
        \inq_ary[6][14] ) );
  LATCHX1_RVT \inq_ary_reg[7][14]  ( .CLK(n3484), .D(n3347), .Q(
        \inq_ary[7][14] ) );
  LATCHX1_RVT \inq_ary_reg[8][14]  ( .CLK(n3483), .D(n3347), .Q(
        \inq_ary[8][14] ) );
  LATCHX1_RVT \inq_ary_reg[9][14]  ( .CLK(n3482), .D(n3347), .Q(
        \inq_ary[9][14] ) );
  LATCHX1_RVT \inq_ary_reg[10][14]  ( .CLK(n3481), .D(n3347), .Q(
        \inq_ary[10][14] ) );
  LATCHX1_RVT \inq_ary_reg[11][14]  ( .CLK(n3480), .D(n3347), .Q(
        \inq_ary[11][14] ) );
  LATCHX1_RVT \inq_ary_reg[12][14]  ( .CLK(n3479), .D(n3347), .Q(
        \inq_ary[12][14] ) );
  LATCHX1_RVT \inq_ary_reg[13][14]  ( .CLK(n3478), .D(n3347), .Q(
        \inq_ary[13][14] ) );
  LATCHX1_RVT \inq_ary_reg[14][14]  ( .CLK(n3477), .D(n3347), .Q(
        \inq_ary[14][14] ) );
  LATCHX1_RVT \inq_ary_reg[15][14]  ( .CLK(n3476), .D(n3347), .Q(
        \inq_ary[15][14] ) );
  LATCHX1_RVT \dout_reg[14]  ( .CLK(n3492), .D(N275), .Q(dout[14]) );
  LATCHX1_RVT \inq_ary_reg[0][13]  ( .CLK(n3491), .D(n3345), .Q(
        \inq_ary[0][13] ) );
  LATCHX1_RVT \inq_ary_reg[1][13]  ( .CLK(n3490), .D(n3345), .Q(
        \inq_ary[1][13] ) );
  LATCHX1_RVT \inq_ary_reg[2][13]  ( .CLK(n3489), .D(n3345), .Q(
        \inq_ary[2][13] ) );
  LATCHX1_RVT \inq_ary_reg[3][13]  ( .CLK(n3488), .D(n3345), .Q(
        \inq_ary[3][13] ) );
  LATCHX1_RVT \inq_ary_reg[4][13]  ( .CLK(n3487), .D(n3345), .Q(
        \inq_ary[4][13] ) );
  LATCHX1_RVT \inq_ary_reg[5][13]  ( .CLK(n3486), .D(n3345), .Q(
        \inq_ary[5][13] ) );
  LATCHX1_RVT \inq_ary_reg[6][13]  ( .CLK(n3485), .D(n3345), .Q(
        \inq_ary[6][13] ) );
  LATCHX1_RVT \inq_ary_reg[7][13]  ( .CLK(n3484), .D(n3345), .Q(
        \inq_ary[7][13] ) );
  LATCHX1_RVT \inq_ary_reg[8][13]  ( .CLK(n3483), .D(n3345), .Q(
        \inq_ary[8][13] ) );
  LATCHX1_RVT \inq_ary_reg[9][13]  ( .CLK(n3482), .D(n3345), .Q(
        \inq_ary[9][13] ) );
  LATCHX1_RVT \inq_ary_reg[10][13]  ( .CLK(n3481), .D(n3345), .Q(
        \inq_ary[10][13] ) );
  LATCHX1_RVT \inq_ary_reg[11][13]  ( .CLK(n3480), .D(n3345), .Q(
        \inq_ary[11][13] ) );
  LATCHX1_RVT \inq_ary_reg[12][13]  ( .CLK(n3479), .D(n3345), .Q(
        \inq_ary[12][13] ) );
  LATCHX1_RVT \inq_ary_reg[13][13]  ( .CLK(n3478), .D(n3345), .Q(
        \inq_ary[13][13] ) );
  LATCHX1_RVT \inq_ary_reg[14][13]  ( .CLK(n3477), .D(n3345), .Q(
        \inq_ary[14][13] ) );
  LATCHX1_RVT \inq_ary_reg[15][13]  ( .CLK(n3476), .D(n3345), .Q(
        \inq_ary[15][13] ) );
  LATCHX1_RVT \dout_reg[13]  ( .CLK(n3492), .D(N274), .Q(dout[13]) );
  LATCHX1_RVT \inq_ary_reg[0][12]  ( .CLK(n3491), .D(n3343), .Q(
        \inq_ary[0][12] ) );
  LATCHX1_RVT \inq_ary_reg[1][12]  ( .CLK(n3490), .D(n3343), .Q(
        \inq_ary[1][12] ) );
  LATCHX1_RVT \inq_ary_reg[2][12]  ( .CLK(n3489), .D(n3343), .Q(
        \inq_ary[2][12] ) );
  LATCHX1_RVT \inq_ary_reg[3][12]  ( .CLK(n3488), .D(n3343), .Q(
        \inq_ary[3][12] ) );
  LATCHX1_RVT \inq_ary_reg[4][12]  ( .CLK(n3487), .D(n3343), .Q(
        \inq_ary[4][12] ) );
  LATCHX1_RVT \inq_ary_reg[5][12]  ( .CLK(n3486), .D(n3343), .Q(
        \inq_ary[5][12] ) );
  LATCHX1_RVT \inq_ary_reg[6][12]  ( .CLK(n3485), .D(n3343), .Q(
        \inq_ary[6][12] ) );
  LATCHX1_RVT \inq_ary_reg[7][12]  ( .CLK(n3484), .D(n3343), .Q(
        \inq_ary[7][12] ) );
  LATCHX1_RVT \inq_ary_reg[8][12]  ( .CLK(n3483), .D(n3343), .Q(
        \inq_ary[8][12] ) );
  LATCHX1_RVT \inq_ary_reg[9][12]  ( .CLK(n3482), .D(n3343), .Q(
        \inq_ary[9][12] ) );
  LATCHX1_RVT \inq_ary_reg[10][12]  ( .CLK(n3481), .D(n3343), .Q(
        \inq_ary[10][12] ) );
  LATCHX1_RVT \inq_ary_reg[11][12]  ( .CLK(n3480), .D(n3343), .Q(
        \inq_ary[11][12] ) );
  LATCHX1_RVT \inq_ary_reg[12][12]  ( .CLK(n3479), .D(n3343), .Q(
        \inq_ary[12][12] ) );
  LATCHX1_RVT \inq_ary_reg[13][12]  ( .CLK(n3478), .D(n3343), .Q(
        \inq_ary[13][12] ) );
  LATCHX1_RVT \inq_ary_reg[14][12]  ( .CLK(n3477), .D(n3343), .Q(
        \inq_ary[14][12] ) );
  LATCHX1_RVT \inq_ary_reg[15][12]  ( .CLK(n3476), .D(n3343), .Q(
        \inq_ary[15][12] ) );
  LATCHX1_RVT \dout_reg[12]  ( .CLK(n3492), .D(N273), .Q(dout[12]) );
  LATCHX1_RVT \inq_ary_reg[0][11]  ( .CLK(n3491), .D(n3350), .Q(
        \inq_ary[0][11] ) );
  LATCHX1_RVT \inq_ary_reg[1][11]  ( .CLK(n3490), .D(n3350), .Q(
        \inq_ary[1][11] ) );
  LATCHX1_RVT \inq_ary_reg[2][11]  ( .CLK(n3489), .D(n3350), .Q(
        \inq_ary[2][11] ) );
  LATCHX1_RVT \inq_ary_reg[3][11]  ( .CLK(n3488), .D(n3350), .Q(
        \inq_ary[3][11] ) );
  LATCHX1_RVT \inq_ary_reg[4][11]  ( .CLK(n3487), .D(n3350), .Q(
        \inq_ary[4][11] ) );
  LATCHX1_RVT \inq_ary_reg[5][11]  ( .CLK(n3486), .D(n3350), .Q(
        \inq_ary[5][11] ) );
  LATCHX1_RVT \inq_ary_reg[6][11]  ( .CLK(n3485), .D(n3350), .Q(
        \inq_ary[6][11] ) );
  LATCHX1_RVT \inq_ary_reg[7][11]  ( .CLK(n3484), .D(n3350), .Q(
        \inq_ary[7][11] ) );
  LATCHX1_RVT \inq_ary_reg[8][11]  ( .CLK(n3483), .D(n3350), .Q(
        \inq_ary[8][11] ) );
  LATCHX1_RVT \inq_ary_reg[9][11]  ( .CLK(n3482), .D(n3350), .Q(
        \inq_ary[9][11] ) );
  LATCHX1_RVT \inq_ary_reg[10][11]  ( .CLK(n3481), .D(n3350), .Q(
        \inq_ary[10][11] ) );
  LATCHX1_RVT \inq_ary_reg[11][11]  ( .CLK(n3480), .D(n3350), .Q(
        \inq_ary[11][11] ) );
  LATCHX1_RVT \inq_ary_reg[12][11]  ( .CLK(n3479), .D(n3350), .Q(
        \inq_ary[12][11] ) );
  LATCHX1_RVT \inq_ary_reg[13][11]  ( .CLK(n3478), .D(n3350), .Q(
        \inq_ary[13][11] ) );
  LATCHX1_RVT \inq_ary_reg[14][11]  ( .CLK(n3477), .D(n3350), .Q(
        \inq_ary[14][11] ) );
  LATCHX1_RVT \inq_ary_reg[15][11]  ( .CLK(n3476), .D(n3350), .Q(
        \inq_ary[15][11] ) );
  LATCHX1_RVT \dout_reg[11]  ( .CLK(n3492), .D(N272), .Q(dout[11]) );
  LATCHX1_RVT \inq_ary_reg[0][10]  ( .CLK(n3491), .D(n3348), .Q(
        \inq_ary[0][10] ) );
  LATCHX1_RVT \inq_ary_reg[1][10]  ( .CLK(n3490), .D(n3348), .Q(
        \inq_ary[1][10] ) );
  LATCHX1_RVT \inq_ary_reg[2][10]  ( .CLK(n3489), .D(n3348), .Q(
        \inq_ary[2][10] ) );
  LATCHX1_RVT \inq_ary_reg[3][10]  ( .CLK(n3488), .D(n3348), .Q(
        \inq_ary[3][10] ) );
  LATCHX1_RVT \inq_ary_reg[4][10]  ( .CLK(n3487), .D(n3348), .Q(
        \inq_ary[4][10] ) );
  LATCHX1_RVT \inq_ary_reg[5][10]  ( .CLK(n3486), .D(n3348), .Q(
        \inq_ary[5][10] ) );
  LATCHX1_RVT \inq_ary_reg[6][10]  ( .CLK(n3485), .D(n3348), .Q(
        \inq_ary[6][10] ) );
  LATCHX1_RVT \inq_ary_reg[7][10]  ( .CLK(n3484), .D(n3348), .Q(
        \inq_ary[7][10] ) );
  LATCHX1_RVT \inq_ary_reg[8][10]  ( .CLK(n3483), .D(n3348), .Q(
        \inq_ary[8][10] ) );
  LATCHX1_RVT \inq_ary_reg[9][10]  ( .CLK(n3482), .D(n3348), .Q(
        \inq_ary[9][10] ) );
  LATCHX1_RVT \inq_ary_reg[10][10]  ( .CLK(n3481), .D(n3348), .Q(
        \inq_ary[10][10] ) );
  LATCHX1_RVT \inq_ary_reg[11][10]  ( .CLK(n3480), .D(n3348), .Q(
        \inq_ary[11][10] ) );
  LATCHX1_RVT \inq_ary_reg[12][10]  ( .CLK(n3479), .D(n3348), .Q(
        \inq_ary[12][10] ) );
  LATCHX1_RVT \inq_ary_reg[13][10]  ( .CLK(n3478), .D(n3348), .Q(
        \inq_ary[13][10] ) );
  LATCHX1_RVT \inq_ary_reg[14][10]  ( .CLK(n3477), .D(n3348), .Q(
        \inq_ary[14][10] ) );
  LATCHX1_RVT \inq_ary_reg[15][10]  ( .CLK(n3476), .D(n3348), .Q(
        \inq_ary[15][10] ) );
  LATCHX1_RVT \dout_reg[10]  ( .CLK(n3492), .D(N271), .Q(dout[10]) );
  LATCHX1_RVT \inq_ary_reg[0][9]  ( .CLK(n3491), .D(n3346), .Q(\inq_ary[0][9] ) );
  LATCHX1_RVT \inq_ary_reg[1][9]  ( .CLK(n3490), .D(n3346), .Q(\inq_ary[1][9] ) );
  LATCHX1_RVT \inq_ary_reg[2][9]  ( .CLK(n3489), .D(n3346), .Q(\inq_ary[2][9] ) );
  LATCHX1_RVT \inq_ary_reg[3][9]  ( .CLK(n3488), .D(n3346), .Q(\inq_ary[3][9] ) );
  LATCHX1_RVT \inq_ary_reg[4][9]  ( .CLK(n3487), .D(n3346), .Q(\inq_ary[4][9] ) );
  LATCHX1_RVT \inq_ary_reg[5][9]  ( .CLK(n3486), .D(n3346), .Q(\inq_ary[5][9] ) );
  LATCHX1_RVT \inq_ary_reg[6][9]  ( .CLK(n3485), .D(n3346), .Q(\inq_ary[6][9] ) );
  LATCHX1_RVT \inq_ary_reg[7][9]  ( .CLK(n3484), .D(n3346), .Q(\inq_ary[7][9] ) );
  LATCHX1_RVT \inq_ary_reg[8][9]  ( .CLK(n3483), .D(n3346), .Q(\inq_ary[8][9] ) );
  LATCHX1_RVT \inq_ary_reg[9][9]  ( .CLK(n3482), .D(n3346), .Q(\inq_ary[9][9] ) );
  LATCHX1_RVT \inq_ary_reg[10][9]  ( .CLK(n3481), .D(n3346), .Q(
        \inq_ary[10][9] ) );
  LATCHX1_RVT \inq_ary_reg[11][9]  ( .CLK(n3480), .D(n3346), .Q(
        \inq_ary[11][9] ) );
  LATCHX1_RVT \inq_ary_reg[12][9]  ( .CLK(n3479), .D(n3346), .Q(
        \inq_ary[12][9] ) );
  LATCHX1_RVT \inq_ary_reg[13][9]  ( .CLK(n3478), .D(n3346), .Q(
        \inq_ary[13][9] ) );
  LATCHX1_RVT \inq_ary_reg[14][9]  ( .CLK(n3477), .D(n3346), .Q(
        \inq_ary[14][9] ) );
  LATCHX1_RVT \inq_ary_reg[15][9]  ( .CLK(n3476), .D(n3346), .Q(
        \inq_ary[15][9] ) );
  LATCHX1_RVT \dout_reg[9]  ( .CLK(n3492), .D(N270), .Q(dout[9]) );
  LATCHX1_RVT \inq_ary_reg[0][8]  ( .CLK(n3491), .D(n3344), .Q(\inq_ary[0][8] ) );
  LATCHX1_RVT \inq_ary_reg[1][8]  ( .CLK(n3490), .D(n3344), .Q(\inq_ary[1][8] ) );
  LATCHX1_RVT \inq_ary_reg[2][8]  ( .CLK(n3489), .D(n3344), .Q(\inq_ary[2][8] ) );
  LATCHX1_RVT \inq_ary_reg[3][8]  ( .CLK(n3488), .D(n3344), .Q(\inq_ary[3][8] ) );
  LATCHX1_RVT \inq_ary_reg[4][8]  ( .CLK(n3487), .D(n3344), .Q(\inq_ary[4][8] ) );
  LATCHX1_RVT \inq_ary_reg[5][8]  ( .CLK(n3486), .D(n3344), .Q(\inq_ary[5][8] ) );
  LATCHX1_RVT \inq_ary_reg[6][8]  ( .CLK(n3485), .D(n3344), .Q(\inq_ary[6][8] ) );
  LATCHX1_RVT \inq_ary_reg[7][8]  ( .CLK(n3484), .D(n3344), .Q(\inq_ary[7][8] ) );
  LATCHX1_RVT \inq_ary_reg[8][8]  ( .CLK(n3483), .D(n3344), .Q(\inq_ary[8][8] ) );
  LATCHX1_RVT \inq_ary_reg[9][8]  ( .CLK(n3482), .D(n3344), .Q(\inq_ary[9][8] ) );
  LATCHX1_RVT \inq_ary_reg[10][8]  ( .CLK(n3481), .D(n3344), .Q(
        \inq_ary[10][8] ) );
  LATCHX1_RVT \inq_ary_reg[11][8]  ( .CLK(n3480), .D(n3344), .Q(
        \inq_ary[11][8] ) );
  LATCHX1_RVT \inq_ary_reg[12][8]  ( .CLK(n3479), .D(n3344), .Q(
        \inq_ary[12][8] ) );
  LATCHX1_RVT \inq_ary_reg[13][8]  ( .CLK(n3478), .D(n3344), .Q(
        \inq_ary[13][8] ) );
  LATCHX1_RVT \inq_ary_reg[14][8]  ( .CLK(n3477), .D(n3344), .Q(
        \inq_ary[14][8] ) );
  LATCHX1_RVT \inq_ary_reg[15][8]  ( .CLK(n3476), .D(n3344), .Q(
        \inq_ary[15][8] ) );
  LATCHX1_RVT \dout_reg[8]  ( .CLK(n3492), .D(N269), .Q(dout[8]) );
  LATCHX1_RVT \inq_ary_reg[0][7]  ( .CLK(n3491), .D(n3342), .Q(\inq_ary[0][7] ) );
  LATCHX1_RVT \inq_ary_reg[1][7]  ( .CLK(n3490), .D(n3342), .Q(\inq_ary[1][7] ) );
  LATCHX1_RVT \inq_ary_reg[2][7]  ( .CLK(n3489), .D(n3342), .Q(\inq_ary[2][7] ) );
  LATCHX1_RVT \inq_ary_reg[3][7]  ( .CLK(n3488), .D(n3342), .Q(\inq_ary[3][7] ) );
  LATCHX1_RVT \inq_ary_reg[4][7]  ( .CLK(n3487), .D(n3342), .Q(\inq_ary[4][7] ) );
  LATCHX1_RVT \inq_ary_reg[5][7]  ( .CLK(n3486), .D(n3342), .Q(\inq_ary[5][7] ) );
  LATCHX1_RVT \inq_ary_reg[6][7]  ( .CLK(n3485), .D(n3342), .Q(\inq_ary[6][7] ) );
  LATCHX1_RVT \inq_ary_reg[7][7]  ( .CLK(n3484), .D(n3342), .Q(\inq_ary[7][7] ) );
  LATCHX1_RVT \inq_ary_reg[8][7]  ( .CLK(n3483), .D(n3342), .Q(\inq_ary[8][7] ) );
  LATCHX1_RVT \inq_ary_reg[9][7]  ( .CLK(n3482), .D(n3342), .Q(\inq_ary[9][7] ) );
  LATCHX1_RVT \inq_ary_reg[10][7]  ( .CLK(n3481), .D(n3342), .Q(
        \inq_ary[10][7] ) );
  LATCHX1_RVT \inq_ary_reg[11][7]  ( .CLK(n3480), .D(n3342), .Q(
        \inq_ary[11][7] ) );
  LATCHX1_RVT \inq_ary_reg[12][7]  ( .CLK(n3479), .D(n3342), .Q(
        \inq_ary[12][7] ) );
  LATCHX1_RVT \inq_ary_reg[13][7]  ( .CLK(n3478), .D(n3342), .Q(
        \inq_ary[13][7] ) );
  LATCHX1_RVT \inq_ary_reg[14][7]  ( .CLK(n3477), .D(n3342), .Q(
        \inq_ary[14][7] ) );
  LATCHX1_RVT \inq_ary_reg[15][7]  ( .CLK(n3476), .D(n3342), .Q(
        \inq_ary[15][7] ) );
  LATCHX1_RVT \dout_reg[7]  ( .CLK(n3492), .D(N268), .Q(dout[7]) );
  LATCHX1_RVT \inq_ary_reg[0][6]  ( .CLK(n3491), .D(n3341), .Q(\inq_ary[0][6] ) );
  LATCHX1_RVT \inq_ary_reg[1][6]  ( .CLK(n3490), .D(n3341), .Q(\inq_ary[1][6] ) );
  LATCHX1_RVT \inq_ary_reg[2][6]  ( .CLK(n3489), .D(n3341), .Q(\inq_ary[2][6] ) );
  LATCHX1_RVT \inq_ary_reg[3][6]  ( .CLK(n3488), .D(n3341), .Q(\inq_ary[3][6] ) );
  LATCHX1_RVT \inq_ary_reg[4][6]  ( .CLK(n3487), .D(n3341), .Q(\inq_ary[4][6] ) );
  LATCHX1_RVT \inq_ary_reg[5][6]  ( .CLK(n3486), .D(n3341), .Q(\inq_ary[5][6] ) );
  LATCHX1_RVT \inq_ary_reg[6][6]  ( .CLK(n3485), .D(n3341), .Q(\inq_ary[6][6] ) );
  LATCHX1_RVT \inq_ary_reg[7][6]  ( .CLK(n3484), .D(n3341), .Q(\inq_ary[7][6] ) );
  LATCHX1_RVT \inq_ary_reg[8][6]  ( .CLK(n3483), .D(n3341), .Q(\inq_ary[8][6] ) );
  LATCHX1_RVT \inq_ary_reg[9][6]  ( .CLK(n3482), .D(n3341), .Q(\inq_ary[9][6] ) );
  LATCHX1_RVT \inq_ary_reg[10][6]  ( .CLK(n3481), .D(n3341), .Q(
        \inq_ary[10][6] ) );
  LATCHX1_RVT \inq_ary_reg[11][6]  ( .CLK(n3480), .D(n3341), .Q(
        \inq_ary[11][6] ) );
  LATCHX1_RVT \inq_ary_reg[12][6]  ( .CLK(n3479), .D(n3341), .Q(
        \inq_ary[12][6] ) );
  LATCHX1_RVT \inq_ary_reg[13][6]  ( .CLK(n3478), .D(n3341), .Q(
        \inq_ary[13][6] ) );
  LATCHX1_RVT \inq_ary_reg[14][6]  ( .CLK(n3477), .D(n3341), .Q(
        \inq_ary[14][6] ) );
  LATCHX1_RVT \inq_ary_reg[15][6]  ( .CLK(n3476), .D(n3341), .Q(
        \inq_ary[15][6] ) );
  LATCHX1_RVT \dout_reg[6]  ( .CLK(n3492), .D(N267), .Q(dout[6]) );
  LATCHX1_RVT \inq_ary_reg[0][5]  ( .CLK(n3491), .D(n3340), .Q(\inq_ary[0][5] ) );
  LATCHX1_RVT \inq_ary_reg[1][5]  ( .CLK(n3490), .D(n3340), .Q(\inq_ary[1][5] ) );
  LATCHX1_RVT \inq_ary_reg[2][5]  ( .CLK(n3489), .D(n3340), .Q(\inq_ary[2][5] ) );
  LATCHX1_RVT \inq_ary_reg[3][5]  ( .CLK(n3488), .D(n3340), .Q(\inq_ary[3][5] ) );
  LATCHX1_RVT \inq_ary_reg[4][5]  ( .CLK(n3487), .D(n3340), .Q(\inq_ary[4][5] ) );
  LATCHX1_RVT \inq_ary_reg[5][5]  ( .CLK(n3486), .D(n3340), .Q(\inq_ary[5][5] ) );
  LATCHX1_RVT \inq_ary_reg[6][5]  ( .CLK(n3485), .D(n3340), .Q(\inq_ary[6][5] ) );
  LATCHX1_RVT \inq_ary_reg[7][5]  ( .CLK(n3484), .D(n3340), .Q(\inq_ary[7][5] ) );
  LATCHX1_RVT \inq_ary_reg[8][5]  ( .CLK(n3483), .D(n3340), .Q(\inq_ary[8][5] ) );
  LATCHX1_RVT \inq_ary_reg[9][5]  ( .CLK(n3482), .D(n3340), .Q(\inq_ary[9][5] ) );
  LATCHX1_RVT \inq_ary_reg[10][5]  ( .CLK(n3481), .D(n3340), .Q(
        \inq_ary[10][5] ) );
  LATCHX1_RVT \inq_ary_reg[11][5]  ( .CLK(n3480), .D(n3340), .Q(
        \inq_ary[11][5] ) );
  LATCHX1_RVT \inq_ary_reg[12][5]  ( .CLK(n3479), .D(n3340), .Q(
        \inq_ary[12][5] ) );
  LATCHX1_RVT \inq_ary_reg[13][5]  ( .CLK(n3478), .D(n3340), .Q(
        \inq_ary[13][5] ) );
  LATCHX1_RVT \inq_ary_reg[14][5]  ( .CLK(n3477), .D(n3340), .Q(
        \inq_ary[14][5] ) );
  LATCHX1_RVT \inq_ary_reg[15][5]  ( .CLK(n3476), .D(n3340), .Q(
        \inq_ary[15][5] ) );
  LATCHX1_RVT \dout_reg[5]  ( .CLK(n3492), .D(N266), .Q(dout[5]) );
  DFFX1_RVT \rdptr_d1_reg[1]  ( .D(rd_adr[1]), .CLK(net24660), .Q(rdptr_d1[1]), 
        .QN(n3337) );
  DFFX1_RVT \wrptr_d1_reg[2]  ( .D(wr_adr[2]), .CLK(net24660), .Q(wrptr_d1[2]), 
        .QN(n3336) );
  DFFX1_RVT \wrptr_d1_reg[3]  ( .D(wr_adr[3]), .CLK(net24660), .Q(wrptr_d1[3]), 
        .QN(n3335) );
  DFFX1_RVT \rdptr_d1_reg[0]  ( .D(rd_adr[0]), .CLK(net24660), .Q(rdptr_d1[0]), 
        .QN(n3334) );
  DFFX1_RVT \wrptr_d1_reg[1]  ( .D(wr_adr[1]), .CLK(net24660), .Q(wrptr_d1[1]), 
        .QN(n6) );
  DFFX1_RVT \rdptr_d1_reg[3]  ( .D(rd_adr[3]), .CLK(net24660), .Q(rdptr_d1[3]), 
        .QN(n5) );
  DFFX1_RVT \wrptr_d1_reg[0]  ( .D(wr_adr[0]), .CLK(net24660), .Q(wrptr_d1[0]), 
        .QN(n4) );
  DFFSSRX1_RVT ren_d1_reg ( .D(1'b0), .SETB(1'b0), .RSTB(read_en), .CLK(
        net24660), .QN(n3339) );
  INVX1_RVT U3 ( .A(n1760), .Y(n1) );
  INVX1_RVT U4 ( .A(n1598), .Y(n2) );
  NAND2X1_RVT U5 ( .A1(n3339), .A2(reset_l), .Y(n3492) );
  INVX1_RVT U6 ( .A(n946), .Y(n3) );
  INVX1_RVT U8 ( .A(rst_tri_en), .Y(n7) );
  NAND2X0_RVT U9 ( .A1(wr_en_d1), .A2(n7), .Y(n946) );
  INVX1_RVT U10 ( .A(n946), .Y(n758) );
  INVX1_RVT U11 ( .A(n946), .Y(n1598) );
  INVX1_RVT U12 ( .A(n1598), .Y(n969) );
  AND4X1_RVT U13 ( .A1(wrptr_d1[0]), .A2(wrptr_d1[1]), .A3(n3335), .A4(n3336), 
        .Y(n1742) );
  AND4X1_RVT U14 ( .A1(n4), .A2(n3335), .A3(n6), .A4(n3336), .Y(n1686) );
  AO22X1_RVT U15 ( .A1(n1742), .A2(\inq_ary[3][96] ), .A3(n1686), .A4(
        \inq_ary[0][96] ), .Y(n11) );
  AND4X1_RVT U16 ( .A1(wrptr_d1[0]), .A2(wrptr_d1[3]), .A3(wrptr_d1[1]), .A4(
        wrptr_d1[2]), .Y(n1537) );
  AND2X1_RVT U17 ( .A1(n4), .A2(n3335), .Y(n13) );
  AND3X1_RVT U18 ( .A1(n13), .A2(wrptr_d1[1]), .A3(wrptr_d1[2]), .Y(n1738) );
  AO22X1_RVT U19 ( .A1(n1537), .A2(\inq_ary[15][96] ), .A3(n1738), .A4(
        \inq_ary[6][96] ), .Y(n10) );
  AND4X1_RVT U20 ( .A1(wrptr_d1[3]), .A2(wrptr_d1[1]), .A3(n4), .A4(n3336), 
        .Y(n1748) );
  AND2X1_RVT U21 ( .A1(n6), .A2(n3336), .Y(n12) );
  AND3X1_RVT U22 ( .A1(wrptr_d1[0]), .A2(wrptr_d1[3]), .A3(n12), .Y(n1751) );
  AO22X1_RVT U23 ( .A1(n1748), .A2(\inq_ary[10][96] ), .A3(n1751), .A4(
        \inq_ary[9][96] ), .Y(n9) );
  AND4X1_RVT U24 ( .A1(wrptr_d1[0]), .A2(wrptr_d1[2]), .A3(n6), .A4(n3335), 
        .Y(n1747) );
  AND4X1_RVT U25 ( .A1(wrptr_d1[3]), .A2(wrptr_d1[0]), .A3(wrptr_d1[2]), .A4(
        n6), .Y(n1711) );
  AO22X1_RVT U26 ( .A1(n1747), .A2(\inq_ary[5][96] ), .A3(n1711), .A4(
        \inq_ary[13][96] ), .Y(n8) );
  NOR4X1_RVT U27 ( .A1(n11), .A2(n10), .A3(n9), .A4(n8), .Y(n19) );
  AND4X1_RVT U28 ( .A1(wrptr_d1[3]), .A2(wrptr_d1[2]), .A3(n4), .A4(n6), .Y(
        n1740) );
  AND3X1_RVT U29 ( .A1(wrptr_d1[0]), .A2(n12), .A3(n3335), .Y(n1749) );
  AO22X1_RVT U30 ( .A1(n1740), .A2(\inq_ary[12][96] ), .A3(n1749), .A4(
        \inq_ary[1][96] ), .Y(n17) );
  AND4X1_RVT U31 ( .A1(wrptr_d1[3]), .A2(wrptr_d1[1]), .A3(wrptr_d1[2]), .A4(
        n4), .Y(n1554) );
  AND4X1_RVT U32 ( .A1(wrptr_d1[3]), .A2(wrptr_d1[0]), .A3(wrptr_d1[1]), .A4(
        n3336), .Y(n1750) );
  AO22X1_RVT U33 ( .A1(n1554), .A2(\inq_ary[14][96] ), .A3(n1750), .A4(
        \inq_ary[11][96] ), .Y(n16) );
  AND3X1_RVT U34 ( .A1(wrptr_d1[3]), .A2(n12), .A3(n4), .Y(n1612) );
  AND4X1_RVT U35 ( .A1(wrptr_d1[0]), .A2(wrptr_d1[1]), .A3(wrptr_d1[2]), .A4(
        n3335), .Y(n1741) );
  AO22X1_RVT U36 ( .A1(n1612), .A2(\inq_ary[8][96] ), .A3(n1741), .A4(
        \inq_ary[7][96] ), .Y(n15) );
  AND3X1_RVT U37 ( .A1(wrptr_d1[1]), .A2(n13), .A3(n3336), .Y(n1739) );
  AND3X1_RVT U38 ( .A1(n13), .A2(wrptr_d1[2]), .A3(n6), .Y(n1729) );
  AO22X1_RVT U39 ( .A1(n1739), .A2(\inq_ary[2][96] ), .A3(n1729), .A4(
        \inq_ary[4][96] ), .Y(n14) );
  NOR4X1_RVT U40 ( .A1(n17), .A2(n16), .A3(n15), .A4(n14), .Y(n18) );
  NAND2X0_RVT U41 ( .A1(n19), .A2(n18), .Y(n20) );
  AO22X1_RVT U42 ( .A1(n758), .A2(wrdata_d1[96]), .A3(n969), .A4(n20), .Y(
        n3425) );
  AO22X1_RVT U43 ( .A1(n1749), .A2(\inq_ary[1][97] ), .A3(n1747), .A4(
        \inq_ary[5][97] ), .Y(n24) );
  AO22X1_RVT U44 ( .A1(n1554), .A2(\inq_ary[14][97] ), .A3(n1537), .A4(
        \inq_ary[15][97] ), .Y(n23) );
  AO22X1_RVT U45 ( .A1(n1729), .A2(\inq_ary[4][97] ), .A3(n1740), .A4(
        \inq_ary[12][97] ), .Y(n22) );
  AO22X1_RVT U46 ( .A1(n1612), .A2(\inq_ary[8][97] ), .A3(n1750), .A4(
        \inq_ary[11][97] ), .Y(n21) );
  NOR4X1_RVT U47 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .Y(n30) );
  AO22X1_RVT U48 ( .A1(n1742), .A2(\inq_ary[3][97] ), .A3(n1738), .A4(
        \inq_ary[6][97] ), .Y(n28) );
  AO22X1_RVT U49 ( .A1(n1711), .A2(\inq_ary[13][97] ), .A3(n1751), .A4(
        \inq_ary[9][97] ), .Y(n27) );
  AO22X1_RVT U50 ( .A1(n1739), .A2(\inq_ary[2][97] ), .A3(n1686), .A4(
        \inq_ary[0][97] ), .Y(n26) );
  AO22X1_RVT U51 ( .A1(n1741), .A2(\inq_ary[7][97] ), .A3(n1748), .A4(
        \inq_ary[10][97] ), .Y(n25) );
  NOR4X1_RVT U52 ( .A1(n28), .A2(n27), .A3(n26), .A4(n25), .Y(n29) );
  NAND2X0_RVT U53 ( .A1(n30), .A2(n29), .Y(n31) );
  AO22X1_RVT U54 ( .A1(n758), .A2(wrdata_d1[97]), .A3(n1), .A4(n31), .Y(n3427)
         );
  AO22X1_RVT U55 ( .A1(n1612), .A2(\inq_ary[8][41] ), .A3(n1738), .A4(
        \inq_ary[6][41] ), .Y(n35) );
  AO22X1_RVT U56 ( .A1(n1741), .A2(\inq_ary[7][41] ), .A3(n1748), .A4(
        \inq_ary[10][41] ), .Y(n34) );
  AO22X1_RVT U57 ( .A1(n1749), .A2(\inq_ary[1][41] ), .A3(n1751), .A4(
        \inq_ary[9][41] ), .Y(n33) );
  AO22X1_RVT U58 ( .A1(n1740), .A2(\inq_ary[12][41] ), .A3(n1747), .A4(
        \inq_ary[5][41] ), .Y(n32) );
  NOR4X1_RVT U59 ( .A1(n35), .A2(n34), .A3(n33), .A4(n32), .Y(n41) );
  AO22X1_RVT U60 ( .A1(n1739), .A2(\inq_ary[2][41] ), .A3(n1742), .A4(
        \inq_ary[3][41] ), .Y(n39) );
  AO22X1_RVT U61 ( .A1(n1686), .A2(\inq_ary[0][41] ), .A3(n1711), .A4(
        \inq_ary[13][41] ), .Y(n38) );
  AO22X1_RVT U62 ( .A1(n1729), .A2(\inq_ary[4][41] ), .A3(n1537), .A4(
        \inq_ary[15][41] ), .Y(n37) );
  AO22X1_RVT U63 ( .A1(n1554), .A2(\inq_ary[14][41] ), .A3(n1750), .A4(
        \inq_ary[11][41] ), .Y(n36) );
  NOR4X1_RVT U64 ( .A1(n39), .A2(n38), .A3(n37), .A4(n36), .Y(n40) );
  NAND2X0_RVT U65 ( .A1(n41), .A2(n40), .Y(n42) );
  AO22X1_RVT U66 ( .A1(n1598), .A2(wrdata_d1[41]), .A3(n2), .A4(n42), .Y(n3378) );
  INVX1_RVT U67 ( .A(n946), .Y(n1760) );
  AO22X1_RVT U68 ( .A1(n1537), .A2(\inq_ary[15][98] ), .A3(n1612), .A4(
        \inq_ary[8][98] ), .Y(n46) );
  AO22X1_RVT U69 ( .A1(n1554), .A2(\inq_ary[14][98] ), .A3(n1750), .A4(
        \inq_ary[11][98] ), .Y(n45) );
  AO22X1_RVT U70 ( .A1(n1740), .A2(\inq_ary[12][98] ), .A3(n1738), .A4(
        \inq_ary[6][98] ), .Y(n44) );
  AO22X1_RVT U71 ( .A1(n1729), .A2(\inq_ary[4][98] ), .A3(n1751), .A4(
        \inq_ary[9][98] ), .Y(n43) );
  NOR4X1_RVT U72 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .Y(n52) );
  AO22X1_RVT U73 ( .A1(n1747), .A2(\inq_ary[5][98] ), .A3(n1711), .A4(
        \inq_ary[13][98] ), .Y(n50) );
  AO22X1_RVT U74 ( .A1(n1686), .A2(\inq_ary[0][98] ), .A3(n1749), .A4(
        \inq_ary[1][98] ), .Y(n49) );
  AO22X1_RVT U75 ( .A1(n1741), .A2(\inq_ary[7][98] ), .A3(n1748), .A4(
        \inq_ary[10][98] ), .Y(n48) );
  AO22X1_RVT U76 ( .A1(n1739), .A2(\inq_ary[2][98] ), .A3(n1742), .A4(
        \inq_ary[3][98] ), .Y(n47) );
  NOR4X1_RVT U77 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .Y(n51) );
  NAND2X0_RVT U78 ( .A1(n52), .A2(n51), .Y(n53) );
  AO22X1_RVT U79 ( .A1(n758), .A2(wrdata_d1[98]), .A3(n1), .A4(n53), .Y(n3429)
         );
  AO22X1_RVT U80 ( .A1(n1554), .A2(\inq_ary[14][99] ), .A3(n1711), .A4(
        \inq_ary[13][99] ), .Y(n57) );
  AO22X1_RVT U81 ( .A1(n1740), .A2(\inq_ary[12][99] ), .A3(n1741), .A4(
        \inq_ary[7][99] ), .Y(n56) );
  AO22X1_RVT U82 ( .A1(n1742), .A2(\inq_ary[3][99] ), .A3(n1686), .A4(
        \inq_ary[0][99] ), .Y(n55) );
  AO22X1_RVT U83 ( .A1(n1739), .A2(\inq_ary[2][99] ), .A3(n1729), .A4(
        \inq_ary[4][99] ), .Y(n54) );
  NOR4X1_RVT U84 ( .A1(n57), .A2(n56), .A3(n55), .A4(n54), .Y(n63) );
  AO22X1_RVT U85 ( .A1(n1749), .A2(\inq_ary[1][99] ), .A3(n1751), .A4(
        \inq_ary[9][99] ), .Y(n61) );
  AO22X1_RVT U86 ( .A1(n1537), .A2(\inq_ary[15][99] ), .A3(n1747), .A4(
        \inq_ary[5][99] ), .Y(n60) );
  AO22X1_RVT U87 ( .A1(n1750), .A2(\inq_ary[11][99] ), .A3(n1748), .A4(
        \inq_ary[10][99] ), .Y(n59) );
  AO22X1_RVT U88 ( .A1(n1612), .A2(\inq_ary[8][99] ), .A3(n1738), .A4(
        \inq_ary[6][99] ), .Y(n58) );
  NOR4X1_RVT U89 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .Y(n62) );
  NAND2X0_RVT U90 ( .A1(n63), .A2(n62), .Y(n64) );
  AO22X1_RVT U91 ( .A1(n1684), .A2(wrdata_d1[99]), .A3(n1), .A4(n64), .Y(n3431) );
  AO22X1_RVT U92 ( .A1(n1537), .A2(\inq_ary[15][40] ), .A3(n1751), .A4(
        \inq_ary[9][40] ), .Y(n68) );
  AO22X1_RVT U93 ( .A1(n1686), .A2(\inq_ary[0][40] ), .A3(n1738), .A4(
        \inq_ary[6][40] ), .Y(n67) );
  AO22X1_RVT U94 ( .A1(n1739), .A2(\inq_ary[2][40] ), .A3(n1747), .A4(
        \inq_ary[5][40] ), .Y(n66) );
  AO22X1_RVT U95 ( .A1(n1749), .A2(\inq_ary[1][40] ), .A3(n1748), .A4(
        \inq_ary[10][40] ), .Y(n65) );
  NOR4X1_RVT U96 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .Y(n74) );
  AO22X1_RVT U97 ( .A1(n1729), .A2(\inq_ary[4][40] ), .A3(n1612), .A4(
        \inq_ary[8][40] ), .Y(n72) );
  AO22X1_RVT U98 ( .A1(n1740), .A2(\inq_ary[12][40] ), .A3(n1741), .A4(
        \inq_ary[7][40] ), .Y(n71) );
  AO22X1_RVT U99 ( .A1(n1554), .A2(\inq_ary[14][40] ), .A3(n1742), .A4(
        \inq_ary[3][40] ), .Y(n70) );
  AO22X1_RVT U100 ( .A1(n1750), .A2(\inq_ary[11][40] ), .A3(n1711), .A4(
        \inq_ary[13][40] ), .Y(n69) );
  NOR4X1_RVT U101 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .Y(n73) );
  NAND2X0_RVT U102 ( .A1(n74), .A2(n73), .Y(n75) );
  AO22X1_RVT U103 ( .A1(n1598), .A2(wrdata_d1[40]), .A3(n969), .A4(n75), .Y(
        n3376) );
  AO22X1_RVT U104 ( .A1(n1686), .A2(\inq_ary[0][100] ), .A3(n1751), .A4(
        \inq_ary[9][100] ), .Y(n79) );
  AO22X1_RVT U105 ( .A1(n1554), .A2(\inq_ary[14][100] ), .A3(n1748), .A4(
        \inq_ary[10][100] ), .Y(n78) );
  AO22X1_RVT U106 ( .A1(n1537), .A2(\inq_ary[15][100] ), .A3(n1741), .A4(
        \inq_ary[7][100] ), .Y(n77) );
  AO22X1_RVT U107 ( .A1(n1739), .A2(\inq_ary[2][100] ), .A3(n1711), .A4(
        \inq_ary[13][100] ), .Y(n76) );
  NOR4X1_RVT U108 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .Y(n85) );
  AO22X1_RVT U109 ( .A1(n1612), .A2(\inq_ary[8][100] ), .A3(n1749), .A4(
        \inq_ary[1][100] ), .Y(n83) );
  AO22X1_RVT U110 ( .A1(n1742), .A2(\inq_ary[3][100] ), .A3(n1740), .A4(
        \inq_ary[12][100] ), .Y(n82) );
  AO22X1_RVT U111 ( .A1(n1747), .A2(\inq_ary[5][100] ), .A3(n1738), .A4(
        \inq_ary[6][100] ), .Y(n81) );
  AO22X1_RVT U112 ( .A1(n1729), .A2(\inq_ary[4][100] ), .A3(n1750), .A4(
        \inq_ary[11][100] ), .Y(n80) );
  NOR4X1_RVT U113 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .Y(n84) );
  NAND2X0_RVT U114 ( .A1(n85), .A2(n84), .Y(n86) );
  AO22X1_RVT U115 ( .A1(n758), .A2(wrdata_d1[100]), .A3(n1759), .A4(n86), .Y(
        n3424) );
  AO22X1_RVT U116 ( .A1(n1537), .A2(\inq_ary[15][101] ), .A3(n1749), .A4(
        \inq_ary[1][101] ), .Y(n90) );
  AO22X1_RVT U117 ( .A1(n1729), .A2(\inq_ary[4][101] ), .A3(n1738), .A4(
        \inq_ary[6][101] ), .Y(n89) );
  AO22X1_RVT U118 ( .A1(n1686), .A2(\inq_ary[0][101] ), .A3(n1612), .A4(
        \inq_ary[8][101] ), .Y(n88) );
  AO22X1_RVT U119 ( .A1(n1741), .A2(\inq_ary[7][101] ), .A3(n1751), .A4(
        \inq_ary[9][101] ), .Y(n87) );
  NOR4X1_RVT U120 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .Y(n96) );
  AO22X1_RVT U121 ( .A1(n1739), .A2(\inq_ary[2][101] ), .A3(n1740), .A4(
        \inq_ary[12][101] ), .Y(n94) );
  AO22X1_RVT U122 ( .A1(n1750), .A2(\inq_ary[11][101] ), .A3(n1748), .A4(
        \inq_ary[10][101] ), .Y(n93) );
  AO22X1_RVT U123 ( .A1(n1742), .A2(\inq_ary[3][101] ), .A3(n1747), .A4(
        \inq_ary[5][101] ), .Y(n92) );
  AO22X1_RVT U124 ( .A1(n1554), .A2(\inq_ary[14][101] ), .A3(n1711), .A4(
        \inq_ary[13][101] ), .Y(n91) );
  NOR4X1_RVT U125 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .Y(n95) );
  NAND2X0_RVT U126 ( .A1(n96), .A2(n95), .Y(n97) );
  AO22X1_RVT U127 ( .A1(n758), .A2(wrdata_d1[101]), .A3(n2), .A4(n97), .Y(
        n3426) );
  AO22X1_RVT U128 ( .A1(n1741), .A2(\inq_ary[7][39] ), .A3(n1711), .A4(
        \inq_ary[13][39] ), .Y(n101) );
  AO22X1_RVT U129 ( .A1(n1739), .A2(\inq_ary[2][39] ), .A3(n1747), .A4(
        \inq_ary[5][39] ), .Y(n100) );
  AO22X1_RVT U130 ( .A1(n1686), .A2(\inq_ary[0][39] ), .A3(n1748), .A4(
        \inq_ary[10][39] ), .Y(n99) );
  AO22X1_RVT U131 ( .A1(n1612), .A2(\inq_ary[8][39] ), .A3(n1751), .A4(
        \inq_ary[9][39] ), .Y(n98) );
  NOR4X1_RVT U132 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .Y(n107) );
  AO22X1_RVT U133 ( .A1(n1554), .A2(\inq_ary[14][39] ), .A3(n1742), .A4(
        \inq_ary[3][39] ), .Y(n105) );
  AO22X1_RVT U134 ( .A1(n1729), .A2(\inq_ary[4][39] ), .A3(n1749), .A4(
        \inq_ary[1][39] ), .Y(n104) );
  AO22X1_RVT U135 ( .A1(n1537), .A2(\inq_ary[15][39] ), .A3(n1738), .A4(
        \inq_ary[6][39] ), .Y(n103) );
  AO22X1_RVT U136 ( .A1(n1740), .A2(\inq_ary[12][39] ), .A3(n1750), .A4(
        \inq_ary[11][39] ), .Y(n102) );
  NOR4X1_RVT U137 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .Y(n106) );
  NAND2X0_RVT U138 ( .A1(n107), .A2(n106), .Y(n108) );
  AO22X1_RVT U139 ( .A1(n3), .A2(wrdata_d1[39]), .A3(n2), .A4(n108), .Y(n3373)
         );
  AO22X1_RVT U140 ( .A1(n1741), .A2(\inq_ary[7][89] ), .A3(n1748), .A4(
        \inq_ary[10][89] ), .Y(n112) );
  AO22X1_RVT U141 ( .A1(n1749), .A2(\inq_ary[1][89] ), .A3(n1711), .A4(
        \inq_ary[13][89] ), .Y(n111) );
  AO22X1_RVT U142 ( .A1(n1739), .A2(\inq_ary[2][89] ), .A3(n1750), .A4(
        \inq_ary[11][89] ), .Y(n110) );
  AO22X1_RVT U143 ( .A1(n1537), .A2(\inq_ary[15][89] ), .A3(n1738), .A4(
        \inq_ary[6][89] ), .Y(n109) );
  NOR4X1_RVT U144 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .Y(n118) );
  AO22X1_RVT U145 ( .A1(n1686), .A2(\inq_ary[0][89] ), .A3(n1612), .A4(
        \inq_ary[8][89] ), .Y(n116) );
  AO22X1_RVT U146 ( .A1(n1554), .A2(\inq_ary[14][89] ), .A3(n1747), .A4(
        \inq_ary[5][89] ), .Y(n115) );
  AO22X1_RVT U147 ( .A1(n1729), .A2(\inq_ary[4][89] ), .A3(n1740), .A4(
        \inq_ary[12][89] ), .Y(n114) );
  AO22X1_RVT U148 ( .A1(n1742), .A2(\inq_ary[3][89] ), .A3(n1751), .A4(
        \inq_ary[9][89] ), .Y(n113) );
  NOR4X1_RVT U149 ( .A1(n116), .A2(n115), .A3(n114), .A4(n113), .Y(n117) );
  NAND2X0_RVT U150 ( .A1(n118), .A2(n117), .Y(n119) );
  AO22X1_RVT U151 ( .A1(n3), .A2(wrdata_d1[89]), .A3(n969), .A4(n119), .Y(
        n3419) );
  AO22X1_RVT U152 ( .A1(n1537), .A2(\inq_ary[15][90] ), .A3(n1750), .A4(
        \inq_ary[11][90] ), .Y(n123) );
  AO22X1_RVT U153 ( .A1(n1742), .A2(\inq_ary[3][90] ), .A3(n1729), .A4(
        \inq_ary[4][90] ), .Y(n122) );
  AO22X1_RVT U154 ( .A1(n1612), .A2(\inq_ary[8][90] ), .A3(n1740), .A4(
        \inq_ary[12][90] ), .Y(n121) );
  AO22X1_RVT U155 ( .A1(n1749), .A2(\inq_ary[1][90] ), .A3(n1738), .A4(
        \inq_ary[6][90] ), .Y(n120) );
  NOR4X1_RVT U156 ( .A1(n123), .A2(n122), .A3(n121), .A4(n120), .Y(n129) );
  AO22X1_RVT U157 ( .A1(n1741), .A2(\inq_ary[7][90] ), .A3(n1747), .A4(
        \inq_ary[5][90] ), .Y(n127) );
  AO22X1_RVT U158 ( .A1(n1739), .A2(\inq_ary[2][90] ), .A3(n1554), .A4(
        \inq_ary[14][90] ), .Y(n126) );
  AO22X1_RVT U159 ( .A1(n1711), .A2(\inq_ary[13][90] ), .A3(n1748), .A4(
        \inq_ary[10][90] ), .Y(n125) );
  AO22X1_RVT U160 ( .A1(n1686), .A2(\inq_ary[0][90] ), .A3(n1751), .A4(
        \inq_ary[9][90] ), .Y(n124) );
  NOR4X1_RVT U161 ( .A1(n127), .A2(n126), .A3(n125), .A4(n124), .Y(n128) );
  NAND2X0_RVT U162 ( .A1(n129), .A2(n128), .Y(n130) );
  AO22X1_RVT U163 ( .A1(n1723), .A2(wrdata_d1[90]), .A3(n969), .A4(n130), .Y(
        n3421) );
  AO22X1_RVT U164 ( .A1(n1554), .A2(\inq_ary[14][91] ), .A3(n1711), .A4(
        \inq_ary[13][91] ), .Y(n134) );
  AO22X1_RVT U165 ( .A1(n1537), .A2(\inq_ary[15][91] ), .A3(n1741), .A4(
        \inq_ary[7][91] ), .Y(n133) );
  AO22X1_RVT U166 ( .A1(n1739), .A2(\inq_ary[2][91] ), .A3(n1751), .A4(
        \inq_ary[9][91] ), .Y(n132) );
  AO22X1_RVT U167 ( .A1(n1740), .A2(\inq_ary[12][91] ), .A3(n1747), .A4(
        \inq_ary[5][91] ), .Y(n131) );
  NOR4X1_RVT U168 ( .A1(n134), .A2(n133), .A3(n132), .A4(n131), .Y(n140) );
  AO22X1_RVT U169 ( .A1(n1612), .A2(\inq_ary[8][91] ), .A3(n1748), .A4(
        \inq_ary[10][91] ), .Y(n138) );
  AO22X1_RVT U170 ( .A1(n1742), .A2(\inq_ary[3][91] ), .A3(n1686), .A4(
        \inq_ary[0][91] ), .Y(n137) );
  AO22X1_RVT U171 ( .A1(n1750), .A2(\inq_ary[11][91] ), .A3(n1738), .A4(
        \inq_ary[6][91] ), .Y(n136) );
  AO22X1_RVT U172 ( .A1(n1729), .A2(\inq_ary[4][91] ), .A3(n1749), .A4(
        \inq_ary[1][91] ), .Y(n135) );
  NOR4X1_RVT U173 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .Y(n139) );
  NAND2X0_RVT U174 ( .A1(n140), .A2(n139), .Y(n141) );
  AO22X1_RVT U175 ( .A1(n1684), .A2(wrdata_d1[91]), .A3(n969), .A4(n141), .Y(
        n3423) );
  AO22X1_RVT U176 ( .A1(n1741), .A2(\inq_ary[7][44] ), .A3(n1747), .A4(
        \inq_ary[5][44] ), .Y(n145) );
  AO22X1_RVT U177 ( .A1(n1554), .A2(\inq_ary[14][44] ), .A3(n1751), .A4(
        \inq_ary[9][44] ), .Y(n144) );
  AO22X1_RVT U178 ( .A1(n1612), .A2(\inq_ary[8][44] ), .A3(n1711), .A4(
        \inq_ary[13][44] ), .Y(n143) );
  AO22X1_RVT U179 ( .A1(n1739), .A2(\inq_ary[2][44] ), .A3(n1686), .A4(
        \inq_ary[0][44] ), .Y(n142) );
  NOR4X1_RVT U180 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .Y(n151) );
  AO22X1_RVT U181 ( .A1(n1742), .A2(\inq_ary[3][44] ), .A3(n1750), .A4(
        \inq_ary[11][44] ), .Y(n149) );
  AO22X1_RVT U182 ( .A1(n1729), .A2(\inq_ary[4][44] ), .A3(n1749), .A4(
        \inq_ary[1][44] ), .Y(n148) );
  AO22X1_RVT U183 ( .A1(n1537), .A2(\inq_ary[15][44] ), .A3(n1748), .A4(
        \inq_ary[10][44] ), .Y(n147) );
  AO22X1_RVT U184 ( .A1(n1740), .A2(\inq_ary[12][44] ), .A3(n1738), .A4(
        \inq_ary[6][44] ), .Y(n146) );
  NOR4X1_RVT U185 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .Y(n150) );
  NAND2X0_RVT U186 ( .A1(n151), .A2(n150), .Y(n152) );
  AO22X1_RVT U187 ( .A1(n1598), .A2(wrdata_d1[44]), .A3(n2), .A4(n152), .Y(
        n3375) );
  INVX1_RVT U188 ( .A(n946), .Y(n1025) );
  AO22X1_RVT U189 ( .A1(n1686), .A2(\inq_ary[0][92] ), .A3(n1537), .A4(
        \inq_ary[15][92] ), .Y(n156) );
  AO22X1_RVT U190 ( .A1(n1739), .A2(\inq_ary[2][92] ), .A3(n1747), .A4(
        \inq_ary[5][92] ), .Y(n155) );
  AO22X1_RVT U191 ( .A1(n1742), .A2(\inq_ary[3][92] ), .A3(n1749), .A4(
        \inq_ary[1][92] ), .Y(n154) );
  AO22X1_RVT U192 ( .A1(n1750), .A2(\inq_ary[11][92] ), .A3(n1738), .A4(
        \inq_ary[6][92] ), .Y(n153) );
  NOR4X1_RVT U193 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .Y(n162) );
  AO22X1_RVT U194 ( .A1(n1729), .A2(\inq_ary[4][92] ), .A3(n1748), .A4(
        \inq_ary[10][92] ), .Y(n160) );
  AO22X1_RVT U195 ( .A1(n1741), .A2(\inq_ary[7][92] ), .A3(n1711), .A4(
        \inq_ary[13][92] ), .Y(n159) );
  AO22X1_RVT U196 ( .A1(n1554), .A2(\inq_ary[14][92] ), .A3(n1751), .A4(
        \inq_ary[9][92] ), .Y(n158) );
  AO22X1_RVT U197 ( .A1(n1612), .A2(\inq_ary[8][92] ), .A3(n1740), .A4(
        \inq_ary[12][92] ), .Y(n157) );
  NOR4X1_RVT U198 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .Y(n161) );
  NAND2X0_RVT U199 ( .A1(n162), .A2(n161), .Y(n163) );
  AO22X1_RVT U200 ( .A1(n1025), .A2(wrdata_d1[92]), .A3(n969), .A4(n163), .Y(
        n3416) );
  AO22X1_RVT U201 ( .A1(n1749), .A2(\inq_ary[1][93] ), .A3(n1748), .A4(
        \inq_ary[10][93] ), .Y(n167) );
  AO22X1_RVT U202 ( .A1(n1729), .A2(\inq_ary[4][93] ), .A3(n1740), .A4(
        \inq_ary[12][93] ), .Y(n166) );
  AO22X1_RVT U203 ( .A1(n1686), .A2(\inq_ary[0][93] ), .A3(n1741), .A4(
        \inq_ary[7][93] ), .Y(n165) );
  AO22X1_RVT U204 ( .A1(n1537), .A2(\inq_ary[15][93] ), .A3(n1612), .A4(
        \inq_ary[8][93] ), .Y(n164) );
  NOR4X1_RVT U205 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .Y(n173) );
  AO22X1_RVT U206 ( .A1(n1739), .A2(\inq_ary[2][93] ), .A3(n1751), .A4(
        \inq_ary[9][93] ), .Y(n171) );
  AO22X1_RVT U207 ( .A1(n1554), .A2(\inq_ary[14][93] ), .A3(n1711), .A4(
        \inq_ary[13][93] ), .Y(n170) );
  AO22X1_RVT U208 ( .A1(n1747), .A2(\inq_ary[5][93] ), .A3(n1750), .A4(
        \inq_ary[11][93] ), .Y(n169) );
  AO22X1_RVT U209 ( .A1(n1742), .A2(\inq_ary[3][93] ), .A3(n1738), .A4(
        \inq_ary[6][93] ), .Y(n168) );
  NOR4X1_RVT U210 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .Y(n172) );
  NAND2X0_RVT U211 ( .A1(n173), .A2(n172), .Y(n174) );
  AO22X1_RVT U212 ( .A1(n3), .A2(wrdata_d1[93]), .A3(n946), .A4(n174), .Y(
        n3418) );
  AO22X1_RVT U213 ( .A1(n1554), .A2(\inq_ary[14][43] ), .A3(n1711), .A4(
        \inq_ary[13][43] ), .Y(n178) );
  AO22X1_RVT U214 ( .A1(n1750), .A2(\inq_ary[11][43] ), .A3(n1751), .A4(
        \inq_ary[9][43] ), .Y(n177) );
  AO22X1_RVT U215 ( .A1(n1740), .A2(\inq_ary[12][43] ), .A3(n1741), .A4(
        \inq_ary[7][43] ), .Y(n176) );
  AO22X1_RVT U216 ( .A1(n1749), .A2(\inq_ary[1][43] ), .A3(n1747), .A4(
        \inq_ary[5][43] ), .Y(n175) );
  NOR4X1_RVT U217 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .Y(n184) );
  AO22X1_RVT U218 ( .A1(n1739), .A2(\inq_ary[2][43] ), .A3(n1729), .A4(
        \inq_ary[4][43] ), .Y(n182) );
  AO22X1_RVT U219 ( .A1(n1742), .A2(\inq_ary[3][43] ), .A3(n1686), .A4(
        \inq_ary[0][43] ), .Y(n181) );
  AO22X1_RVT U220 ( .A1(n1738), .A2(\inq_ary[6][43] ), .A3(n1748), .A4(
        \inq_ary[10][43] ), .Y(n180) );
  AO22X1_RVT U221 ( .A1(n1537), .A2(\inq_ary[15][43] ), .A3(n1612), .A4(
        \inq_ary[8][43] ), .Y(n179) );
  NOR4X1_RVT U222 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .Y(n183) );
  NAND2X0_RVT U223 ( .A1(n184), .A2(n183), .Y(n185) );
  AO22X1_RVT U224 ( .A1(n1598), .A2(wrdata_d1[43]), .A3(n2), .A4(n185), .Y(
        n3382) );
  AO22X1_RVT U225 ( .A1(n1554), .A2(\inq_ary[14][94] ), .A3(n1742), .A4(
        \inq_ary[3][94] ), .Y(n189) );
  AO22X1_RVT U226 ( .A1(n1740), .A2(\inq_ary[12][94] ), .A3(n1748), .A4(
        \inq_ary[10][94] ), .Y(n188) );
  AO22X1_RVT U227 ( .A1(n1612), .A2(\inq_ary[8][94] ), .A3(n1747), .A4(
        \inq_ary[5][94] ), .Y(n187) );
  AO22X1_RVT U228 ( .A1(n1686), .A2(\inq_ary[0][94] ), .A3(n1751), .A4(
        \inq_ary[9][94] ), .Y(n186) );
  NOR4X1_RVT U229 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .Y(n195) );
  AO22X1_RVT U230 ( .A1(n1739), .A2(\inq_ary[2][94] ), .A3(n1738), .A4(
        \inq_ary[6][94] ), .Y(n193) );
  AO22X1_RVT U231 ( .A1(n1749), .A2(\inq_ary[1][94] ), .A3(n1711), .A4(
        \inq_ary[13][94] ), .Y(n192) );
  AO22X1_RVT U232 ( .A1(n1729), .A2(\inq_ary[4][94] ), .A3(n1741), .A4(
        \inq_ary[7][94] ), .Y(n191) );
  AO22X1_RVT U233 ( .A1(n1537), .A2(\inq_ary[15][94] ), .A3(n1750), .A4(
        \inq_ary[11][94] ), .Y(n190) );
  NOR4X1_RVT U234 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .Y(n194) );
  NAND2X0_RVT U235 ( .A1(n195), .A2(n194), .Y(n196) );
  AO22X1_RVT U236 ( .A1(n758), .A2(wrdata_d1[94]), .A3(n969), .A4(n196), .Y(
        n3420) );
  AO22X1_RVT U237 ( .A1(n1729), .A2(\inq_ary[4][95] ), .A3(n1711), .A4(
        \inq_ary[13][95] ), .Y(n200) );
  AO22X1_RVT U238 ( .A1(n1537), .A2(\inq_ary[15][95] ), .A3(n1738), .A4(
        \inq_ary[6][95] ), .Y(n199) );
  AO22X1_RVT U239 ( .A1(n1686), .A2(\inq_ary[0][95] ), .A3(n1748), .A4(
        \inq_ary[10][95] ), .Y(n198) );
  AO22X1_RVT U240 ( .A1(n1554), .A2(\inq_ary[14][95] ), .A3(n1751), .A4(
        \inq_ary[9][95] ), .Y(n197) );
  NOR4X1_RVT U241 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .Y(n206) );
  AO22X1_RVT U242 ( .A1(n1749), .A2(\inq_ary[1][95] ), .A3(n1741), .A4(
        \inq_ary[7][95] ), .Y(n204) );
  AO22X1_RVT U243 ( .A1(n1739), .A2(\inq_ary[2][95] ), .A3(n1747), .A4(
        \inq_ary[5][95] ), .Y(n203) );
  AO22X1_RVT U244 ( .A1(n1742), .A2(\inq_ary[3][95] ), .A3(n1740), .A4(
        \inq_ary[12][95] ), .Y(n202) );
  AO22X1_RVT U245 ( .A1(n1612), .A2(\inq_ary[8][95] ), .A3(n1750), .A4(
        \inq_ary[11][95] ), .Y(n201) );
  NOR4X1_RVT U246 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .Y(n205) );
  NAND2X0_RVT U247 ( .A1(n206), .A2(n205), .Y(n207) );
  AO22X1_RVT U248 ( .A1(n1025), .A2(wrdata_d1[95]), .A3(n2), .A4(n207), .Y(
        n3422) );
  AO22X1_RVT U249 ( .A1(n1686), .A2(\inq_ary[0][42] ), .A3(n1612), .A4(
        \inq_ary[8][42] ), .Y(n211) );
  AO22X1_RVT U250 ( .A1(n1750), .A2(\inq_ary[11][42] ), .A3(n1711), .A4(
        \inq_ary[13][42] ), .Y(n210) );
  AO22X1_RVT U251 ( .A1(n1749), .A2(\inq_ary[1][42] ), .A3(n1741), .A4(
        \inq_ary[7][42] ), .Y(n209) );
  AO22X1_RVT U252 ( .A1(n1742), .A2(\inq_ary[3][42] ), .A3(n1537), .A4(
        \inq_ary[15][42] ), .Y(n208) );
  NOR4X1_RVT U253 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .Y(n217) );
  AO22X1_RVT U254 ( .A1(n1729), .A2(\inq_ary[4][42] ), .A3(n1748), .A4(
        \inq_ary[10][42] ), .Y(n215) );
  AO22X1_RVT U255 ( .A1(n1738), .A2(\inq_ary[6][42] ), .A3(n1751), .A4(
        \inq_ary[9][42] ), .Y(n214) );
  AO22X1_RVT U256 ( .A1(n1554), .A2(\inq_ary[14][42] ), .A3(n1747), .A4(
        \inq_ary[5][42] ), .Y(n213) );
  AO22X1_RVT U257 ( .A1(n1739), .A2(\inq_ary[2][42] ), .A3(n1740), .A4(
        \inq_ary[12][42] ), .Y(n212) );
  NOR4X1_RVT U258 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .Y(n216) );
  NAND2X0_RVT U259 ( .A1(n217), .A2(n216), .Y(n218) );
  AO22X1_RVT U260 ( .A1(n1598), .A2(wrdata_d1[42]), .A3(n1489), .A4(n218), .Y(
        n3380) );
  AO22X1_RVT U261 ( .A1(n1739), .A2(\inq_ary[2][102] ), .A3(n1751), .A4(
        \inq_ary[9][102] ), .Y(n222) );
  AO22X1_RVT U262 ( .A1(n1554), .A2(\inq_ary[14][102] ), .A3(n1537), .A4(
        \inq_ary[15][102] ), .Y(n221) );
  AO22X1_RVT U263 ( .A1(n1740), .A2(\inq_ary[12][102] ), .A3(n1748), .A4(
        \inq_ary[10][102] ), .Y(n220) );
  AO22X1_RVT U264 ( .A1(n1747), .A2(\inq_ary[5][102] ), .A3(n1711), .A4(
        \inq_ary[13][102] ), .Y(n219) );
  NOR4X1_RVT U265 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .Y(n228) );
  AO22X1_RVT U266 ( .A1(n1729), .A2(\inq_ary[4][102] ), .A3(n1749), .A4(
        \inq_ary[1][102] ), .Y(n226) );
  AO22X1_RVT U267 ( .A1(n1742), .A2(\inq_ary[3][102] ), .A3(n1612), .A4(
        \inq_ary[8][102] ), .Y(n225) );
  AO22X1_RVT U268 ( .A1(n1686), .A2(\inq_ary[0][102] ), .A3(n1738), .A4(
        \inq_ary[6][102] ), .Y(n224) );
  AO22X1_RVT U269 ( .A1(n1741), .A2(\inq_ary[7][102] ), .A3(n1750), .A4(
        \inq_ary[11][102] ), .Y(n223) );
  NOR4X1_RVT U270 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .Y(n227) );
  NAND2X0_RVT U271 ( .A1(n228), .A2(n227), .Y(n229) );
  AO22X1_RVT U272 ( .A1(n758), .A2(wrdata_d1[102]), .A3(n2), .A4(n229), .Y(
        n3428) );
  AO22X1_RVT U273 ( .A1(n1729), .A2(\inq_ary[4][110] ), .A3(n1612), .A4(
        \inq_ary[8][110] ), .Y(n233) );
  AO22X1_RVT U274 ( .A1(n1739), .A2(\inq_ary[2][110] ), .A3(n1686), .A4(
        \inq_ary[0][110] ), .Y(n232) );
  AO22X1_RVT U275 ( .A1(n1740), .A2(\inq_ary[12][110] ), .A3(n1711), .A4(
        \inq_ary[13][110] ), .Y(n231) );
  AO22X1_RVT U276 ( .A1(n1749), .A2(\inq_ary[1][110] ), .A3(n1741), .A4(
        \inq_ary[7][110] ), .Y(n230) );
  NOR4X1_RVT U277 ( .A1(n233), .A2(n232), .A3(n231), .A4(n230), .Y(n239) );
  AO22X1_RVT U278 ( .A1(n1554), .A2(\inq_ary[14][110] ), .A3(n1537), .A4(
        \inq_ary[15][110] ), .Y(n237) );
  AO22X1_RVT U279 ( .A1(n1747), .A2(\inq_ary[5][110] ), .A3(n1748), .A4(
        \inq_ary[10][110] ), .Y(n236) );
  AO22X1_RVT U280 ( .A1(n1750), .A2(\inq_ary[11][110] ), .A3(n1738), .A4(
        \inq_ary[6][110] ), .Y(n235) );
  AO22X1_RVT U281 ( .A1(n1742), .A2(\inq_ary[3][110] ), .A3(n1751), .A4(
        \inq_ary[9][110] ), .Y(n234) );
  NOR4X1_RVT U282 ( .A1(n237), .A2(n236), .A3(n235), .A4(n234), .Y(n238) );
  NAND2X0_RVT U283 ( .A1(n239), .A2(n238), .Y(n240) );
  AO22X1_RVT U284 ( .A1(n3), .A2(wrdata_d1[110]), .A3(n1), .A4(n240), .Y(n3436) );
  AO22X1_RVT U285 ( .A1(n1742), .A2(\inq_ary[3][111] ), .A3(n1748), .A4(
        \inq_ary[10][111] ), .Y(n244) );
  AO22X1_RVT U286 ( .A1(n1537), .A2(\inq_ary[15][111] ), .A3(n1612), .A4(
        \inq_ary[8][111] ), .Y(n243) );
  AO22X1_RVT U287 ( .A1(n1749), .A2(\inq_ary[1][111] ), .A3(n1711), .A4(
        \inq_ary[13][111] ), .Y(n242) );
  AO22X1_RVT U288 ( .A1(n1739), .A2(\inq_ary[2][111] ), .A3(n1751), .A4(
        \inq_ary[9][111] ), .Y(n241) );
  NOR4X1_RVT U289 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .Y(n250) );
  AO22X1_RVT U290 ( .A1(n1686), .A2(\inq_ary[0][111] ), .A3(n1738), .A4(
        \inq_ary[6][111] ), .Y(n248) );
  AO22X1_RVT U291 ( .A1(n1741), .A2(\inq_ary[7][111] ), .A3(n1747), .A4(
        \inq_ary[5][111] ), .Y(n247) );
  AO22X1_RVT U292 ( .A1(n1554), .A2(\inq_ary[14][111] ), .A3(n1740), .A4(
        \inq_ary[12][111] ), .Y(n246) );
  AO22X1_RVT U293 ( .A1(n1729), .A2(\inq_ary[4][111] ), .A3(n1750), .A4(
        \inq_ary[11][111] ), .Y(n245) );
  NOR4X1_RVT U294 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .Y(n249) );
  NAND2X0_RVT U295 ( .A1(n250), .A2(n249), .Y(n251) );
  AO22X1_RVT U296 ( .A1(n1684), .A2(wrdata_d1[111]), .A3(n1), .A4(n251), .Y(
        n3438) );
  AO22X1_RVT U297 ( .A1(n1729), .A2(\inq_ary[4][34] ), .A3(n1749), .A4(
        \inq_ary[1][34] ), .Y(n255) );
  AO22X1_RVT U298 ( .A1(n1554), .A2(\inq_ary[14][34] ), .A3(n1738), .A4(
        \inq_ary[6][34] ), .Y(n254) );
  AO22X1_RVT U299 ( .A1(n1537), .A2(\inq_ary[15][34] ), .A3(n1740), .A4(
        \inq_ary[12][34] ), .Y(n253) );
  AO22X1_RVT U300 ( .A1(n1747), .A2(\inq_ary[5][34] ), .A3(n1748), .A4(
        \inq_ary[10][34] ), .Y(n252) );
  NOR4X1_RVT U301 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .Y(n261) );
  AO22X1_RVT U302 ( .A1(n1686), .A2(\inq_ary[0][34] ), .A3(n1741), .A4(
        \inq_ary[7][34] ), .Y(n259) );
  AO22X1_RVT U303 ( .A1(n1742), .A2(\inq_ary[3][34] ), .A3(n1750), .A4(
        \inq_ary[11][34] ), .Y(n258) );
  AO22X1_RVT U304 ( .A1(n1739), .A2(\inq_ary[2][34] ), .A3(n1612), .A4(
        \inq_ary[8][34] ), .Y(n257) );
  AO22X1_RVT U305 ( .A1(n1711), .A2(\inq_ary[13][34] ), .A3(n1751), .A4(
        \inq_ary[9][34] ), .Y(n256) );
  NOR4X1_RVT U306 ( .A1(n259), .A2(n258), .A3(n257), .A4(n256), .Y(n260) );
  NAND2X0_RVT U307 ( .A1(n261), .A2(n260), .Y(n262) );
  AO22X1_RVT U308 ( .A1(n1477), .A2(wrdata_d1[34]), .A3(n2), .A4(n262), .Y(
        n3372) );
  INVX1_RVT U309 ( .A(n946), .Y(n1477) );
  AO22X1_RVT U310 ( .A1(n1729), .A2(\inq_ary[4][112] ), .A3(n1749), .A4(
        \inq_ary[1][112] ), .Y(n266) );
  AO22X1_RVT U311 ( .A1(n1554), .A2(\inq_ary[14][112] ), .A3(n1740), .A4(
        \inq_ary[12][112] ), .Y(n265) );
  AO22X1_RVT U312 ( .A1(n1742), .A2(\inq_ary[3][112] ), .A3(n1751), .A4(
        \inq_ary[9][112] ), .Y(n264) );
  AO22X1_RVT U313 ( .A1(n1612), .A2(\inq_ary[8][112] ), .A3(n1738), .A4(
        \inq_ary[6][112] ), .Y(n263) );
  NOR4X1_RVT U314 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .Y(n272) );
  AO22X1_RVT U315 ( .A1(n1686), .A2(\inq_ary[0][112] ), .A3(n1748), .A4(
        \inq_ary[10][112] ), .Y(n270) );
  AO22X1_RVT U316 ( .A1(n1739), .A2(\inq_ary[2][112] ), .A3(n1537), .A4(
        \inq_ary[15][112] ), .Y(n269) );
  AO22X1_RVT U317 ( .A1(n1741), .A2(\inq_ary[7][112] ), .A3(n1711), .A4(
        \inq_ary[13][112] ), .Y(n268) );
  AO22X1_RVT U318 ( .A1(n1747), .A2(\inq_ary[5][112] ), .A3(n1750), .A4(
        \inq_ary[11][112] ), .Y(n267) );
  NOR4X1_RVT U319 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .Y(n271) );
  NAND2X0_RVT U320 ( .A1(n272), .A2(n271), .Y(n273) );
  AO22X1_RVT U321 ( .A1(n1477), .A2(wrdata_d1[112]), .A3(n1), .A4(n273), .Y(
        n3441) );
  AO22X1_RVT U322 ( .A1(n1742), .A2(\inq_ary[3][113] ), .A3(n1686), .A4(
        \inq_ary[0][113] ), .Y(n277) );
  AO22X1_RVT U323 ( .A1(n1739), .A2(\inq_ary[2][113] ), .A3(n1740), .A4(
        \inq_ary[12][113] ), .Y(n276) );
  AO22X1_RVT U324 ( .A1(n1729), .A2(\inq_ary[4][113] ), .A3(n1751), .A4(
        \inq_ary[9][113] ), .Y(n275) );
  AO22X1_RVT U325 ( .A1(n1554), .A2(\inq_ary[14][113] ), .A3(n1750), .A4(
        \inq_ary[11][113] ), .Y(n274) );
  NOR4X1_RVT U326 ( .A1(n277), .A2(n276), .A3(n275), .A4(n274), .Y(n283) );
  AO22X1_RVT U327 ( .A1(n1612), .A2(\inq_ary[8][113] ), .A3(n1738), .A4(
        \inq_ary[6][113] ), .Y(n281) );
  AO22X1_RVT U328 ( .A1(n1749), .A2(\inq_ary[1][113] ), .A3(n1741), .A4(
        \inq_ary[7][113] ), .Y(n280) );
  AO22X1_RVT U329 ( .A1(n1747), .A2(\inq_ary[5][113] ), .A3(n1748), .A4(
        \inq_ary[10][113] ), .Y(n279) );
  AO22X1_RVT U330 ( .A1(n1537), .A2(\inq_ary[15][113] ), .A3(n1711), .A4(
        \inq_ary[13][113] ), .Y(n278) );
  NOR4X1_RVT U331 ( .A1(n281), .A2(n280), .A3(n279), .A4(n278), .Y(n282) );
  NAND2X0_RVT U332 ( .A1(n283), .A2(n282), .Y(n284) );
  AO22X1_RVT U333 ( .A1(n1477), .A2(wrdata_d1[113]), .A3(n1), .A4(n284), .Y(
        n3443) );
  AO22X1_RVT U334 ( .A1(n1742), .A2(\inq_ary[3][33] ), .A3(n1740), .A4(
        \inq_ary[12][33] ), .Y(n288) );
  AO22X1_RVT U335 ( .A1(n1738), .A2(\inq_ary[6][33] ), .A3(n1751), .A4(
        \inq_ary[9][33] ), .Y(n287) );
  AO22X1_RVT U336 ( .A1(n1741), .A2(\inq_ary[7][33] ), .A3(n1750), .A4(
        \inq_ary[11][33] ), .Y(n286) );
  AO22X1_RVT U337 ( .A1(n1686), .A2(\inq_ary[0][33] ), .A3(n1748), .A4(
        \inq_ary[10][33] ), .Y(n285) );
  NOR4X1_RVT U338 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .Y(n294) );
  AO22X1_RVT U339 ( .A1(n1749), .A2(\inq_ary[1][33] ), .A3(n1711), .A4(
        \inq_ary[13][33] ), .Y(n292) );
  AO22X1_RVT U340 ( .A1(n1739), .A2(\inq_ary[2][33] ), .A3(n1612), .A4(
        \inq_ary[8][33] ), .Y(n291) );
  AO22X1_RVT U341 ( .A1(n1729), .A2(\inq_ary[4][33] ), .A3(n1537), .A4(
        \inq_ary[15][33] ), .Y(n290) );
  AO22X1_RVT U342 ( .A1(n1554), .A2(\inq_ary[14][33] ), .A3(n1747), .A4(
        \inq_ary[5][33] ), .Y(n289) );
  NOR4X1_RVT U343 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .Y(n293) );
  NAND2X0_RVT U344 ( .A1(n294), .A2(n293), .Y(n295) );
  AO22X1_RVT U345 ( .A1(n3), .A2(wrdata_d1[33]), .A3(n2), .A4(n295), .Y(n3370)
         );
  INVX1_RVT U346 ( .A(n946), .Y(n1684) );
  AO22X1_RVT U347 ( .A1(n1741), .A2(\inq_ary[7][114] ), .A3(n1748), .A4(
        \inq_ary[10][114] ), .Y(n299) );
  AO22X1_RVT U348 ( .A1(n1537), .A2(\inq_ary[15][114] ), .A3(n1749), .A4(
        \inq_ary[1][114] ), .Y(n298) );
  AO22X1_RVT U349 ( .A1(n1686), .A2(\inq_ary[0][114] ), .A3(n1740), .A4(
        \inq_ary[12][114] ), .Y(n297) );
  AO22X1_RVT U350 ( .A1(n1747), .A2(\inq_ary[5][114] ), .A3(n1750), .A4(
        \inq_ary[11][114] ), .Y(n296) );
  NOR4X1_RVT U351 ( .A1(n299), .A2(n298), .A3(n297), .A4(n296), .Y(n305) );
  AO22X1_RVT U352 ( .A1(n1729), .A2(\inq_ary[4][114] ), .A3(n1751), .A4(
        \inq_ary[9][114] ), .Y(n303) );
  AO22X1_RVT U353 ( .A1(n1554), .A2(\inq_ary[14][114] ), .A3(n1742), .A4(
        \inq_ary[3][114] ), .Y(n302) );
  AO22X1_RVT U354 ( .A1(n1739), .A2(\inq_ary[2][114] ), .A3(n1738), .A4(
        \inq_ary[6][114] ), .Y(n301) );
  AO22X1_RVT U355 ( .A1(n1612), .A2(\inq_ary[8][114] ), .A3(n1711), .A4(
        \inq_ary[13][114] ), .Y(n300) );
  NOR4X1_RVT U356 ( .A1(n303), .A2(n302), .A3(n301), .A4(n300), .Y(n304) );
  NAND2X0_RVT U357 ( .A1(n305), .A2(n304), .Y(n306) );
  AO22X1_RVT U358 ( .A1(n1684), .A2(wrdata_d1[114]), .A3(n1), .A4(n306), .Y(
        n3445) );
  AO22X1_RVT U359 ( .A1(n1739), .A2(\inq_ary[2][115] ), .A3(n1742), .A4(
        \inq_ary[3][115] ), .Y(n310) );
  AO22X1_RVT U360 ( .A1(n1749), .A2(\inq_ary[1][115] ), .A3(n1738), .A4(
        \inq_ary[6][115] ), .Y(n309) );
  AO22X1_RVT U361 ( .A1(n1729), .A2(\inq_ary[4][115] ), .A3(n1686), .A4(
        \inq_ary[0][115] ), .Y(n308) );
  AO22X1_RVT U362 ( .A1(n1711), .A2(\inq_ary[13][115] ), .A3(n1748), .A4(
        \inq_ary[10][115] ), .Y(n307) );
  NOR4X1_RVT U363 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .Y(n316) );
  AO22X1_RVT U364 ( .A1(n1554), .A2(\inq_ary[14][115] ), .A3(n1612), .A4(
        \inq_ary[8][115] ), .Y(n314) );
  AO22X1_RVT U365 ( .A1(n1750), .A2(\inq_ary[11][115] ), .A3(n1751), .A4(
        \inq_ary[9][115] ), .Y(n313) );
  AO22X1_RVT U366 ( .A1(n1740), .A2(\inq_ary[12][115] ), .A3(n1747), .A4(
        \inq_ary[5][115] ), .Y(n312) );
  AO22X1_RVT U367 ( .A1(n1537), .A2(\inq_ary[15][115] ), .A3(n1741), .A4(
        \inq_ary[7][115] ), .Y(n311) );
  NOR4X1_RVT U368 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .Y(n315) );
  NAND2X0_RVT U369 ( .A1(n316), .A2(n315), .Y(n317) );
  AO22X1_RVT U370 ( .A1(n1684), .A2(wrdata_d1[115]), .A3(n1), .A4(n317), .Y(
        n3447) );
  AO22X1_RVT U371 ( .A1(n1749), .A2(\inq_ary[1][32] ), .A3(n1747), .A4(
        \inq_ary[5][32] ), .Y(n321) );
  AO22X1_RVT U372 ( .A1(n1739), .A2(\inq_ary[2][32] ), .A3(n1738), .A4(
        \inq_ary[6][32] ), .Y(n320) );
  AO22X1_RVT U373 ( .A1(n1612), .A2(\inq_ary[8][32] ), .A3(n1711), .A4(
        \inq_ary[13][32] ), .Y(n319) );
  AO22X1_RVT U374 ( .A1(n1729), .A2(\inq_ary[4][32] ), .A3(n1740), .A4(
        \inq_ary[12][32] ), .Y(n318) );
  NOR4X1_RVT U375 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .Y(n327) );
  AO22X1_RVT U376 ( .A1(n1554), .A2(\inq_ary[14][32] ), .A3(n1741), .A4(
        \inq_ary[7][32] ), .Y(n325) );
  AO22X1_RVT U377 ( .A1(n1742), .A2(\inq_ary[3][32] ), .A3(n1751), .A4(
        \inq_ary[9][32] ), .Y(n324) );
  AO22X1_RVT U378 ( .A1(n1686), .A2(\inq_ary[0][32] ), .A3(n1750), .A4(
        \inq_ary[11][32] ), .Y(n323) );
  AO22X1_RVT U379 ( .A1(n1537), .A2(\inq_ary[15][32] ), .A3(n1748), .A4(
        \inq_ary[10][32] ), .Y(n322) );
  NOR4X1_RVT U380 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .Y(n326) );
  NAND2X0_RVT U381 ( .A1(n327), .A2(n326), .Y(n328) );
  AO22X1_RVT U382 ( .A1(n1025), .A2(wrdata_d1[32]), .A3(n2), .A4(n328), .Y(
        n3368) );
  AO22X1_RVT U383 ( .A1(n1740), .A2(\inq_ary[12][116] ), .A3(n1741), .A4(
        \inq_ary[7][116] ), .Y(n332) );
  AO22X1_RVT U384 ( .A1(n1739), .A2(\inq_ary[2][116] ), .A3(n1686), .A4(
        \inq_ary[0][116] ), .Y(n331) );
  AO22X1_RVT U385 ( .A1(n1554), .A2(\inq_ary[14][116] ), .A3(n1729), .A4(
        \inq_ary[4][116] ), .Y(n330) );
  AO22X1_RVT U386 ( .A1(n1749), .A2(\inq_ary[1][116] ), .A3(n1751), .A4(
        \inq_ary[9][116] ), .Y(n329) );
  NOR4X1_RVT U387 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .Y(n338) );
  AO22X1_RVT U388 ( .A1(n1537), .A2(\inq_ary[15][116] ), .A3(n1750), .A4(
        \inq_ary[11][116] ), .Y(n336) );
  AO22X1_RVT U389 ( .A1(n1612), .A2(\inq_ary[8][116] ), .A3(n1748), .A4(
        \inq_ary[10][116] ), .Y(n335) );
  AO22X1_RVT U390 ( .A1(n1742), .A2(\inq_ary[3][116] ), .A3(n1738), .A4(
        \inq_ary[6][116] ), .Y(n334) );
  AO22X1_RVT U391 ( .A1(n1747), .A2(\inq_ary[5][116] ), .A3(n1711), .A4(
        \inq_ary[13][116] ), .Y(n333) );
  NOR4X1_RVT U392 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .Y(n337) );
  NAND2X0_RVT U393 ( .A1(n338), .A2(n337), .Y(n339) );
  AO22X1_RVT U394 ( .A1(n1477), .A2(wrdata_d1[116]), .A3(n1), .A4(n339), .Y(
        n3440) );
  AO22X1_RVT U395 ( .A1(n1738), .A2(\inq_ary[6][103] ), .A3(n1751), .A4(
        \inq_ary[9][103] ), .Y(n343) );
  AO22X1_RVT U396 ( .A1(n1741), .A2(\inq_ary[7][103] ), .A3(n1747), .A4(
        \inq_ary[5][103] ), .Y(n342) );
  AO22X1_RVT U397 ( .A1(n1554), .A2(\inq_ary[14][103] ), .A3(n1742), .A4(
        \inq_ary[3][103] ), .Y(n341) );
  AO22X1_RVT U398 ( .A1(n1711), .A2(\inq_ary[13][103] ), .A3(n1748), .A4(
        \inq_ary[10][103] ), .Y(n340) );
  NOR4X1_RVT U399 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .Y(n349) );
  AO22X1_RVT U400 ( .A1(n1740), .A2(\inq_ary[12][103] ), .A3(n1749), .A4(
        \inq_ary[1][103] ), .Y(n347) );
  AO22X1_RVT U401 ( .A1(n1729), .A2(\inq_ary[4][103] ), .A3(n1537), .A4(
        \inq_ary[15][103] ), .Y(n346) );
  AO22X1_RVT U402 ( .A1(n1739), .A2(\inq_ary[2][103] ), .A3(n1686), .A4(
        \inq_ary[0][103] ), .Y(n345) );
  AO22X1_RVT U403 ( .A1(n1612), .A2(\inq_ary[8][103] ), .A3(n1750), .A4(
        \inq_ary[11][103] ), .Y(n344) );
  NOR4X1_RVT U404 ( .A1(n347), .A2(n346), .A3(n345), .A4(n344), .Y(n348) );
  NAND2X0_RVT U405 ( .A1(n349), .A2(n348), .Y(n350) );
  AO22X1_RVT U406 ( .A1(n3), .A2(wrdata_d1[103]), .A3(n1), .A4(n350), .Y(n3430) );
  AO22X1_RVT U407 ( .A1(n1612), .A2(\inq_ary[8][104] ), .A3(n1748), .A4(
        \inq_ary[10][104] ), .Y(n354) );
  AO22X1_RVT U408 ( .A1(n1742), .A2(\inq_ary[3][104] ), .A3(n1741), .A4(
        \inq_ary[7][104] ), .Y(n353) );
  AO22X1_RVT U409 ( .A1(n1729), .A2(\inq_ary[4][104] ), .A3(n1738), .A4(
        \inq_ary[6][104] ), .Y(n352) );
  AO22X1_RVT U410 ( .A1(n1554), .A2(\inq_ary[14][104] ), .A3(n1686), .A4(
        \inq_ary[0][104] ), .Y(n351) );
  NOR4X1_RVT U411 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .Y(n360) );
  AO22X1_RVT U412 ( .A1(n1739), .A2(\inq_ary[2][104] ), .A3(n1711), .A4(
        \inq_ary[13][104] ), .Y(n358) );
  AO22X1_RVT U413 ( .A1(n1740), .A2(\inq_ary[12][104] ), .A3(n1750), .A4(
        \inq_ary[11][104] ), .Y(n357) );
  AO22X1_RVT U414 ( .A1(n1749), .A2(\inq_ary[1][104] ), .A3(n1751), .A4(
        \inq_ary[9][104] ), .Y(n356) );
  AO22X1_RVT U415 ( .A1(n1537), .A2(\inq_ary[15][104] ), .A3(n1747), .A4(
        \inq_ary[5][104] ), .Y(n355) );
  NOR4X1_RVT U416 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .Y(n359) );
  NAND2X0_RVT U417 ( .A1(n360), .A2(n359), .Y(n361) );
  AO22X1_RVT U418 ( .A1(n1723), .A2(wrdata_d1[104]), .A3(n1), .A4(n361), .Y(
        n3433) );
  AO22X1_RVT U419 ( .A1(n1729), .A2(\inq_ary[4][105] ), .A3(n1686), .A4(
        \inq_ary[0][105] ), .Y(n365) );
  AO22X1_RVT U420 ( .A1(n1740), .A2(\inq_ary[12][105] ), .A3(n1751), .A4(
        \inq_ary[9][105] ), .Y(n364) );
  AO22X1_RVT U421 ( .A1(n1739), .A2(\inq_ary[2][105] ), .A3(n1750), .A4(
        \inq_ary[11][105] ), .Y(n363) );
  AO22X1_RVT U422 ( .A1(n1612), .A2(\inq_ary[8][105] ), .A3(n1748), .A4(
        \inq_ary[10][105] ), .Y(n362) );
  NOR4X1_RVT U423 ( .A1(n365), .A2(n364), .A3(n363), .A4(n362), .Y(n371) );
  AO22X1_RVT U424 ( .A1(n1554), .A2(\inq_ary[14][105] ), .A3(n1711), .A4(
        \inq_ary[13][105] ), .Y(n369) );
  AO22X1_RVT U425 ( .A1(n1537), .A2(\inq_ary[15][105] ), .A3(n1747), .A4(
        \inq_ary[5][105] ), .Y(n368) );
  AO22X1_RVT U426 ( .A1(n1741), .A2(\inq_ary[7][105] ), .A3(n1738), .A4(
        \inq_ary[6][105] ), .Y(n367) );
  AO22X1_RVT U427 ( .A1(n1742), .A2(\inq_ary[3][105] ), .A3(n1749), .A4(
        \inq_ary[1][105] ), .Y(n366) );
  NOR4X1_RVT U428 ( .A1(n369), .A2(n368), .A3(n367), .A4(n366), .Y(n370) );
  NAND2X0_RVT U429 ( .A1(n371), .A2(n370), .Y(n372) );
  AO22X1_RVT U430 ( .A1(n3), .A2(wrdata_d1[105]), .A3(n1), .A4(n372), .Y(n3435) );
  AO22X1_RVT U431 ( .A1(n1686), .A2(\inq_ary[0][37] ), .A3(n1537), .A4(
        \inq_ary[15][37] ), .Y(n376) );
  AO22X1_RVT U432 ( .A1(n1740), .A2(\inq_ary[12][37] ), .A3(n1750), .A4(
        \inq_ary[11][37] ), .Y(n375) );
  AO22X1_RVT U433 ( .A1(n1741), .A2(\inq_ary[7][37] ), .A3(n1748), .A4(
        \inq_ary[10][37] ), .Y(n374) );
  AO22X1_RVT U434 ( .A1(n1612), .A2(\inq_ary[8][37] ), .A3(n1751), .A4(
        \inq_ary[9][37] ), .Y(n373) );
  NOR4X1_RVT U435 ( .A1(n376), .A2(n375), .A3(n374), .A4(n373), .Y(n382) );
  AO22X1_RVT U436 ( .A1(n1738), .A2(\inq_ary[6][37] ), .A3(n1711), .A4(
        \inq_ary[13][37] ), .Y(n380) );
  AO22X1_RVT U437 ( .A1(n1739), .A2(\inq_ary[2][37] ), .A3(n1554), .A4(
        \inq_ary[14][37] ), .Y(n379) );
  AO22X1_RVT U438 ( .A1(n1729), .A2(\inq_ary[4][37] ), .A3(n1749), .A4(
        \inq_ary[1][37] ), .Y(n378) );
  AO22X1_RVT U439 ( .A1(n1742), .A2(\inq_ary[3][37] ), .A3(n1747), .A4(
        \inq_ary[5][37] ), .Y(n377) );
  NOR4X1_RVT U440 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .Y(n381) );
  NAND2X0_RVT U441 ( .A1(n382), .A2(n381), .Y(n383) );
  AO22X1_RVT U442 ( .A1(n1723), .A2(wrdata_d1[37]), .A3(n2), .A4(n383), .Y(
        n3369) );
  AO22X1_RVT U443 ( .A1(n1729), .A2(\inq_ary[4][38] ), .A3(n1738), .A4(
        \inq_ary[6][38] ), .Y(n387) );
  AO22X1_RVT U444 ( .A1(n1742), .A2(\inq_ary[3][38] ), .A3(n1751), .A4(
        \inq_ary[9][38] ), .Y(n386) );
  AO22X1_RVT U445 ( .A1(n1686), .A2(\inq_ary[0][38] ), .A3(n1612), .A4(
        \inq_ary[8][38] ), .Y(n385) );
  AO22X1_RVT U446 ( .A1(n1739), .A2(\inq_ary[2][38] ), .A3(n1740), .A4(
        \inq_ary[12][38] ), .Y(n384) );
  NOR4X1_RVT U447 ( .A1(n387), .A2(n386), .A3(n385), .A4(n384), .Y(n393) );
  AO22X1_RVT U448 ( .A1(n1537), .A2(\inq_ary[15][38] ), .A3(n1749), .A4(
        \inq_ary[1][38] ), .Y(n391) );
  AO22X1_RVT U449 ( .A1(n1750), .A2(\inq_ary[11][38] ), .A3(n1748), .A4(
        \inq_ary[10][38] ), .Y(n390) );
  AO22X1_RVT U450 ( .A1(n1554), .A2(\inq_ary[14][38] ), .A3(n1741), .A4(
        \inq_ary[7][38] ), .Y(n389) );
  AO22X1_RVT U451 ( .A1(n1747), .A2(\inq_ary[5][38] ), .A3(n1711), .A4(
        \inq_ary[13][38] ), .Y(n388) );
  NOR4X1_RVT U452 ( .A1(n391), .A2(n390), .A3(n389), .A4(n388), .Y(n392) );
  NAND2X0_RVT U453 ( .A1(n393), .A2(n392), .Y(n394) );
  AO22X1_RVT U454 ( .A1(n1760), .A2(wrdata_d1[38]), .A3(n2), .A4(n394), .Y(
        n3371) );
  AO22X1_RVT U455 ( .A1(n1612), .A2(\inq_ary[8][106] ), .A3(n1747), .A4(
        \inq_ary[5][106] ), .Y(n398) );
  AO22X1_RVT U456 ( .A1(n1739), .A2(\inq_ary[2][106] ), .A3(n1537), .A4(
        \inq_ary[15][106] ), .Y(n397) );
  AO22X1_RVT U457 ( .A1(n1742), .A2(\inq_ary[3][106] ), .A3(n1738), .A4(
        \inq_ary[6][106] ), .Y(n396) );
  AO22X1_RVT U458 ( .A1(n1750), .A2(\inq_ary[11][106] ), .A3(n1748), .A4(
        \inq_ary[10][106] ), .Y(n395) );
  NOR4X1_RVT U459 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .Y(n404) );
  AO22X1_RVT U460 ( .A1(n1686), .A2(\inq_ary[0][106] ), .A3(n1751), .A4(
        \inq_ary[9][106] ), .Y(n402) );
  AO22X1_RVT U461 ( .A1(n1554), .A2(\inq_ary[14][106] ), .A3(n1729), .A4(
        \inq_ary[4][106] ), .Y(n401) );
  AO22X1_RVT U462 ( .A1(n1740), .A2(\inq_ary[12][106] ), .A3(n1741), .A4(
        \inq_ary[7][106] ), .Y(n400) );
  AO22X1_RVT U463 ( .A1(n1749), .A2(\inq_ary[1][106] ), .A3(n1711), .A4(
        \inq_ary[13][106] ), .Y(n399) );
  NOR4X1_RVT U464 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .Y(n403) );
  NAND2X0_RVT U465 ( .A1(n404), .A2(n403), .Y(n405) );
  AO22X1_RVT U466 ( .A1(n758), .A2(wrdata_d1[106]), .A3(n1), .A4(n405), .Y(
        n3437) );
  AO22X1_RVT U467 ( .A1(n1742), .A2(\inq_ary[3][107] ), .A3(n1750), .A4(
        \inq_ary[11][107] ), .Y(n409) );
  AO22X1_RVT U468 ( .A1(n1612), .A2(\inq_ary[8][107] ), .A3(n1747), .A4(
        \inq_ary[5][107] ), .Y(n408) );
  AO22X1_RVT U469 ( .A1(n1686), .A2(\inq_ary[0][107] ), .A3(n1537), .A4(
        \inq_ary[15][107] ), .Y(n407) );
  AO22X1_RVT U470 ( .A1(n1739), .A2(\inq_ary[2][107] ), .A3(n1711), .A4(
        \inq_ary[13][107] ), .Y(n406) );
  NOR4X1_RVT U471 ( .A1(n409), .A2(n408), .A3(n407), .A4(n406), .Y(n415) );
  AO22X1_RVT U472 ( .A1(n1554), .A2(\inq_ary[14][107] ), .A3(n1751), .A4(
        \inq_ary[9][107] ), .Y(n413) );
  AO22X1_RVT U473 ( .A1(n1741), .A2(\inq_ary[7][107] ), .A3(n1738), .A4(
        \inq_ary[6][107] ), .Y(n412) );
  AO22X1_RVT U474 ( .A1(n1740), .A2(\inq_ary[12][107] ), .A3(n1748), .A4(
        \inq_ary[10][107] ), .Y(n411) );
  AO22X1_RVT U475 ( .A1(n1729), .A2(\inq_ary[4][107] ), .A3(n1749), .A4(
        \inq_ary[1][107] ), .Y(n410) );
  NOR4X1_RVT U476 ( .A1(n413), .A2(n412), .A3(n411), .A4(n410), .Y(n414) );
  NAND2X0_RVT U477 ( .A1(n415), .A2(n414), .Y(n416) );
  AO22X1_RVT U478 ( .A1(n1477), .A2(wrdata_d1[107]), .A3(n1), .A4(n416), .Y(
        n3439) );
  AO22X1_RVT U479 ( .A1(n1742), .A2(\inq_ary[3][36] ), .A3(n1749), .A4(
        \inq_ary[1][36] ), .Y(n420) );
  AO22X1_RVT U480 ( .A1(n1729), .A2(\inq_ary[4][36] ), .A3(n1711), .A4(
        \inq_ary[13][36] ), .Y(n419) );
  AO22X1_RVT U481 ( .A1(n1554), .A2(\inq_ary[14][36] ), .A3(n1751), .A4(
        \inq_ary[9][36] ), .Y(n418) );
  AO22X1_RVT U482 ( .A1(n1747), .A2(\inq_ary[5][36] ), .A3(n1748), .A4(
        \inq_ary[10][36] ), .Y(n417) );
  NOR4X1_RVT U483 ( .A1(n420), .A2(n419), .A3(n418), .A4(n417), .Y(n426) );
  AO22X1_RVT U484 ( .A1(n1739), .A2(\inq_ary[2][36] ), .A3(n1750), .A4(
        \inq_ary[11][36] ), .Y(n424) );
  AO22X1_RVT U485 ( .A1(n1686), .A2(\inq_ary[0][36] ), .A3(n1740), .A4(
        \inq_ary[12][36] ), .Y(n423) );
  AO22X1_RVT U486 ( .A1(n1612), .A2(\inq_ary[8][36] ), .A3(n1738), .A4(
        \inq_ary[6][36] ), .Y(n422) );
  AO22X1_RVT U487 ( .A1(n1537), .A2(\inq_ary[15][36] ), .A3(n1741), .A4(
        \inq_ary[7][36] ), .Y(n421) );
  NOR4X1_RVT U488 ( .A1(n424), .A2(n423), .A3(n422), .A4(n421), .Y(n425) );
  NAND2X0_RVT U489 ( .A1(n426), .A2(n425), .Y(n427) );
  AO22X1_RVT U490 ( .A1(n1477), .A2(wrdata_d1[36]), .A3(n2), .A4(n427), .Y(
        n3367) );
  AO22X1_RVT U491 ( .A1(n1686), .A2(\inq_ary[0][108] ), .A3(n1741), .A4(
        \inq_ary[7][108] ), .Y(n431) );
  AO22X1_RVT U492 ( .A1(n1747), .A2(\inq_ary[5][108] ), .A3(n1738), .A4(
        \inq_ary[6][108] ), .Y(n430) );
  AO22X1_RVT U493 ( .A1(n1742), .A2(\inq_ary[3][108] ), .A3(n1748), .A4(
        \inq_ary[10][108] ), .Y(n429) );
  AO22X1_RVT U494 ( .A1(n1740), .A2(\inq_ary[12][108] ), .A3(n1749), .A4(
        \inq_ary[1][108] ), .Y(n428) );
  NOR4X1_RVT U495 ( .A1(n431), .A2(n430), .A3(n429), .A4(n428), .Y(n437) );
  AO22X1_RVT U496 ( .A1(n1750), .A2(\inq_ary[11][108] ), .A3(n1751), .A4(
        \inq_ary[9][108] ), .Y(n435) );
  AO22X1_RVT U497 ( .A1(n1729), .A2(\inq_ary[4][108] ), .A3(n1612), .A4(
        \inq_ary[8][108] ), .Y(n434) );
  AO22X1_RVT U498 ( .A1(n1554), .A2(\inq_ary[14][108] ), .A3(n1537), .A4(
        \inq_ary[15][108] ), .Y(n433) );
  AO22X1_RVT U499 ( .A1(n1739), .A2(\inq_ary[2][108] ), .A3(n1711), .A4(
        \inq_ary[13][108] ), .Y(n432) );
  NOR4X1_RVT U500 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .Y(n436) );
  NAND2X0_RVT U501 ( .A1(n437), .A2(n436), .Y(n438) );
  AO22X1_RVT U502 ( .A1(n1025), .A2(wrdata_d1[108]), .A3(n1), .A4(n438), .Y(
        n3432) );
  AO22X1_RVT U503 ( .A1(n1741), .A2(\inq_ary[7][109] ), .A3(n1748), .A4(
        \inq_ary[10][109] ), .Y(n442) );
  AO22X1_RVT U504 ( .A1(n1742), .A2(\inq_ary[3][109] ), .A3(n1612), .A4(
        \inq_ary[8][109] ), .Y(n441) );
  AO22X1_RVT U505 ( .A1(n1739), .A2(\inq_ary[2][109] ), .A3(n1751), .A4(
        \inq_ary[9][109] ), .Y(n440) );
  AO22X1_RVT U506 ( .A1(n1537), .A2(\inq_ary[15][109] ), .A3(n1747), .A4(
        \inq_ary[5][109] ), .Y(n439) );
  NOR4X1_RVT U507 ( .A1(n442), .A2(n441), .A3(n440), .A4(n439), .Y(n448) );
  AO22X1_RVT U508 ( .A1(n1554), .A2(\inq_ary[14][109] ), .A3(n1686), .A4(
        \inq_ary[0][109] ), .Y(n446) );
  AO22X1_RVT U509 ( .A1(n1740), .A2(\inq_ary[12][109] ), .A3(n1749), .A4(
        \inq_ary[1][109] ), .Y(n445) );
  AO22X1_RVT U510 ( .A1(n1750), .A2(\inq_ary[11][109] ), .A3(n1711), .A4(
        \inq_ary[13][109] ), .Y(n444) );
  AO22X1_RVT U511 ( .A1(n1729), .A2(\inq_ary[4][109] ), .A3(n1738), .A4(
        \inq_ary[6][109] ), .Y(n443) );
  NOR4X1_RVT U512 ( .A1(n446), .A2(n445), .A3(n444), .A4(n443), .Y(n447) );
  NAND2X0_RVT U513 ( .A1(n448), .A2(n447), .Y(n449) );
  AO22X1_RVT U514 ( .A1(n1477), .A2(wrdata_d1[109]), .A3(n1), .A4(n449), .Y(
        n3434) );
  AO22X1_RVT U515 ( .A1(n1686), .A2(\inq_ary[0][35] ), .A3(n1750), .A4(
        \inq_ary[11][35] ), .Y(n453) );
  AO22X1_RVT U516 ( .A1(n1729), .A2(\inq_ary[4][35] ), .A3(n1738), .A4(
        \inq_ary[6][35] ), .Y(n452) );
  AO22X1_RVT U517 ( .A1(n1537), .A2(\inq_ary[15][35] ), .A3(n1749), .A4(
        \inq_ary[1][35] ), .Y(n451) );
  AO22X1_RVT U518 ( .A1(n1612), .A2(\inq_ary[8][35] ), .A3(n1747), .A4(
        \inq_ary[5][35] ), .Y(n450) );
  NOR4X1_RVT U519 ( .A1(n453), .A2(n452), .A3(n451), .A4(n450), .Y(n459) );
  AO22X1_RVT U520 ( .A1(n1739), .A2(\inq_ary[2][35] ), .A3(n1711), .A4(
        \inq_ary[13][35] ), .Y(n457) );
  AO22X1_RVT U521 ( .A1(n1742), .A2(\inq_ary[3][35] ), .A3(n1751), .A4(
        \inq_ary[9][35] ), .Y(n456) );
  AO22X1_RVT U522 ( .A1(n1554), .A2(\inq_ary[14][35] ), .A3(n1740), .A4(
        \inq_ary[12][35] ), .Y(n455) );
  AO22X1_RVT U523 ( .A1(n1741), .A2(\inq_ary[7][35] ), .A3(n1748), .A4(
        \inq_ary[10][35] ), .Y(n454) );
  NOR4X1_RVT U524 ( .A1(n457), .A2(n456), .A3(n455), .A4(n454), .Y(n458) );
  NAND2X0_RVT U525 ( .A1(n459), .A2(n458), .Y(n460) );
  AO22X1_RVT U526 ( .A1(n1684), .A2(wrdata_d1[35]), .A3(n2), .A4(n460), .Y(
        n3374) );
  AO22X1_RVT U527 ( .A1(n1554), .A2(\inq_ary[14][68] ), .A3(n1747), .A4(
        \inq_ary[5][68] ), .Y(n464) );
  AO22X1_RVT U528 ( .A1(n1612), .A2(\inq_ary[8][68] ), .A3(n1750), .A4(
        \inq_ary[11][68] ), .Y(n463) );
  AO22X1_RVT U529 ( .A1(n1729), .A2(\inq_ary[4][68] ), .A3(n1537), .A4(
        \inq_ary[15][68] ), .Y(n462) );
  AO22X1_RVT U530 ( .A1(n1739), .A2(\inq_ary[2][68] ), .A3(n1751), .A4(
        \inq_ary[9][68] ), .Y(n461) );
  NOR4X1_RVT U531 ( .A1(n464), .A2(n463), .A3(n462), .A4(n461), .Y(n470) );
  AO22X1_RVT U532 ( .A1(n1686), .A2(\inq_ary[0][68] ), .A3(n1741), .A4(
        \inq_ary[7][68] ), .Y(n468) );
  AO22X1_RVT U533 ( .A1(n1749), .A2(\inq_ary[1][68] ), .A3(n1748), .A4(
        \inq_ary[10][68] ), .Y(n467) );
  AO22X1_RVT U534 ( .A1(n1740), .A2(\inq_ary[12][68] ), .A3(n1711), .A4(
        \inq_ary[13][68] ), .Y(n466) );
  AO22X1_RVT U535 ( .A1(n1742), .A2(\inq_ary[3][68] ), .A3(n1738), .A4(
        \inq_ary[6][68] ), .Y(n465) );
  NOR4X1_RVT U536 ( .A1(n468), .A2(n467), .A3(n466), .A4(n465), .Y(n469) );
  NAND2X0_RVT U537 ( .A1(n470), .A2(n469), .Y(n471) );
  AO22X1_RVT U538 ( .A1(n3), .A2(wrdata_d1[68]), .A3(n1), .A4(n471), .Y(n3392)
         );
  AO22X1_RVT U539 ( .A1(n1554), .A2(\inq_ary[14][69] ), .A3(n1748), .A4(
        \inq_ary[10][69] ), .Y(n475) );
  AO22X1_RVT U540 ( .A1(n1742), .A2(\inq_ary[3][69] ), .A3(n1711), .A4(
        \inq_ary[13][69] ), .Y(n474) );
  AO22X1_RVT U541 ( .A1(n1612), .A2(\inq_ary[8][69] ), .A3(n1738), .A4(
        \inq_ary[6][69] ), .Y(n473) );
  AO22X1_RVT U542 ( .A1(n1739), .A2(\inq_ary[2][69] ), .A3(n1750), .A4(
        \inq_ary[11][69] ), .Y(n472) );
  NOR4X1_RVT U543 ( .A1(n475), .A2(n474), .A3(n473), .A4(n472), .Y(n481) );
  AO22X1_RVT U544 ( .A1(n1740), .A2(\inq_ary[12][69] ), .A3(n1751), .A4(
        \inq_ary[9][69] ), .Y(n479) );
  AO22X1_RVT U545 ( .A1(n1749), .A2(\inq_ary[1][69] ), .A3(n1741), .A4(
        \inq_ary[7][69] ), .Y(n478) );
  AO22X1_RVT U546 ( .A1(n1686), .A2(\inq_ary[0][69] ), .A3(n1537), .A4(
        \inq_ary[15][69] ), .Y(n477) );
  AO22X1_RVT U547 ( .A1(n1729), .A2(\inq_ary[4][69] ), .A3(n1747), .A4(
        \inq_ary[5][69] ), .Y(n476) );
  NOR4X1_RVT U548 ( .A1(n479), .A2(n478), .A3(n477), .A4(n476), .Y(n480) );
  NAND2X0_RVT U549 ( .A1(n481), .A2(n480), .Y(n482) );
  AO22X1_RVT U550 ( .A1(n3), .A2(wrdata_d1[69]), .A3(n1489), .A4(n482), .Y(
        n3394) );
  AO22X1_RVT U551 ( .A1(n1729), .A2(\inq_ary[4][55] ), .A3(n1740), .A4(
        \inq_ary[12][55] ), .Y(n486) );
  AO22X1_RVT U552 ( .A1(n1612), .A2(\inq_ary[8][55] ), .A3(n1749), .A4(
        \inq_ary[1][55] ), .Y(n485) );
  AO22X1_RVT U553 ( .A1(n1739), .A2(\inq_ary[2][55] ), .A3(n1751), .A4(
        \inq_ary[9][55] ), .Y(n484) );
  AO22X1_RVT U554 ( .A1(n1741), .A2(\inq_ary[7][55] ), .A3(n1711), .A4(
        \inq_ary[13][55] ), .Y(n483) );
  NOR4X1_RVT U555 ( .A1(n486), .A2(n485), .A3(n484), .A4(n483), .Y(n492) );
  AO22X1_RVT U556 ( .A1(n1750), .A2(\inq_ary[11][55] ), .A3(n1748), .A4(
        \inq_ary[10][55] ), .Y(n490) );
  AO22X1_RVT U557 ( .A1(n1554), .A2(\inq_ary[14][55] ), .A3(n1686), .A4(
        \inq_ary[0][55] ), .Y(n489) );
  AO22X1_RVT U558 ( .A1(n1742), .A2(\inq_ary[3][55] ), .A3(n1537), .A4(
        \inq_ary[15][55] ), .Y(n488) );
  AO22X1_RVT U559 ( .A1(n1747), .A2(\inq_ary[5][55] ), .A3(n1738), .A4(
        \inq_ary[6][55] ), .Y(n487) );
  NOR4X1_RVT U560 ( .A1(n490), .A2(n489), .A3(n488), .A4(n487), .Y(n491) );
  NAND2X0_RVT U561 ( .A1(n492), .A2(n491), .Y(n493) );
  AO22X1_RVT U562 ( .A1(n1598), .A2(wrdata_d1[55]), .A3(n1759), .A4(n493), .Y(
        n3388) );
  AO22X1_RVT U563 ( .A1(n1742), .A2(\inq_ary[3][70] ), .A3(n1741), .A4(
        \inq_ary[7][70] ), .Y(n497) );
  AO22X1_RVT U564 ( .A1(n1749), .A2(\inq_ary[1][70] ), .A3(n1748), .A4(
        \inq_ary[10][70] ), .Y(n496) );
  AO22X1_RVT U565 ( .A1(n1554), .A2(\inq_ary[14][70] ), .A3(n1750), .A4(
        \inq_ary[11][70] ), .Y(n495) );
  AO22X1_RVT U566 ( .A1(n1612), .A2(\inq_ary[8][70] ), .A3(n1751), .A4(
        \inq_ary[9][70] ), .Y(n494) );
  NOR4X1_RVT U567 ( .A1(n497), .A2(n496), .A3(n495), .A4(n494), .Y(n503) );
  AO22X1_RVT U568 ( .A1(n1738), .A2(\inq_ary[6][70] ), .A3(n1711), .A4(
        \inq_ary[13][70] ), .Y(n501) );
  AO22X1_RVT U569 ( .A1(n1729), .A2(\inq_ary[4][70] ), .A3(n1740), .A4(
        \inq_ary[12][70] ), .Y(n500) );
  AO22X1_RVT U570 ( .A1(n1686), .A2(\inq_ary[0][70] ), .A3(n1537), .A4(
        \inq_ary[15][70] ), .Y(n499) );
  AO22X1_RVT U571 ( .A1(n1739), .A2(\inq_ary[2][70] ), .A3(n1747), .A4(
        \inq_ary[5][70] ), .Y(n498) );
  NOR4X1_RVT U572 ( .A1(n501), .A2(n500), .A3(n499), .A4(n498), .Y(n502) );
  NAND2X0_RVT U573 ( .A1(n503), .A2(n502), .Y(n504) );
  AO22X1_RVT U574 ( .A1(n3), .A2(wrdata_d1[70]), .A3(n1), .A4(n504), .Y(n3396)
         );
  AO22X1_RVT U575 ( .A1(n1742), .A2(\inq_ary[3][71] ), .A3(n1711), .A4(
        \inq_ary[13][71] ), .Y(n508) );
  AO22X1_RVT U576 ( .A1(n1729), .A2(\inq_ary[4][71] ), .A3(n1738), .A4(
        \inq_ary[6][71] ), .Y(n507) );
  AO22X1_RVT U577 ( .A1(n1739), .A2(\inq_ary[2][71] ), .A3(n1740), .A4(
        \inq_ary[12][71] ), .Y(n506) );
  AO22X1_RVT U578 ( .A1(n1554), .A2(\inq_ary[14][71] ), .A3(n1747), .A4(
        \inq_ary[5][71] ), .Y(n505) );
  NOR4X1_RVT U579 ( .A1(n508), .A2(n507), .A3(n506), .A4(n505), .Y(n514) );
  AO22X1_RVT U580 ( .A1(n1750), .A2(\inq_ary[11][71] ), .A3(n1751), .A4(
        \inq_ary[9][71] ), .Y(n512) );
  AO22X1_RVT U581 ( .A1(n1537), .A2(\inq_ary[15][71] ), .A3(n1612), .A4(
        \inq_ary[8][71] ), .Y(n511) );
  AO22X1_RVT U582 ( .A1(n1749), .A2(\inq_ary[1][71] ), .A3(n1748), .A4(
        \inq_ary[10][71] ), .Y(n510) );
  AO22X1_RVT U583 ( .A1(n1686), .A2(\inq_ary[0][71] ), .A3(n1741), .A4(
        \inq_ary[7][71] ), .Y(n509) );
  NOR4X1_RVT U584 ( .A1(n512), .A2(n511), .A3(n510), .A4(n509), .Y(n513) );
  NAND2X0_RVT U585 ( .A1(n514), .A2(n513), .Y(n515) );
  AO22X1_RVT U586 ( .A1(n1723), .A2(wrdata_d1[71]), .A3(n1), .A4(n515), .Y(
        n3398) );
  AO22X1_RVT U587 ( .A1(n1537), .A2(\inq_ary[15][54] ), .A3(n1740), .A4(
        \inq_ary[12][54] ), .Y(n519) );
  AO22X1_RVT U588 ( .A1(n1686), .A2(\inq_ary[0][54] ), .A3(n1741), .A4(
        \inq_ary[7][54] ), .Y(n518) );
  AO22X1_RVT U589 ( .A1(n1742), .A2(\inq_ary[3][54] ), .A3(n1612), .A4(
        \inq_ary[8][54] ), .Y(n517) );
  AO22X1_RVT U590 ( .A1(n1750), .A2(\inq_ary[11][54] ), .A3(n1711), .A4(
        \inq_ary[13][54] ), .Y(n516) );
  NOR4X1_RVT U591 ( .A1(n519), .A2(n518), .A3(n517), .A4(n516), .Y(n525) );
  AO22X1_RVT U592 ( .A1(n1554), .A2(\inq_ary[14][54] ), .A3(n1729), .A4(
        \inq_ary[4][54] ), .Y(n523) );
  AO22X1_RVT U593 ( .A1(n1738), .A2(\inq_ary[6][54] ), .A3(n1748), .A4(
        \inq_ary[10][54] ), .Y(n522) );
  AO22X1_RVT U594 ( .A1(n1739), .A2(\inq_ary[2][54] ), .A3(n1747), .A4(
        \inq_ary[5][54] ), .Y(n521) );
  AO22X1_RVT U595 ( .A1(n1749), .A2(\inq_ary[1][54] ), .A3(n1751), .A4(
        \inq_ary[9][54] ), .Y(n520) );
  NOR4X1_RVT U596 ( .A1(n523), .A2(n522), .A3(n521), .A4(n520), .Y(n524) );
  NAND2X0_RVT U597 ( .A1(n525), .A2(n524), .Y(n526) );
  AO22X1_RVT U598 ( .A1(n1723), .A2(wrdata_d1[54]), .A3(n1), .A4(n526), .Y(
        n3386) );
  AO22X1_RVT U599 ( .A1(n1750), .A2(\inq_ary[11][72] ), .A3(n1748), .A4(
        \inq_ary[10][72] ), .Y(n530) );
  AO22X1_RVT U600 ( .A1(n1554), .A2(\inq_ary[14][72] ), .A3(n1729), .A4(
        \inq_ary[4][72] ), .Y(n529) );
  AO22X1_RVT U601 ( .A1(n1711), .A2(\inq_ary[13][72] ), .A3(n1751), .A4(
        \inq_ary[9][72] ), .Y(n528) );
  AO22X1_RVT U602 ( .A1(n1612), .A2(\inq_ary[8][72] ), .A3(n1741), .A4(
        \inq_ary[7][72] ), .Y(n527) );
  NOR4X1_RVT U603 ( .A1(n530), .A2(n529), .A3(n528), .A4(n527), .Y(n536) );
  AO22X1_RVT U604 ( .A1(n1537), .A2(\inq_ary[15][72] ), .A3(n1749), .A4(
        \inq_ary[1][72] ), .Y(n534) );
  AO22X1_RVT U605 ( .A1(n1747), .A2(\inq_ary[5][72] ), .A3(n1738), .A4(
        \inq_ary[6][72] ), .Y(n533) );
  AO22X1_RVT U606 ( .A1(n1739), .A2(\inq_ary[2][72] ), .A3(n1742), .A4(
        \inq_ary[3][72] ), .Y(n532) );
  AO22X1_RVT U607 ( .A1(n1686), .A2(\inq_ary[0][72] ), .A3(n1740), .A4(
        \inq_ary[12][72] ), .Y(n531) );
  NOR4X1_RVT U608 ( .A1(n534), .A2(n533), .A3(n532), .A4(n531), .Y(n535) );
  NAND2X0_RVT U609 ( .A1(n536), .A2(n535), .Y(n537) );
  AO22X1_RVT U610 ( .A1(n3), .A2(wrdata_d1[72]), .A3(n1759), .A4(n537), .Y(
        n3401) );
  AO22X1_RVT U611 ( .A1(n1747), .A2(\inq_ary[5][73] ), .A3(n1750), .A4(
        \inq_ary[11][73] ), .Y(n541) );
  AO22X1_RVT U612 ( .A1(n1739), .A2(\inq_ary[2][73] ), .A3(n1742), .A4(
        \inq_ary[3][73] ), .Y(n540) );
  AO22X1_RVT U613 ( .A1(n1554), .A2(\inq_ary[14][73] ), .A3(n1748), .A4(
        \inq_ary[10][73] ), .Y(n539) );
  AO22X1_RVT U614 ( .A1(n1686), .A2(\inq_ary[0][73] ), .A3(n1749), .A4(
        \inq_ary[1][73] ), .Y(n538) );
  NOR4X1_RVT U615 ( .A1(n541), .A2(n540), .A3(n539), .A4(n538), .Y(n547) );
  AO22X1_RVT U616 ( .A1(n1729), .A2(\inq_ary[4][73] ), .A3(n1612), .A4(
        \inq_ary[8][73] ), .Y(n545) );
  AO22X1_RVT U617 ( .A1(n1738), .A2(\inq_ary[6][73] ), .A3(n1751), .A4(
        \inq_ary[9][73] ), .Y(n544) );
  AO22X1_RVT U618 ( .A1(n1740), .A2(\inq_ary[12][73] ), .A3(n1711), .A4(
        \inq_ary[13][73] ), .Y(n543) );
  AO22X1_RVT U619 ( .A1(n1537), .A2(\inq_ary[15][73] ), .A3(n1741), .A4(
        \inq_ary[7][73] ), .Y(n542) );
  NOR4X1_RVT U620 ( .A1(n545), .A2(n544), .A3(n543), .A4(n542), .Y(n546) );
  NAND2X0_RVT U621 ( .A1(n547), .A2(n546), .Y(n548) );
  AO22X1_RVT U622 ( .A1(n3), .A2(wrdata_d1[73]), .A3(n946), .A4(n548), .Y(
        n3403) );
  AO22X1_RVT U623 ( .A1(n1729), .A2(\inq_ary[4][53] ), .A3(n1747), .A4(
        \inq_ary[5][53] ), .Y(n552) );
  AO22X1_RVT U624 ( .A1(n1686), .A2(\inq_ary[0][53] ), .A3(n1537), .A4(
        \inq_ary[15][53] ), .Y(n551) );
  AO22X1_RVT U625 ( .A1(n1741), .A2(\inq_ary[7][53] ), .A3(n1750), .A4(
        \inq_ary[11][53] ), .Y(n550) );
  AO22X1_RVT U626 ( .A1(n1612), .A2(\inq_ary[8][53] ), .A3(n1740), .A4(
        \inq_ary[12][53] ), .Y(n549) );
  NOR4X1_RVT U627 ( .A1(n552), .A2(n551), .A3(n550), .A4(n549), .Y(n558) );
  AO22X1_RVT U628 ( .A1(n1711), .A2(\inq_ary[13][53] ), .A3(n1748), .A4(
        \inq_ary[10][53] ), .Y(n556) );
  AO22X1_RVT U629 ( .A1(n1554), .A2(\inq_ary[14][53] ), .A3(n1749), .A4(
        \inq_ary[1][53] ), .Y(n555) );
  AO22X1_RVT U630 ( .A1(n1742), .A2(\inq_ary[3][53] ), .A3(n1738), .A4(
        \inq_ary[6][53] ), .Y(n554) );
  AO22X1_RVT U631 ( .A1(n1739), .A2(\inq_ary[2][53] ), .A3(n1751), .A4(
        \inq_ary[9][53] ), .Y(n553) );
  NOR4X1_RVT U632 ( .A1(n556), .A2(n555), .A3(n554), .A4(n553), .Y(n557) );
  NAND2X0_RVT U633 ( .A1(n558), .A2(n557), .Y(n559) );
  AO22X1_RVT U634 ( .A1(n758), .A2(wrdata_d1[53]), .A3(n1), .A4(n559), .Y(
        n3384) );
  AO22X1_RVT U635 ( .A1(n1742), .A2(\inq_ary[3][61] ), .A3(n1741), .A4(
        \inq_ary[7][61] ), .Y(n563) );
  AO22X1_RVT U636 ( .A1(n1537), .A2(\inq_ary[15][61] ), .A3(n1738), .A4(
        \inq_ary[6][61] ), .Y(n562) );
  AO22X1_RVT U637 ( .A1(n1739), .A2(\inq_ary[2][61] ), .A3(n1686), .A4(
        \inq_ary[0][61] ), .Y(n561) );
  AO22X1_RVT U638 ( .A1(n1749), .A2(\inq_ary[1][61] ), .A3(n1711), .A4(
        \inq_ary[13][61] ), .Y(n560) );
  NOR4X1_RVT U639 ( .A1(n563), .A2(n562), .A3(n561), .A4(n560), .Y(n569) );
  AO22X1_RVT U640 ( .A1(n1747), .A2(\inq_ary[5][61] ), .A3(n1751), .A4(
        \inq_ary[9][61] ), .Y(n567) );
  AO22X1_RVT U641 ( .A1(n1750), .A2(\inq_ary[11][61] ), .A3(n1748), .A4(
        \inq_ary[10][61] ), .Y(n566) );
  AO22X1_RVT U642 ( .A1(n1729), .A2(\inq_ary[4][61] ), .A3(n1612), .A4(
        \inq_ary[8][61] ), .Y(n565) );
  AO22X1_RVT U643 ( .A1(n1554), .A2(\inq_ary[14][61] ), .A3(n1740), .A4(
        \inq_ary[12][61] ), .Y(n564) );
  NOR4X1_RVT U644 ( .A1(n567), .A2(n566), .A3(n565), .A4(n564), .Y(n568) );
  NAND2X0_RVT U645 ( .A1(n569), .A2(n568), .Y(n570) );
  AO22X1_RVT U646 ( .A1(n1684), .A2(wrdata_d1[61]), .A3(n946), .A4(n570), .Y(
        n3391) );
  AO22X1_RVT U647 ( .A1(n1740), .A2(\inq_ary[12][64] ), .A3(n1748), .A4(
        \inq_ary[10][64] ), .Y(n574) );
  AO22X1_RVT U648 ( .A1(n1742), .A2(\inq_ary[3][64] ), .A3(n1729), .A4(
        \inq_ary[4][64] ), .Y(n573) );
  AO22X1_RVT U649 ( .A1(n1738), .A2(\inq_ary[6][64] ), .A3(n1751), .A4(
        \inq_ary[9][64] ), .Y(n572) );
  AO22X1_RVT U650 ( .A1(n1554), .A2(\inq_ary[14][64] ), .A3(n1741), .A4(
        \inq_ary[7][64] ), .Y(n571) );
  NOR4X1_RVT U651 ( .A1(n574), .A2(n573), .A3(n572), .A4(n571), .Y(n580) );
  AO22X1_RVT U652 ( .A1(n1537), .A2(\inq_ary[15][64] ), .A3(n1749), .A4(
        \inq_ary[1][64] ), .Y(n578) );
  AO22X1_RVT U653 ( .A1(n1739), .A2(\inq_ary[2][64] ), .A3(n1686), .A4(
        \inq_ary[0][64] ), .Y(n577) );
  AO22X1_RVT U654 ( .A1(n1612), .A2(\inq_ary[8][64] ), .A3(n1711), .A4(
        \inq_ary[13][64] ), .Y(n576) );
  AO22X1_RVT U655 ( .A1(n1747), .A2(\inq_ary[5][64] ), .A3(n1750), .A4(
        \inq_ary[11][64] ), .Y(n575) );
  NOR4X1_RVT U656 ( .A1(n578), .A2(n577), .A3(n576), .A4(n575), .Y(n579) );
  NAND2X0_RVT U657 ( .A1(n580), .A2(n579), .Y(n581) );
  AO22X1_RVT U658 ( .A1(n3), .A2(wrdata_d1[64]), .A3(n2), .A4(n581), .Y(n3393)
         );
  AO22X1_RVT U659 ( .A1(n1740), .A2(\inq_ary[12][65] ), .A3(n1750), .A4(
        \inq_ary[11][65] ), .Y(n585) );
  AO22X1_RVT U660 ( .A1(n1686), .A2(\inq_ary[0][65] ), .A3(n1749), .A4(
        \inq_ary[1][65] ), .Y(n584) );
  AO22X1_RVT U661 ( .A1(n1554), .A2(\inq_ary[14][65] ), .A3(n1747), .A4(
        \inq_ary[5][65] ), .Y(n583) );
  AO22X1_RVT U662 ( .A1(n1738), .A2(\inq_ary[6][65] ), .A3(n1751), .A4(
        \inq_ary[9][65] ), .Y(n582) );
  NOR4X1_RVT U663 ( .A1(n585), .A2(n584), .A3(n583), .A4(n582), .Y(n591) );
  AO22X1_RVT U664 ( .A1(n1739), .A2(\inq_ary[2][65] ), .A3(n1729), .A4(
        \inq_ary[4][65] ), .Y(n589) );
  AO22X1_RVT U665 ( .A1(n1742), .A2(\inq_ary[3][65] ), .A3(n1612), .A4(
        \inq_ary[8][65] ), .Y(n588) );
  AO22X1_RVT U666 ( .A1(n1537), .A2(\inq_ary[15][65] ), .A3(n1711), .A4(
        \inq_ary[13][65] ), .Y(n587) );
  AO22X1_RVT U667 ( .A1(n1741), .A2(\inq_ary[7][65] ), .A3(n1748), .A4(
        \inq_ary[10][65] ), .Y(n586) );
  NOR4X1_RVT U668 ( .A1(n589), .A2(n588), .A3(n587), .A4(n586), .Y(n590) );
  NAND2X0_RVT U669 ( .A1(n591), .A2(n590), .Y(n592) );
  AO22X1_RVT U670 ( .A1(n1477), .A2(wrdata_d1[65]), .A3(n969), .A4(n592), .Y(
        n3395) );
  AO22X1_RVT U671 ( .A1(n1729), .A2(\inq_ary[4][66] ), .A3(n1749), .A4(
        \inq_ary[1][66] ), .Y(n596) );
  AO22X1_RVT U672 ( .A1(n1739), .A2(\inq_ary[2][66] ), .A3(n1554), .A4(
        \inq_ary[14][66] ), .Y(n595) );
  AO22X1_RVT U673 ( .A1(n1686), .A2(\inq_ary[0][66] ), .A3(n1740), .A4(
        \inq_ary[12][66] ), .Y(n594) );
  AO22X1_RVT U674 ( .A1(n1742), .A2(\inq_ary[3][66] ), .A3(n1748), .A4(
        \inq_ary[10][66] ), .Y(n593) );
  NOR4X1_RVT U675 ( .A1(n596), .A2(n595), .A3(n594), .A4(n593), .Y(n602) );
  AO22X1_RVT U676 ( .A1(n1612), .A2(\inq_ary[8][66] ), .A3(n1741), .A4(
        \inq_ary[7][66] ), .Y(n600) );
  AO22X1_RVT U677 ( .A1(n1750), .A2(\inq_ary[11][66] ), .A3(n1711), .A4(
        \inq_ary[13][66] ), .Y(n599) );
  AO22X1_RVT U678 ( .A1(n1738), .A2(\inq_ary[6][66] ), .A3(n1751), .A4(
        \inq_ary[9][66] ), .Y(n598) );
  AO22X1_RVT U679 ( .A1(n1537), .A2(\inq_ary[15][66] ), .A3(n1747), .A4(
        \inq_ary[5][66] ), .Y(n597) );
  NOR4X1_RVT U680 ( .A1(n600), .A2(n599), .A3(n598), .A4(n597), .Y(n601) );
  NAND2X0_RVT U681 ( .A1(n602), .A2(n601), .Y(n603) );
  AO22X1_RVT U682 ( .A1(n3), .A2(wrdata_d1[66]), .A3(n2), .A4(n603), .Y(n3397)
         );
  AO22X1_RVT U683 ( .A1(n1537), .A2(\inq_ary[15][67] ), .A3(n1748), .A4(
        \inq_ary[10][67] ), .Y(n607) );
  AO22X1_RVT U684 ( .A1(n1740), .A2(\inq_ary[12][67] ), .A3(n1751), .A4(
        \inq_ary[9][67] ), .Y(n606) );
  AO22X1_RVT U685 ( .A1(n1686), .A2(\inq_ary[0][67] ), .A3(n1711), .A4(
        \inq_ary[13][67] ), .Y(n605) );
  AO22X1_RVT U686 ( .A1(n1739), .A2(\inq_ary[2][67] ), .A3(n1749), .A4(
        \inq_ary[1][67] ), .Y(n604) );
  NOR4X1_RVT U687 ( .A1(n607), .A2(n606), .A3(n605), .A4(n604), .Y(n613) );
  AO22X1_RVT U688 ( .A1(n1742), .A2(\inq_ary[3][67] ), .A3(n1729), .A4(
        \inq_ary[4][67] ), .Y(n611) );
  AO22X1_RVT U689 ( .A1(n1612), .A2(\inq_ary[8][67] ), .A3(n1741), .A4(
        \inq_ary[7][67] ), .Y(n610) );
  AO22X1_RVT U690 ( .A1(n1747), .A2(\inq_ary[5][67] ), .A3(n1738), .A4(
        \inq_ary[6][67] ), .Y(n609) );
  AO22X1_RVT U691 ( .A1(n1554), .A2(\inq_ary[14][67] ), .A3(n1750), .A4(
        \inq_ary[11][67] ), .Y(n608) );
  NOR4X1_RVT U692 ( .A1(n611), .A2(n610), .A3(n609), .A4(n608), .Y(n612) );
  NAND2X0_RVT U693 ( .A1(n613), .A2(n612), .Y(n614) );
  AO22X1_RVT U694 ( .A1(n758), .A2(wrdata_d1[67]), .A3(n1489), .A4(n614), .Y(
        n3399) );
  AO22X1_RVT U695 ( .A1(n1738), .A2(\inq_ary[6][82] ), .A3(n1748), .A4(
        \inq_ary[10][82] ), .Y(n618) );
  AO22X1_RVT U696 ( .A1(n1686), .A2(\inq_ary[0][82] ), .A3(n1612), .A4(
        \inq_ary[8][82] ), .Y(n617) );
  AO22X1_RVT U697 ( .A1(n1742), .A2(\inq_ary[3][82] ), .A3(n1750), .A4(
        \inq_ary[11][82] ), .Y(n616) );
  AO22X1_RVT U698 ( .A1(n1739), .A2(\inq_ary[2][82] ), .A3(n1747), .A4(
        \inq_ary[5][82] ), .Y(n615) );
  NOR4X1_RVT U699 ( .A1(n618), .A2(n617), .A3(n616), .A4(n615), .Y(n624) );
  AO22X1_RVT U700 ( .A1(n1554), .A2(\inq_ary[14][82] ), .A3(n1751), .A4(
        \inq_ary[9][82] ), .Y(n622) );
  AO22X1_RVT U701 ( .A1(n1729), .A2(\inq_ary[4][82] ), .A3(n1537), .A4(
        \inq_ary[15][82] ), .Y(n621) );
  AO22X1_RVT U702 ( .A1(n1741), .A2(\inq_ary[7][82] ), .A3(n1711), .A4(
        \inq_ary[13][82] ), .Y(n620) );
  AO22X1_RVT U703 ( .A1(n1740), .A2(\inq_ary[12][82] ), .A3(n1749), .A4(
        \inq_ary[1][82] ), .Y(n619) );
  NOR4X1_RVT U704 ( .A1(n622), .A2(n621), .A3(n620), .A4(n619), .Y(n623) );
  NAND2X0_RVT U705 ( .A1(n624), .A2(n623), .Y(n625) );
  AO22X1_RVT U706 ( .A1(n3), .A2(wrdata_d1[82]), .A3(n969), .A4(n625), .Y(
        n3413) );
  AO22X1_RVT U707 ( .A1(n1747), .A2(\inq_ary[5][83] ), .A3(n1751), .A4(
        \inq_ary[9][83] ), .Y(n629) );
  AO22X1_RVT U708 ( .A1(n1749), .A2(\inq_ary[1][83] ), .A3(n1738), .A4(
        \inq_ary[6][83] ), .Y(n628) );
  AO22X1_RVT U709 ( .A1(n1686), .A2(\inq_ary[0][83] ), .A3(n1612), .A4(
        \inq_ary[8][83] ), .Y(n627) );
  AO22X1_RVT U710 ( .A1(n1729), .A2(\inq_ary[4][83] ), .A3(n1748), .A4(
        \inq_ary[10][83] ), .Y(n626) );
  NOR4X1_RVT U711 ( .A1(n629), .A2(n628), .A3(n627), .A4(n626), .Y(n635) );
  AO22X1_RVT U712 ( .A1(n1742), .A2(\inq_ary[3][83] ), .A3(n1750), .A4(
        \inq_ary[11][83] ), .Y(n633) );
  AO22X1_RVT U713 ( .A1(n1740), .A2(\inq_ary[12][83] ), .A3(n1741), .A4(
        \inq_ary[7][83] ), .Y(n632) );
  AO22X1_RVT U714 ( .A1(n1537), .A2(\inq_ary[15][83] ), .A3(n1711), .A4(
        \inq_ary[13][83] ), .Y(n631) );
  AO22X1_RVT U715 ( .A1(n1739), .A2(\inq_ary[2][83] ), .A3(n1554), .A4(
        \inq_ary[14][83] ), .Y(n630) );
  NOR4X1_RVT U716 ( .A1(n633), .A2(n632), .A3(n631), .A4(n630), .Y(n634) );
  NAND2X0_RVT U717 ( .A1(n635), .A2(n634), .Y(n636) );
  AO22X1_RVT U718 ( .A1(n1477), .A2(wrdata_d1[83]), .A3(n969), .A4(n636), .Y(
        n3415) );
  AO22X1_RVT U719 ( .A1(n1739), .A2(\inq_ary[2][48] ), .A3(n1554), .A4(
        \inq_ary[14][48] ), .Y(n640) );
  AO22X1_RVT U720 ( .A1(n1741), .A2(\inq_ary[7][48] ), .A3(n1711), .A4(
        \inq_ary[13][48] ), .Y(n639) );
  AO22X1_RVT U721 ( .A1(n1747), .A2(\inq_ary[5][48] ), .A3(n1751), .A4(
        \inq_ary[9][48] ), .Y(n638) );
  AO22X1_RVT U722 ( .A1(n1729), .A2(\inq_ary[4][48] ), .A3(n1686), .A4(
        \inq_ary[0][48] ), .Y(n637) );
  NOR4X1_RVT U723 ( .A1(n640), .A2(n639), .A3(n638), .A4(n637), .Y(n646) );
  AO22X1_RVT U724 ( .A1(n1612), .A2(\inq_ary[8][48] ), .A3(n1750), .A4(
        \inq_ary[11][48] ), .Y(n644) );
  AO22X1_RVT U725 ( .A1(n1537), .A2(\inq_ary[15][48] ), .A3(n1749), .A4(
        \inq_ary[1][48] ), .Y(n643) );
  AO22X1_RVT U726 ( .A1(n1740), .A2(\inq_ary[12][48] ), .A3(n1738), .A4(
        \inq_ary[6][48] ), .Y(n642) );
  AO22X1_RVT U727 ( .A1(n1742), .A2(\inq_ary[3][48] ), .A3(n1748), .A4(
        \inq_ary[10][48] ), .Y(n641) );
  NOR4X1_RVT U728 ( .A1(n644), .A2(n643), .A3(n642), .A4(n641), .Y(n645) );
  NAND2X0_RVT U729 ( .A1(n646), .A2(n645), .Y(n647) );
  AO22X1_RVT U730 ( .A1(n1598), .A2(wrdata_d1[48]), .A3(n1759), .A4(n647), .Y(
        n3383) );
  AO22X1_RVT U731 ( .A1(n1750), .A2(\inq_ary[11][84] ), .A3(n1711), .A4(
        \inq_ary[13][84] ), .Y(n651) );
  AO22X1_RVT U732 ( .A1(n1729), .A2(\inq_ary[4][84] ), .A3(n1751), .A4(
        \inq_ary[9][84] ), .Y(n650) );
  AO22X1_RVT U733 ( .A1(n1537), .A2(\inq_ary[15][84] ), .A3(n1748), .A4(
        \inq_ary[10][84] ), .Y(n649) );
  AO22X1_RVT U734 ( .A1(n1612), .A2(\inq_ary[8][84] ), .A3(n1747), .A4(
        \inq_ary[5][84] ), .Y(n648) );
  NOR4X1_RVT U735 ( .A1(n651), .A2(n650), .A3(n649), .A4(n648), .Y(n657) );
  AO22X1_RVT U736 ( .A1(n1554), .A2(\inq_ary[14][84] ), .A3(n1686), .A4(
        \inq_ary[0][84] ), .Y(n655) );
  AO22X1_RVT U737 ( .A1(n1740), .A2(\inq_ary[12][84] ), .A3(n1738), .A4(
        \inq_ary[6][84] ), .Y(n654) );
  AO22X1_RVT U738 ( .A1(n1739), .A2(\inq_ary[2][84] ), .A3(n1749), .A4(
        \inq_ary[1][84] ), .Y(n653) );
  AO22X1_RVT U739 ( .A1(n1742), .A2(\inq_ary[3][84] ), .A3(n1741), .A4(
        \inq_ary[7][84] ), .Y(n652) );
  NOR4X1_RVT U740 ( .A1(n655), .A2(n654), .A3(n653), .A4(n652), .Y(n656) );
  NAND2X0_RVT U741 ( .A1(n657), .A2(n656), .Y(n658) );
  AO22X1_RVT U742 ( .A1(n1723), .A2(wrdata_d1[84]), .A3(n969), .A4(n658), .Y(
        n3408) );
  AO22X1_RVT U743 ( .A1(n1554), .A2(\inq_ary[14][85] ), .A3(n1612), .A4(
        \inq_ary[8][85] ), .Y(n662) );
  AO22X1_RVT U744 ( .A1(n1750), .A2(\inq_ary[11][85] ), .A3(n1711), .A4(
        \inq_ary[13][85] ), .Y(n661) );
  AO22X1_RVT U745 ( .A1(n1729), .A2(\inq_ary[4][85] ), .A3(n1751), .A4(
        \inq_ary[9][85] ), .Y(n660) );
  AO22X1_RVT U746 ( .A1(n1686), .A2(\inq_ary[0][85] ), .A3(n1748), .A4(
        \inq_ary[10][85] ), .Y(n659) );
  NOR4X1_RVT U747 ( .A1(n662), .A2(n661), .A3(n660), .A4(n659), .Y(n668) );
  AO22X1_RVT U748 ( .A1(n1740), .A2(\inq_ary[12][85] ), .A3(n1747), .A4(
        \inq_ary[5][85] ), .Y(n666) );
  AO22X1_RVT U749 ( .A1(n1742), .A2(\inq_ary[3][85] ), .A3(n1738), .A4(
        \inq_ary[6][85] ), .Y(n665) );
  AO22X1_RVT U750 ( .A1(n1537), .A2(\inq_ary[15][85] ), .A3(n1741), .A4(
        \inq_ary[7][85] ), .Y(n664) );
  AO22X1_RVT U751 ( .A1(n1739), .A2(\inq_ary[2][85] ), .A3(n1749), .A4(
        \inq_ary[1][85] ), .Y(n663) );
  NOR4X1_RVT U752 ( .A1(n666), .A2(n665), .A3(n664), .A4(n663), .Y(n667) );
  NAND2X0_RVT U753 ( .A1(n668), .A2(n667), .Y(n669) );
  AO22X1_RVT U754 ( .A1(n1025), .A2(wrdata_d1[85]), .A3(n969), .A4(n669), .Y(
        n3410) );
  AO22X1_RVT U755 ( .A1(n1739), .A2(\inq_ary[2][47] ), .A3(n1537), .A4(
        \inq_ary[15][47] ), .Y(n673) );
  AO22X1_RVT U756 ( .A1(n1740), .A2(\inq_ary[12][47] ), .A3(n1741), .A4(
        \inq_ary[7][47] ), .Y(n672) );
  AO22X1_RVT U757 ( .A1(n1747), .A2(\inq_ary[5][47] ), .A3(n1748), .A4(
        \inq_ary[10][47] ), .Y(n671) );
  AO22X1_RVT U758 ( .A1(n1750), .A2(\inq_ary[11][47] ), .A3(n1751), .A4(
        \inq_ary[9][47] ), .Y(n670) );
  NOR4X1_RVT U759 ( .A1(n673), .A2(n672), .A3(n671), .A4(n670), .Y(n679) );
  AO22X1_RVT U760 ( .A1(n1729), .A2(\inq_ary[4][47] ), .A3(n1612), .A4(
        \inq_ary[8][47] ), .Y(n677) );
  AO22X1_RVT U761 ( .A1(n1686), .A2(\inq_ary[0][47] ), .A3(n1749), .A4(
        \inq_ary[1][47] ), .Y(n676) );
  AO22X1_RVT U762 ( .A1(n1742), .A2(\inq_ary[3][47] ), .A3(n1711), .A4(
        \inq_ary[13][47] ), .Y(n675) );
  AO22X1_RVT U763 ( .A1(n1554), .A2(\inq_ary[14][47] ), .A3(n1738), .A4(
        \inq_ary[6][47] ), .Y(n674) );
  NOR4X1_RVT U764 ( .A1(n677), .A2(n676), .A3(n675), .A4(n674), .Y(n678) );
  NAND2X0_RVT U765 ( .A1(n679), .A2(n678), .Y(n680) );
  AO22X1_RVT U766 ( .A1(n1598), .A2(wrdata_d1[47]), .A3(n2), .A4(n680), .Y(
        n3381) );
  AO22X1_RVT U767 ( .A1(n1749), .A2(\inq_ary[1][86] ), .A3(n1751), .A4(
        \inq_ary[9][86] ), .Y(n684) );
  AO22X1_RVT U768 ( .A1(n1750), .A2(\inq_ary[11][86] ), .A3(n1738), .A4(
        \inq_ary[6][86] ), .Y(n683) );
  AO22X1_RVT U769 ( .A1(n1739), .A2(\inq_ary[2][86] ), .A3(n1748), .A4(
        \inq_ary[10][86] ), .Y(n682) );
  AO22X1_RVT U770 ( .A1(n1747), .A2(\inq_ary[5][86] ), .A3(n1711), .A4(
        \inq_ary[13][86] ), .Y(n681) );
  NOR4X1_RVT U771 ( .A1(n684), .A2(n683), .A3(n682), .A4(n681), .Y(n690) );
  AO22X1_RVT U772 ( .A1(n1612), .A2(\inq_ary[8][86] ), .A3(n1741), .A4(
        \inq_ary[7][86] ), .Y(n688) );
  AO22X1_RVT U773 ( .A1(n1554), .A2(\inq_ary[14][86] ), .A3(n1742), .A4(
        \inq_ary[3][86] ), .Y(n687) );
  AO22X1_RVT U774 ( .A1(n1537), .A2(\inq_ary[15][86] ), .A3(n1740), .A4(
        \inq_ary[12][86] ), .Y(n686) );
  AO22X1_RVT U775 ( .A1(n1729), .A2(\inq_ary[4][86] ), .A3(n1686), .A4(
        \inq_ary[0][86] ), .Y(n685) );
  NOR4X1_RVT U776 ( .A1(n688), .A2(n687), .A3(n686), .A4(n685), .Y(n689) );
  NAND2X0_RVT U777 ( .A1(n690), .A2(n689), .Y(n691) );
  AO22X1_RVT U778 ( .A1(n1684), .A2(wrdata_d1[86]), .A3(n969), .A4(n691), .Y(
        n3412) );
  AO22X1_RVT U779 ( .A1(n1740), .A2(\inq_ary[12][87] ), .A3(n1747), .A4(
        \inq_ary[5][87] ), .Y(n695) );
  AO22X1_RVT U780 ( .A1(n1686), .A2(\inq_ary[0][87] ), .A3(n1749), .A4(
        \inq_ary[1][87] ), .Y(n694) );
  AO22X1_RVT U781 ( .A1(n1739), .A2(\inq_ary[2][87] ), .A3(n1750), .A4(
        \inq_ary[11][87] ), .Y(n693) );
  AO22X1_RVT U782 ( .A1(n1742), .A2(\inq_ary[3][87] ), .A3(n1748), .A4(
        \inq_ary[10][87] ), .Y(n692) );
  NOR4X1_RVT U783 ( .A1(n695), .A2(n694), .A3(n693), .A4(n692), .Y(n701) );
  AO22X1_RVT U784 ( .A1(n1729), .A2(\inq_ary[4][87] ), .A3(n1741), .A4(
        \inq_ary[7][87] ), .Y(n699) );
  AO22X1_RVT U785 ( .A1(n1554), .A2(\inq_ary[14][87] ), .A3(n1751), .A4(
        \inq_ary[9][87] ), .Y(n698) );
  AO22X1_RVT U786 ( .A1(n1612), .A2(\inq_ary[8][87] ), .A3(n1738), .A4(
        \inq_ary[6][87] ), .Y(n697) );
  AO22X1_RVT U787 ( .A1(n1537), .A2(\inq_ary[15][87] ), .A3(n1711), .A4(
        \inq_ary[13][87] ), .Y(n696) );
  NOR4X1_RVT U788 ( .A1(n699), .A2(n698), .A3(n697), .A4(n696), .Y(n700) );
  NAND2X0_RVT U789 ( .A1(n701), .A2(n700), .Y(n702) );
  AO22X1_RVT U790 ( .A1(n1477), .A2(wrdata_d1[87]), .A3(n1759), .A4(n702), .Y(
        n3414) );
  AO22X1_RVT U791 ( .A1(n1748), .A2(\inq_ary[10][46] ), .A3(n1751), .A4(
        \inq_ary[9][46] ), .Y(n706) );
  AO22X1_RVT U792 ( .A1(n1554), .A2(\inq_ary[14][46] ), .A3(n1729), .A4(
        \inq_ary[4][46] ), .Y(n705) );
  AO22X1_RVT U793 ( .A1(n1686), .A2(\inq_ary[0][46] ), .A3(n1747), .A4(
        \inq_ary[5][46] ), .Y(n704) );
  AO22X1_RVT U794 ( .A1(n1742), .A2(\inq_ary[3][46] ), .A3(n1537), .A4(
        \inq_ary[15][46] ), .Y(n703) );
  NOR4X1_RVT U795 ( .A1(n706), .A2(n705), .A3(n704), .A4(n703), .Y(n712) );
  AO22X1_RVT U796 ( .A1(n1612), .A2(\inq_ary[8][46] ), .A3(n1741), .A4(
        \inq_ary[7][46] ), .Y(n710) );
  AO22X1_RVT U797 ( .A1(n1749), .A2(\inq_ary[1][46] ), .A3(n1711), .A4(
        \inq_ary[13][46] ), .Y(n709) );
  AO22X1_RVT U798 ( .A1(n1740), .A2(\inq_ary[12][46] ), .A3(n1738), .A4(
        \inq_ary[6][46] ), .Y(n708) );
  AO22X1_RVT U799 ( .A1(n1739), .A2(\inq_ary[2][46] ), .A3(n1750), .A4(
        \inq_ary[11][46] ), .Y(n707) );
  NOR4X1_RVT U800 ( .A1(n710), .A2(n709), .A3(n708), .A4(n707), .Y(n711) );
  NAND2X0_RVT U801 ( .A1(n712), .A2(n711), .Y(n713) );
  AO22X1_RVT U802 ( .A1(n1598), .A2(wrdata_d1[46]), .A3(n946), .A4(n713), .Y(
        n3379) );
  AO22X1_RVT U803 ( .A1(n1739), .A2(\inq_ary[2][45] ), .A3(n1741), .A4(
        \inq_ary[7][45] ), .Y(n717) );
  AO22X1_RVT U804 ( .A1(n1554), .A2(\inq_ary[14][45] ), .A3(n1751), .A4(
        \inq_ary[9][45] ), .Y(n716) );
  AO22X1_RVT U805 ( .A1(n1749), .A2(\inq_ary[1][45] ), .A3(n1711), .A4(
        \inq_ary[13][45] ), .Y(n715) );
  AO22X1_RVT U806 ( .A1(n1742), .A2(\inq_ary[3][45] ), .A3(n1537), .A4(
        \inq_ary[15][45] ), .Y(n714) );
  NOR4X1_RVT U807 ( .A1(n717), .A2(n716), .A3(n715), .A4(n714), .Y(n723) );
  AO22X1_RVT U808 ( .A1(n1612), .A2(\inq_ary[8][45] ), .A3(n1738), .A4(
        \inq_ary[6][45] ), .Y(n721) );
  AO22X1_RVT U809 ( .A1(n1729), .A2(\inq_ary[4][45] ), .A3(n1740), .A4(
        \inq_ary[12][45] ), .Y(n720) );
  AO22X1_RVT U810 ( .A1(n1747), .A2(\inq_ary[5][45] ), .A3(n1748), .A4(
        \inq_ary[10][45] ), .Y(n719) );
  AO22X1_RVT U811 ( .A1(n1686), .A2(\inq_ary[0][45] ), .A3(n1750), .A4(
        \inq_ary[11][45] ), .Y(n718) );
  NOR4X1_RVT U812 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .Y(n722) );
  NAND2X0_RVT U813 ( .A1(n723), .A2(n722), .Y(n724) );
  AO22X1_RVT U814 ( .A1(n1025), .A2(wrdata_d1[45]), .A3(n2), .A4(n724), .Y(
        n3377) );
  AO22X1_RVT U815 ( .A1(n1729), .A2(\inq_ary[4][74] ), .A3(n1750), .A4(
        \inq_ary[11][74] ), .Y(n728) );
  AO22X1_RVT U816 ( .A1(n1554), .A2(\inq_ary[14][74] ), .A3(n1741), .A4(
        \inq_ary[7][74] ), .Y(n727) );
  AO22X1_RVT U817 ( .A1(n1742), .A2(\inq_ary[3][74] ), .A3(n1751), .A4(
        \inq_ary[9][74] ), .Y(n726) );
  AO22X1_RVT U818 ( .A1(n1739), .A2(\inq_ary[2][74] ), .A3(n1740), .A4(
        \inq_ary[12][74] ), .Y(n725) );
  NOR4X1_RVT U819 ( .A1(n728), .A2(n727), .A3(n726), .A4(n725), .Y(n734) );
  AO22X1_RVT U820 ( .A1(n1686), .A2(\inq_ary[0][74] ), .A3(n1738), .A4(
        \inq_ary[6][74] ), .Y(n732) );
  AO22X1_RVT U821 ( .A1(n1537), .A2(\inq_ary[15][74] ), .A3(n1612), .A4(
        \inq_ary[8][74] ), .Y(n731) );
  AO22X1_RVT U822 ( .A1(n1711), .A2(\inq_ary[13][74] ), .A3(n1748), .A4(
        \inq_ary[10][74] ), .Y(n730) );
  AO22X1_RVT U823 ( .A1(n1749), .A2(\inq_ary[1][74] ), .A3(n1747), .A4(
        \inq_ary[5][74] ), .Y(n729) );
  NOR4X1_RVT U824 ( .A1(n732), .A2(n731), .A3(n730), .A4(n729), .Y(n733) );
  NAND2X0_RVT U825 ( .A1(n734), .A2(n733), .Y(n735) );
  AO22X1_RVT U826 ( .A1(n3), .A2(wrdata_d1[74]), .A3(n969), .A4(n735), .Y(
        n3405) );
  AO22X1_RVT U827 ( .A1(n1748), .A2(\inq_ary[10][75] ), .A3(n1751), .A4(
        \inq_ary[9][75] ), .Y(n739) );
  AO22X1_RVT U828 ( .A1(n1686), .A2(\inq_ary[0][75] ), .A3(n1738), .A4(
        \inq_ary[6][75] ), .Y(n738) );
  AO22X1_RVT U829 ( .A1(n1739), .A2(\inq_ary[2][75] ), .A3(n1747), .A4(
        \inq_ary[5][75] ), .Y(n737) );
  AO22X1_RVT U830 ( .A1(n1742), .A2(\inq_ary[3][75] ), .A3(n1711), .A4(
        \inq_ary[13][75] ), .Y(n736) );
  NOR4X1_RVT U831 ( .A1(n739), .A2(n738), .A3(n737), .A4(n736), .Y(n745) );
  AO22X1_RVT U832 ( .A1(n1554), .A2(\inq_ary[14][75] ), .A3(n1749), .A4(
        \inq_ary[1][75] ), .Y(n743) );
  AO22X1_RVT U833 ( .A1(n1729), .A2(\inq_ary[4][75] ), .A3(n1537), .A4(
        \inq_ary[15][75] ), .Y(n742) );
  AO22X1_RVT U834 ( .A1(n1612), .A2(\inq_ary[8][75] ), .A3(n1740), .A4(
        \inq_ary[12][75] ), .Y(n741) );
  AO22X1_RVT U835 ( .A1(n1741), .A2(\inq_ary[7][75] ), .A3(n1750), .A4(
        \inq_ary[11][75] ), .Y(n740) );
  NOR4X1_RVT U836 ( .A1(n743), .A2(n742), .A3(n741), .A4(n740), .Y(n744) );
  NAND2X0_RVT U837 ( .A1(n745), .A2(n744), .Y(n746) );
  AO22X1_RVT U838 ( .A1(n3), .A2(wrdata_d1[75]), .A3(n2), .A4(n746), .Y(n3407)
         );
  AO22X1_RVT U839 ( .A1(n1742), .A2(\inq_ary[3][76] ), .A3(n1750), .A4(
        \inq_ary[11][76] ), .Y(n750) );
  AO22X1_RVT U840 ( .A1(n1741), .A2(\inq_ary[7][76] ), .A3(n1748), .A4(
        \inq_ary[10][76] ), .Y(n749) );
  AO22X1_RVT U841 ( .A1(n1612), .A2(\inq_ary[8][76] ), .A3(n1740), .A4(
        \inq_ary[12][76] ), .Y(n748) );
  AO22X1_RVT U842 ( .A1(n1729), .A2(\inq_ary[4][76] ), .A3(n1751), .A4(
        \inq_ary[9][76] ), .Y(n747) );
  NOR4X1_RVT U843 ( .A1(n750), .A2(n749), .A3(n748), .A4(n747), .Y(n756) );
  AO22X1_RVT U844 ( .A1(n1686), .A2(\inq_ary[0][76] ), .A3(n1749), .A4(
        \inq_ary[1][76] ), .Y(n754) );
  AO22X1_RVT U845 ( .A1(n1738), .A2(\inq_ary[6][76] ), .A3(n1711), .A4(
        \inq_ary[13][76] ), .Y(n753) );
  AO22X1_RVT U846 ( .A1(n1739), .A2(\inq_ary[2][76] ), .A3(n1554), .A4(
        \inq_ary[14][76] ), .Y(n752) );
  AO22X1_RVT U847 ( .A1(n1537), .A2(\inq_ary[15][76] ), .A3(n1747), .A4(
        \inq_ary[5][76] ), .Y(n751) );
  NOR4X1_RVT U848 ( .A1(n754), .A2(n753), .A3(n752), .A4(n751), .Y(n755) );
  NAND2X0_RVT U849 ( .A1(n756), .A2(n755), .Y(n757) );
  AO22X1_RVT U850 ( .A1(n758), .A2(wrdata_d1[76]), .A3(n1), .A4(n757), .Y(
        n3400) );
  AO22X1_RVT U851 ( .A1(n1750), .A2(\inq_ary[11][77] ), .A3(n1738), .A4(
        \inq_ary[6][77] ), .Y(n762) );
  AO22X1_RVT U852 ( .A1(n1741), .A2(\inq_ary[7][77] ), .A3(n1711), .A4(
        \inq_ary[13][77] ), .Y(n761) );
  AO22X1_RVT U853 ( .A1(n1739), .A2(\inq_ary[2][77] ), .A3(n1554), .A4(
        \inq_ary[14][77] ), .Y(n760) );
  AO22X1_RVT U854 ( .A1(n1729), .A2(\inq_ary[4][77] ), .A3(n1686), .A4(
        \inq_ary[0][77] ), .Y(n759) );
  NOR4X1_RVT U855 ( .A1(n762), .A2(n761), .A3(n760), .A4(n759), .Y(n768) );
  AO22X1_RVT U856 ( .A1(n1742), .A2(\inq_ary[3][77] ), .A3(n1747), .A4(
        \inq_ary[5][77] ), .Y(n766) );
  AO22X1_RVT U857 ( .A1(n1612), .A2(\inq_ary[8][77] ), .A3(n1740), .A4(
        \inq_ary[12][77] ), .Y(n765) );
  AO22X1_RVT U858 ( .A1(n1748), .A2(\inq_ary[10][77] ), .A3(n1751), .A4(
        \inq_ary[9][77] ), .Y(n764) );
  AO22X1_RVT U859 ( .A1(n1537), .A2(\inq_ary[15][77] ), .A3(n1749), .A4(
        \inq_ary[1][77] ), .Y(n763) );
  NOR4X1_RVT U860 ( .A1(n766), .A2(n765), .A3(n764), .A4(n763), .Y(n767) );
  NAND2X0_RVT U861 ( .A1(n768), .A2(n767), .Y(n769) );
  AO22X1_RVT U862 ( .A1(n3), .A2(wrdata_d1[77]), .A3(n1), .A4(n769), .Y(n3402)
         );
  AO22X1_RVT U863 ( .A1(n1748), .A2(\inq_ary[10][51] ), .A3(n1751), .A4(
        \inq_ary[9][51] ), .Y(n773) );
  AO22X1_RVT U864 ( .A1(n1612), .A2(\inq_ary[8][51] ), .A3(n1750), .A4(
        \inq_ary[11][51] ), .Y(n772) );
  AO22X1_RVT U865 ( .A1(n1686), .A2(\inq_ary[0][51] ), .A3(n1738), .A4(
        \inq_ary[6][51] ), .Y(n771) );
  AO22X1_RVT U866 ( .A1(n1554), .A2(\inq_ary[14][51] ), .A3(n1742), .A4(
        \inq_ary[3][51] ), .Y(n770) );
  NOR4X1_RVT U867 ( .A1(n773), .A2(n772), .A3(n771), .A4(n770), .Y(n779) );
  AO22X1_RVT U868 ( .A1(n1741), .A2(\inq_ary[7][51] ), .A3(n1747), .A4(
        \inq_ary[5][51] ), .Y(n777) );
  AO22X1_RVT U869 ( .A1(n1537), .A2(\inq_ary[15][51] ), .A3(n1740), .A4(
        \inq_ary[12][51] ), .Y(n776) );
  AO22X1_RVT U870 ( .A1(n1729), .A2(\inq_ary[4][51] ), .A3(n1711), .A4(
        \inq_ary[13][51] ), .Y(n775) );
  AO22X1_RVT U871 ( .A1(n1739), .A2(\inq_ary[2][51] ), .A3(n1749), .A4(
        \inq_ary[1][51] ), .Y(n774) );
  NOR4X1_RVT U872 ( .A1(n777), .A2(n776), .A3(n775), .A4(n774), .Y(n778) );
  NAND2X0_RVT U873 ( .A1(n779), .A2(n778), .Y(n780) );
  AO22X1_RVT U874 ( .A1(n1025), .A2(wrdata_d1[51]), .A3(n1), .A4(n780), .Y(
        n3389) );
  AO22X1_RVT U875 ( .A1(n1738), .A2(\inq_ary[6][78] ), .A3(n1751), .A4(
        \inq_ary[9][78] ), .Y(n784) );
  AO22X1_RVT U876 ( .A1(n1612), .A2(\inq_ary[8][78] ), .A3(n1750), .A4(
        \inq_ary[11][78] ), .Y(n783) );
  AO22X1_RVT U877 ( .A1(n1739), .A2(\inq_ary[2][78] ), .A3(n1686), .A4(
        \inq_ary[0][78] ), .Y(n782) );
  AO22X1_RVT U878 ( .A1(n1554), .A2(\inq_ary[14][78] ), .A3(n1711), .A4(
        \inq_ary[13][78] ), .Y(n781) );
  NOR4X1_RVT U879 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .Y(n790) );
  AO22X1_RVT U880 ( .A1(n1729), .A2(\inq_ary[4][78] ), .A3(n1537), .A4(
        \inq_ary[15][78] ), .Y(n788) );
  AO22X1_RVT U881 ( .A1(n1747), .A2(\inq_ary[5][78] ), .A3(n1748), .A4(
        \inq_ary[10][78] ), .Y(n787) );
  AO22X1_RVT U882 ( .A1(n1742), .A2(\inq_ary[3][78] ), .A3(n1741), .A4(
        \inq_ary[7][78] ), .Y(n786) );
  AO22X1_RVT U883 ( .A1(n1740), .A2(\inq_ary[12][78] ), .A3(n1749), .A4(
        \inq_ary[1][78] ), .Y(n785) );
  NOR4X1_RVT U884 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .Y(n789) );
  NAND2X0_RVT U885 ( .A1(n790), .A2(n789), .Y(n791) );
  AO22X1_RVT U886 ( .A1(n3), .A2(wrdata_d1[78]), .A3(n1759), .A4(n791), .Y(
        n3404) );
  AO22X1_RVT U887 ( .A1(n1739), .A2(\inq_ary[2][79] ), .A3(n1711), .A4(
        \inq_ary[13][79] ), .Y(n795) );
  AO22X1_RVT U888 ( .A1(n1686), .A2(\inq_ary[0][79] ), .A3(n1537), .A4(
        \inq_ary[15][79] ), .Y(n794) );
  AO22X1_RVT U889 ( .A1(n1554), .A2(\inq_ary[14][79] ), .A3(n1747), .A4(
        \inq_ary[5][79] ), .Y(n793) );
  AO22X1_RVT U890 ( .A1(n1740), .A2(\inq_ary[12][79] ), .A3(n1741), .A4(
        \inq_ary[7][79] ), .Y(n792) );
  NOR4X1_RVT U891 ( .A1(n795), .A2(n794), .A3(n793), .A4(n792), .Y(n801) );
  AO22X1_RVT U892 ( .A1(n1742), .A2(\inq_ary[3][79] ), .A3(n1750), .A4(
        \inq_ary[11][79] ), .Y(n799) );
  AO22X1_RVT U893 ( .A1(n1729), .A2(\inq_ary[4][79] ), .A3(n1738), .A4(
        \inq_ary[6][79] ), .Y(n798) );
  AO22X1_RVT U894 ( .A1(n1749), .A2(\inq_ary[1][79] ), .A3(n1748), .A4(
        \inq_ary[10][79] ), .Y(n797) );
  AO22X1_RVT U895 ( .A1(n1612), .A2(\inq_ary[8][79] ), .A3(n1751), .A4(
        \inq_ary[9][79] ), .Y(n796) );
  NOR4X1_RVT U896 ( .A1(n799), .A2(n798), .A3(n797), .A4(n796), .Y(n800) );
  NAND2X0_RVT U897 ( .A1(n801), .A2(n800), .Y(n802) );
  AO22X1_RVT U898 ( .A1(n3), .A2(wrdata_d1[79]), .A3(n1489), .A4(n802), .Y(
        n3406) );
  AO22X1_RVT U899 ( .A1(n1612), .A2(\inq_ary[8][50] ), .A3(n1747), .A4(
        \inq_ary[5][50] ), .Y(n806) );
  AO22X1_RVT U900 ( .A1(n1554), .A2(\inq_ary[14][50] ), .A3(n1748), .A4(
        \inq_ary[10][50] ), .Y(n805) );
  AO22X1_RVT U901 ( .A1(n1686), .A2(\inq_ary[0][50] ), .A3(n1537), .A4(
        \inq_ary[15][50] ), .Y(n804) );
  AO22X1_RVT U902 ( .A1(n1741), .A2(\inq_ary[7][50] ), .A3(n1738), .A4(
        \inq_ary[6][50] ), .Y(n803) );
  NOR4X1_RVT U903 ( .A1(n806), .A2(n805), .A3(n804), .A4(n803), .Y(n812) );
  AO22X1_RVT U904 ( .A1(n1740), .A2(\inq_ary[12][50] ), .A3(n1711), .A4(
        \inq_ary[13][50] ), .Y(n810) );
  AO22X1_RVT U905 ( .A1(n1729), .A2(\inq_ary[4][50] ), .A3(n1749), .A4(
        \inq_ary[1][50] ), .Y(n809) );
  AO22X1_RVT U906 ( .A1(n1739), .A2(\inq_ary[2][50] ), .A3(n1751), .A4(
        \inq_ary[9][50] ), .Y(n808) );
  AO22X1_RVT U907 ( .A1(n1742), .A2(\inq_ary[3][50] ), .A3(n1750), .A4(
        \inq_ary[11][50] ), .Y(n807) );
  NOR4X1_RVT U908 ( .A1(n810), .A2(n809), .A3(n808), .A4(n807), .Y(n811) );
  NAND2X0_RVT U909 ( .A1(n812), .A2(n811), .Y(n813) );
  AO22X1_RVT U910 ( .A1(n1477), .A2(wrdata_d1[50]), .A3(n946), .A4(n813), .Y(
        n3387) );
  AO22X1_RVT U911 ( .A1(n1686), .A2(\inq_ary[0][80] ), .A3(n1612), .A4(
        \inq_ary[8][80] ), .Y(n817) );
  AO22X1_RVT U912 ( .A1(n1729), .A2(\inq_ary[4][80] ), .A3(n1748), .A4(
        \inq_ary[10][80] ), .Y(n816) );
  AO22X1_RVT U913 ( .A1(n1750), .A2(\inq_ary[11][80] ), .A3(n1751), .A4(
        \inq_ary[9][80] ), .Y(n815) );
  AO22X1_RVT U914 ( .A1(n1740), .A2(\inq_ary[12][80] ), .A3(n1711), .A4(
        \inq_ary[13][80] ), .Y(n814) );
  NOR4X1_RVT U915 ( .A1(n817), .A2(n816), .A3(n815), .A4(n814), .Y(n823) );
  AO22X1_RVT U916 ( .A1(n1742), .A2(\inq_ary[3][80] ), .A3(n1738), .A4(
        \inq_ary[6][80] ), .Y(n821) );
  AO22X1_RVT U917 ( .A1(n1749), .A2(\inq_ary[1][80] ), .A3(n1747), .A4(
        \inq_ary[5][80] ), .Y(n820) );
  AO22X1_RVT U918 ( .A1(n1739), .A2(\inq_ary[2][80] ), .A3(n1537), .A4(
        \inq_ary[15][80] ), .Y(n819) );
  AO22X1_RVT U919 ( .A1(n1554), .A2(\inq_ary[14][80] ), .A3(n1741), .A4(
        \inq_ary[7][80] ), .Y(n818) );
  NOR4X1_RVT U920 ( .A1(n821), .A2(n820), .A3(n819), .A4(n818), .Y(n822) );
  NAND2X0_RVT U921 ( .A1(n823), .A2(n822), .Y(n824) );
  AO22X1_RVT U922 ( .A1(n758), .A2(wrdata_d1[80]), .A3(n1), .A4(n824), .Y(
        n3409) );
  AO22X1_RVT U923 ( .A1(n1612), .A2(\inq_ary[8][81] ), .A3(n1741), .A4(
        \inq_ary[7][81] ), .Y(n828) );
  AO22X1_RVT U924 ( .A1(n1739), .A2(\inq_ary[2][81] ), .A3(n1751), .A4(
        \inq_ary[9][81] ), .Y(n827) );
  AO22X1_RVT U925 ( .A1(n1749), .A2(\inq_ary[1][81] ), .A3(n1750), .A4(
        \inq_ary[11][81] ), .Y(n826) );
  AO22X1_RVT U926 ( .A1(n1747), .A2(\inq_ary[5][81] ), .A3(n1738), .A4(
        \inq_ary[6][81] ), .Y(n825) );
  NOR4X1_RVT U927 ( .A1(n828), .A2(n827), .A3(n826), .A4(n825), .Y(n834) );
  AO22X1_RVT U928 ( .A1(n1742), .A2(\inq_ary[3][81] ), .A3(n1740), .A4(
        \inq_ary[12][81] ), .Y(n832) );
  AO22X1_RVT U929 ( .A1(n1554), .A2(\inq_ary[14][81] ), .A3(n1537), .A4(
        \inq_ary[15][81] ), .Y(n831) );
  AO22X1_RVT U930 ( .A1(n1686), .A2(\inq_ary[0][81] ), .A3(n1711), .A4(
        \inq_ary[13][81] ), .Y(n830) );
  AO22X1_RVT U931 ( .A1(n1729), .A2(\inq_ary[4][81] ), .A3(n1748), .A4(
        \inq_ary[10][81] ), .Y(n829) );
  NOR4X1_RVT U932 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .Y(n833) );
  NAND2X0_RVT U933 ( .A1(n834), .A2(n833), .Y(n835) );
  AO22X1_RVT U934 ( .A1(n1025), .A2(wrdata_d1[81]), .A3(n1), .A4(n835), .Y(
        n3411) );
  AO22X1_RVT U935 ( .A1(n1537), .A2(\inq_ary[15][49] ), .A3(n1750), .A4(
        \inq_ary[11][49] ), .Y(n839) );
  AO22X1_RVT U936 ( .A1(n1742), .A2(\inq_ary[3][49] ), .A3(n1740), .A4(
        \inq_ary[12][49] ), .Y(n838) );
  AO22X1_RVT U937 ( .A1(n1686), .A2(\inq_ary[0][49] ), .A3(n1741), .A4(
        \inq_ary[7][49] ), .Y(n837) );
  AO22X1_RVT U938 ( .A1(n1554), .A2(\inq_ary[14][49] ), .A3(n1612), .A4(
        \inq_ary[8][49] ), .Y(n836) );
  NOR4X1_RVT U939 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .Y(n845) );
  AO22X1_RVT U940 ( .A1(n1729), .A2(\inq_ary[4][49] ), .A3(n1747), .A4(
        \inq_ary[5][49] ), .Y(n843) );
  AO22X1_RVT U941 ( .A1(n1739), .A2(\inq_ary[2][49] ), .A3(n1711), .A4(
        \inq_ary[13][49] ), .Y(n842) );
  AO22X1_RVT U942 ( .A1(n1738), .A2(\inq_ary[6][49] ), .A3(n1748), .A4(
        \inq_ary[10][49] ), .Y(n841) );
  AO22X1_RVT U943 ( .A1(n1749), .A2(\inq_ary[1][49] ), .A3(n1751), .A4(
        \inq_ary[9][49] ), .Y(n840) );
  NOR4X1_RVT U944 ( .A1(n843), .A2(n842), .A3(n841), .A4(n840), .Y(n844) );
  NAND2X0_RVT U945 ( .A1(n845), .A2(n844), .Y(n846) );
  AO22X1_RVT U946 ( .A1(n3), .A2(wrdata_d1[49]), .A3(n946), .A4(n846), .Y(
        n3385) );
  AO22X1_RVT U947 ( .A1(n1742), .A2(\inq_ary[3][88] ), .A3(n1750), .A4(
        \inq_ary[11][88] ), .Y(n850) );
  AO22X1_RVT U948 ( .A1(n1554), .A2(\inq_ary[14][88] ), .A3(n1711), .A4(
        \inq_ary[13][88] ), .Y(n849) );
  AO22X1_RVT U949 ( .A1(n1747), .A2(\inq_ary[5][88] ), .A3(n1738), .A4(
        \inq_ary[6][88] ), .Y(n848) );
  AO22X1_RVT U950 ( .A1(n1537), .A2(\inq_ary[15][88] ), .A3(n1748), .A4(
        \inq_ary[10][88] ), .Y(n847) );
  NOR4X1_RVT U951 ( .A1(n850), .A2(n849), .A3(n848), .A4(n847), .Y(n856) );
  AO22X1_RVT U952 ( .A1(n1729), .A2(\inq_ary[4][88] ), .A3(n1740), .A4(
        \inq_ary[12][88] ), .Y(n854) );
  AO22X1_RVT U953 ( .A1(n1739), .A2(\inq_ary[2][88] ), .A3(n1749), .A4(
        \inq_ary[1][88] ), .Y(n853) );
  AO22X1_RVT U954 ( .A1(n1686), .A2(\inq_ary[0][88] ), .A3(n1612), .A4(
        \inq_ary[8][88] ), .Y(n852) );
  AO22X1_RVT U955 ( .A1(n1741), .A2(\inq_ary[7][88] ), .A3(n1751), .A4(
        \inq_ary[9][88] ), .Y(n851) );
  NOR4X1_RVT U956 ( .A1(n854), .A2(n853), .A3(n852), .A4(n851), .Y(n855) );
  NAND2X0_RVT U957 ( .A1(n856), .A2(n855), .Y(n857) );
  AO22X1_RVT U958 ( .A1(n3), .A2(wrdata_d1[88]), .A3(n969), .A4(n857), .Y(
        n3417) );
  AO22X1_RVT U959 ( .A1(n1729), .A2(\inq_ary[4][60] ), .A3(n1741), .A4(
        \inq_ary[7][60] ), .Y(n861) );
  AO22X1_RVT U960 ( .A1(n1740), .A2(\inq_ary[12][60] ), .A3(n1750), .A4(
        \inq_ary[11][60] ), .Y(n860) );
  AO22X1_RVT U961 ( .A1(n1739), .A2(\inq_ary[2][60] ), .A3(n1686), .A4(
        \inq_ary[0][60] ), .Y(n859) );
  AO22X1_RVT U962 ( .A1(n1554), .A2(\inq_ary[14][60] ), .A3(n1537), .A4(
        \inq_ary[15][60] ), .Y(n858) );
  NOR4X1_RVT U963 ( .A1(n861), .A2(n860), .A3(n859), .A4(n858), .Y(n867) );
  AO22X1_RVT U964 ( .A1(n1749), .A2(\inq_ary[1][60] ), .A3(n1751), .A4(
        \inq_ary[9][60] ), .Y(n865) );
  AO22X1_RVT U965 ( .A1(n1738), .A2(\inq_ary[6][60] ), .A3(n1711), .A4(
        \inq_ary[13][60] ), .Y(n864) );
  AO22X1_RVT U966 ( .A1(n1612), .A2(\inq_ary[8][60] ), .A3(n1747), .A4(
        \inq_ary[5][60] ), .Y(n863) );
  AO22X1_RVT U967 ( .A1(n1742), .A2(\inq_ary[3][60] ), .A3(n1748), .A4(
        \inq_ary[10][60] ), .Y(n862) );
  NOR4X1_RVT U968 ( .A1(n865), .A2(n864), .A3(n863), .A4(n862), .Y(n866) );
  NAND2X0_RVT U969 ( .A1(n867), .A2(n866), .Y(n868) );
  AO22X1_RVT U970 ( .A1(n1723), .A2(wrdata_d1[60]), .A3(n2), .A4(n868), .Y(
        n3390) );
  AO22X1_RVT U971 ( .A1(n1612), .A2(\inq_ary[8][141] ), .A3(n1747), .A4(
        \inq_ary[5][141] ), .Y(n872) );
  AO22X1_RVT U972 ( .A1(n1537), .A2(\inq_ary[15][141] ), .A3(n1748), .A4(
        \inq_ary[10][141] ), .Y(n871) );
  AO22X1_RVT U973 ( .A1(n1750), .A2(\inq_ary[11][141] ), .A3(n1751), .A4(
        \inq_ary[9][141] ), .Y(n870) );
  AO22X1_RVT U974 ( .A1(n1738), .A2(\inq_ary[6][141] ), .A3(n1711), .A4(
        \inq_ary[13][141] ), .Y(n869) );
  NOR4X1_RVT U975 ( .A1(n872), .A2(n871), .A3(n870), .A4(n869), .Y(n878) );
  AO22X1_RVT U976 ( .A1(n1739), .A2(\inq_ary[2][141] ), .A3(n1554), .A4(
        \inq_ary[14][141] ), .Y(n876) );
  AO22X1_RVT U977 ( .A1(n1686), .A2(\inq_ary[0][141] ), .A3(n1741), .A4(
        \inq_ary[7][141] ), .Y(n875) );
  AO22X1_RVT U978 ( .A1(n1742), .A2(\inq_ary[3][141] ), .A3(n1749), .A4(
        \inq_ary[1][141] ), .Y(n874) );
  AO22X1_RVT U979 ( .A1(n1729), .A2(\inq_ary[4][141] ), .A3(n1740), .A4(
        \inq_ary[12][141] ), .Y(n873) );
  NOR4X1_RVT U980 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .Y(n877) );
  NAND2X0_RVT U981 ( .A1(n878), .A2(n877), .Y(n879) );
  AO22X1_RVT U982 ( .A1(n1025), .A2(wrdata_d1[141]), .A3(n2), .A4(n879), .Y(
        n3466) );
  AO22X1_RVT U983 ( .A1(n1711), .A2(\inq_ary[13][142] ), .A3(n1748), .A4(
        \inq_ary[10][142] ), .Y(n883) );
  AO22X1_RVT U984 ( .A1(n1742), .A2(\inq_ary[3][142] ), .A3(n1740), .A4(
        \inq_ary[12][142] ), .Y(n882) );
  AO22X1_RVT U985 ( .A1(n1741), .A2(\inq_ary[7][142] ), .A3(n1747), .A4(
        \inq_ary[5][142] ), .Y(n881) );
  AO22X1_RVT U986 ( .A1(n1686), .A2(\inq_ary[0][142] ), .A3(n1738), .A4(
        \inq_ary[6][142] ), .Y(n880) );
  NOR4X1_RVT U987 ( .A1(n883), .A2(n882), .A3(n881), .A4(n880), .Y(n889) );
  AO22X1_RVT U988 ( .A1(n1749), .A2(\inq_ary[1][142] ), .A3(n1750), .A4(
        \inq_ary[11][142] ), .Y(n887) );
  AO22X1_RVT U989 ( .A1(n1554), .A2(\inq_ary[14][142] ), .A3(n1537), .A4(
        \inq_ary[15][142] ), .Y(n886) );
  AO22X1_RVT U990 ( .A1(n1729), .A2(\inq_ary[4][142] ), .A3(n1751), .A4(
        \inq_ary[9][142] ), .Y(n885) );
  AO22X1_RVT U991 ( .A1(n1739), .A2(\inq_ary[2][142] ), .A3(n1612), .A4(
        \inq_ary[8][142] ), .Y(n884) );
  NOR4X1_RVT U992 ( .A1(n887), .A2(n886), .A3(n885), .A4(n884), .Y(n888) );
  NAND2X0_RVT U993 ( .A1(n889), .A2(n888), .Y(n890) );
  AO22X1_RVT U994 ( .A1(n1025), .A2(wrdata_d1[142]), .A3(n2), .A4(n890), .Y(
        n3468) );
  AO22X1_RVT U995 ( .A1(n1742), .A2(\inq_ary[3][11] ), .A3(n1750), .A4(
        \inq_ary[11][11] ), .Y(n894) );
  AO22X1_RVT U996 ( .A1(n1612), .A2(\inq_ary[8][11] ), .A3(n1738), .A4(
        \inq_ary[6][11] ), .Y(n893) );
  AO22X1_RVT U997 ( .A1(n1537), .A2(\inq_ary[15][11] ), .A3(n1748), .A4(
        \inq_ary[10][11] ), .Y(n892) );
  AO22X1_RVT U998 ( .A1(n1740), .A2(\inq_ary[12][11] ), .A3(n1747), .A4(
        \inq_ary[5][11] ), .Y(n891) );
  NOR4X1_RVT U999 ( .A1(n894), .A2(n893), .A3(n892), .A4(n891), .Y(n900) );
  AO22X1_RVT U1000 ( .A1(n1711), .A2(\inq_ary[13][11] ), .A3(n1751), .A4(
        \inq_ary[9][11] ), .Y(n898) );
  AO22X1_RVT U1001 ( .A1(n1729), .A2(\inq_ary[4][11] ), .A3(n1741), .A4(
        \inq_ary[7][11] ), .Y(n897) );
  AO22X1_RVT U1002 ( .A1(n1686), .A2(\inq_ary[0][11] ), .A3(n1749), .A4(
        \inq_ary[1][11] ), .Y(n896) );
  AO22X1_RVT U1003 ( .A1(n1739), .A2(\inq_ary[2][11] ), .A3(n1554), .A4(
        \inq_ary[14][11] ), .Y(n895) );
  NOR4X1_RVT U1004 ( .A1(n898), .A2(n897), .A3(n896), .A4(n895), .Y(n899) );
  NAND2X0_RVT U1005 ( .A1(n900), .A2(n899), .Y(n901) );
  AO22X1_RVT U1006 ( .A1(n1760), .A2(wrdata_d1[11]), .A3(n969), .A4(n901), .Y(
        n3350) );
  AO22X1_RVT U1007 ( .A1(n1554), .A2(\inq_ary[14][143] ), .A3(n1751), .A4(
        \inq_ary[9][143] ), .Y(n905) );
  AO22X1_RVT U1008 ( .A1(n1739), .A2(\inq_ary[2][143] ), .A3(n1741), .A4(
        \inq_ary[7][143] ), .Y(n904) );
  AO22X1_RVT U1009 ( .A1(n1740), .A2(\inq_ary[12][143] ), .A3(n1747), .A4(
        \inq_ary[5][143] ), .Y(n903) );
  AO22X1_RVT U1010 ( .A1(n1749), .A2(\inq_ary[1][143] ), .A3(n1748), .A4(
        \inq_ary[10][143] ), .Y(n902) );
  NOR4X1_RVT U1011 ( .A1(n905), .A2(n904), .A3(n903), .A4(n902), .Y(n911) );
  AO22X1_RVT U1012 ( .A1(n1537), .A2(\inq_ary[15][143] ), .A3(n1738), .A4(
        \inq_ary[6][143] ), .Y(n909) );
  AO22X1_RVT U1013 ( .A1(n1729), .A2(\inq_ary[4][143] ), .A3(n1750), .A4(
        \inq_ary[11][143] ), .Y(n908) );
  AO22X1_RVT U1014 ( .A1(n1612), .A2(\inq_ary[8][143] ), .A3(n1711), .A4(
        \inq_ary[13][143] ), .Y(n907) );
  AO22X1_RVT U1015 ( .A1(n1742), .A2(\inq_ary[3][143] ), .A3(n1686), .A4(
        \inq_ary[0][143] ), .Y(n906) );
  NOR4X1_RVT U1016 ( .A1(n909), .A2(n908), .A3(n907), .A4(n906), .Y(n910) );
  NAND2X0_RVT U1017 ( .A1(n911), .A2(n910), .Y(n912) );
  AO22X1_RVT U1018 ( .A1(n1025), .A2(wrdata_d1[143]), .A3(n2), .A4(n912), .Y(
        n3470) );
  AO22X1_RVT U1019 ( .A1(n1729), .A2(\inq_ary[4][144] ), .A3(n1749), .A4(
        \inq_ary[1][144] ), .Y(n916) );
  AO22X1_RVT U1020 ( .A1(n1742), .A2(\inq_ary[3][144] ), .A3(n1751), .A4(
        \inq_ary[9][144] ), .Y(n915) );
  AO22X1_RVT U1021 ( .A1(n1612), .A2(\inq_ary[8][144] ), .A3(n1738), .A4(
        \inq_ary[6][144] ), .Y(n914) );
  AO22X1_RVT U1022 ( .A1(n1739), .A2(\inq_ary[2][144] ), .A3(n1711), .A4(
        \inq_ary[13][144] ), .Y(n913) );
  NOR4X1_RVT U1023 ( .A1(n916), .A2(n915), .A3(n914), .A4(n913), .Y(n922) );
  AO22X1_RVT U1024 ( .A1(n1686), .A2(\inq_ary[0][144] ), .A3(n1741), .A4(
        \inq_ary[7][144] ), .Y(n920) );
  AO22X1_RVT U1025 ( .A1(n1740), .A2(\inq_ary[12][144] ), .A3(n1747), .A4(
        \inq_ary[5][144] ), .Y(n919) );
  AO22X1_RVT U1026 ( .A1(n1537), .A2(\inq_ary[15][144] ), .A3(n1748), .A4(
        \inq_ary[10][144] ), .Y(n918) );
  AO22X1_RVT U1027 ( .A1(n1554), .A2(\inq_ary[14][144] ), .A3(n1750), .A4(
        \inq_ary[11][144] ), .Y(n917) );
  NOR4X1_RVT U1028 ( .A1(n920), .A2(n919), .A3(n918), .A4(n917), .Y(n921) );
  NAND2X0_RVT U1029 ( .A1(n922), .A2(n921), .Y(n923) );
  AO22X1_RVT U1030 ( .A1(n1684), .A2(wrdata_d1[144]), .A3(n2), .A4(n923), .Y(
        n3472) );
  AO22X1_RVT U1031 ( .A1(n1686), .A2(\inq_ary[0][24] ), .A3(n1751), .A4(
        \inq_ary[9][24] ), .Y(n927) );
  AO22X1_RVT U1032 ( .A1(n1740), .A2(\inq_ary[12][24] ), .A3(n1749), .A4(
        \inq_ary[1][24] ), .Y(n926) );
  AO22X1_RVT U1033 ( .A1(n1612), .A2(\inq_ary[8][24] ), .A3(n1741), .A4(
        \inq_ary[7][24] ), .Y(n925) );
  AO22X1_RVT U1034 ( .A1(n1747), .A2(\inq_ary[5][24] ), .A3(n1711), .A4(
        \inq_ary[13][24] ), .Y(n924) );
  NOR4X1_RVT U1035 ( .A1(n927), .A2(n926), .A3(n925), .A4(n924), .Y(n933) );
  AO22X1_RVT U1036 ( .A1(n1729), .A2(\inq_ary[4][24] ), .A3(n1537), .A4(
        \inq_ary[15][24] ), .Y(n931) );
  AO22X1_RVT U1037 ( .A1(n1554), .A2(\inq_ary[14][24] ), .A3(n1750), .A4(
        \inq_ary[11][24] ), .Y(n930) );
  AO22X1_RVT U1038 ( .A1(n1739), .A2(\inq_ary[2][24] ), .A3(n1742), .A4(
        \inq_ary[3][24] ), .Y(n929) );
  AO22X1_RVT U1039 ( .A1(n1738), .A2(\inq_ary[6][24] ), .A3(n1748), .A4(
        \inq_ary[10][24] ), .Y(n928) );
  NOR4X1_RVT U1040 ( .A1(n931), .A2(n930), .A3(n929), .A4(n928), .Y(n932) );
  NAND2X0_RVT U1041 ( .A1(n933), .A2(n932), .Y(n934) );
  AO22X1_RVT U1042 ( .A1(n1684), .A2(wrdata_d1[24]), .A3(n969), .A4(n934), .Y(
        n3360) );
  AO22X1_RVT U1043 ( .A1(n1740), .A2(\inq_ary[12][12] ), .A3(n1738), .A4(
        \inq_ary[6][12] ), .Y(n938) );
  AO22X1_RVT U1044 ( .A1(n1686), .A2(\inq_ary[0][12] ), .A3(n1612), .A4(
        \inq_ary[8][12] ), .Y(n937) );
  AO22X1_RVT U1045 ( .A1(n1554), .A2(\inq_ary[14][12] ), .A3(n1747), .A4(
        \inq_ary[5][12] ), .Y(n936) );
  AO22X1_RVT U1046 ( .A1(n1739), .A2(\inq_ary[2][12] ), .A3(n1729), .A4(
        \inq_ary[4][12] ), .Y(n935) );
  NOR4X1_RVT U1047 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .Y(n944) );
  AO22X1_RVT U1048 ( .A1(n1742), .A2(\inq_ary[3][12] ), .A3(n1750), .A4(
        \inq_ary[11][12] ), .Y(n942) );
  AO22X1_RVT U1049 ( .A1(n1748), .A2(\inq_ary[10][12] ), .A3(n1751), .A4(
        \inq_ary[9][12] ), .Y(n941) );
  AO22X1_RVT U1050 ( .A1(n1537), .A2(\inq_ary[15][12] ), .A3(n1749), .A4(
        \inq_ary[1][12] ), .Y(n940) );
  AO22X1_RVT U1051 ( .A1(n1741), .A2(\inq_ary[7][12] ), .A3(n1711), .A4(
        \inq_ary[13][12] ), .Y(n939) );
  NOR4X1_RVT U1052 ( .A1(n942), .A2(n941), .A3(n940), .A4(n939), .Y(n943) );
  NAND2X0_RVT U1053 ( .A1(n944), .A2(n943), .Y(n945) );
  AO22X1_RVT U1054 ( .A1(n1598), .A2(wrdata_d1[12]), .A3(n2), .A4(n945), .Y(
        n3343) );
  INVX1_RVT U1055 ( .A(n946), .Y(n1723) );
  AO22X1_RVT U1056 ( .A1(n1742), .A2(\inq_ary[3][145] ), .A3(n1612), .A4(
        \inq_ary[8][145] ), .Y(n950) );
  AO22X1_RVT U1057 ( .A1(n1729), .A2(\inq_ary[4][145] ), .A3(n1740), .A4(
        \inq_ary[12][145] ), .Y(n949) );
  AO22X1_RVT U1058 ( .A1(n1738), .A2(\inq_ary[6][145] ), .A3(n1711), .A4(
        \inq_ary[13][145] ), .Y(n948) );
  AO22X1_RVT U1059 ( .A1(n1747), .A2(\inq_ary[5][145] ), .A3(n1748), .A4(
        \inq_ary[10][145] ), .Y(n947) );
  NOR4X1_RVT U1060 ( .A1(n950), .A2(n949), .A3(n948), .A4(n947), .Y(n956) );
  AO22X1_RVT U1061 ( .A1(n1554), .A2(\inq_ary[14][145] ), .A3(n1751), .A4(
        \inq_ary[9][145] ), .Y(n954) );
  AO22X1_RVT U1062 ( .A1(n1739), .A2(\inq_ary[2][145] ), .A3(n1686), .A4(
        \inq_ary[0][145] ), .Y(n953) );
  AO22X1_RVT U1063 ( .A1(n1741), .A2(\inq_ary[7][145] ), .A3(n1750), .A4(
        \inq_ary[11][145] ), .Y(n952) );
  AO22X1_RVT U1064 ( .A1(n1537), .A2(\inq_ary[15][145] ), .A3(n1749), .A4(
        \inq_ary[1][145] ), .Y(n951) );
  NOR4X1_RVT U1065 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .Y(n955) );
  NAND2X0_RVT U1066 ( .A1(n956), .A2(n955), .Y(n957) );
  AO22X1_RVT U1067 ( .A1(n1723), .A2(wrdata_d1[145]), .A3(n2), .A4(n957), .Y(
        n3473) );
  INVX1_RVT U1068 ( .A(n1760), .Y(n1759) );
  AO22X1_RVT U1069 ( .A1(n1749), .A2(\inq_ary[1][146] ), .A3(n1747), .A4(
        \inq_ary[5][146] ), .Y(n961) );
  AO22X1_RVT U1070 ( .A1(n1739), .A2(\inq_ary[2][146] ), .A3(n1554), .A4(
        \inq_ary[14][146] ), .Y(n960) );
  AO22X1_RVT U1071 ( .A1(n1537), .A2(\inq_ary[15][146] ), .A3(n1748), .A4(
        \inq_ary[10][146] ), .Y(n959) );
  AO22X1_RVT U1072 ( .A1(n1740), .A2(\inq_ary[12][146] ), .A3(n1738), .A4(
        \inq_ary[6][146] ), .Y(n958) );
  NOR4X1_RVT U1073 ( .A1(n961), .A2(n960), .A3(n959), .A4(n958), .Y(n967) );
  AO22X1_RVT U1074 ( .A1(n1686), .A2(\inq_ary[0][146] ), .A3(n1612), .A4(
        \inq_ary[8][146] ), .Y(n965) );
  AO22X1_RVT U1075 ( .A1(n1729), .A2(\inq_ary[4][146] ), .A3(n1741), .A4(
        \inq_ary[7][146] ), .Y(n964) );
  AO22X1_RVT U1076 ( .A1(n1742), .A2(\inq_ary[3][146] ), .A3(n1751), .A4(
        \inq_ary[9][146] ), .Y(n963) );
  AO22X1_RVT U1077 ( .A1(n1750), .A2(\inq_ary[11][146] ), .A3(n1711), .A4(
        \inq_ary[13][146] ), .Y(n962) );
  NOR4X1_RVT U1078 ( .A1(n965), .A2(n964), .A3(n963), .A4(n962), .Y(n966) );
  NAND2X0_RVT U1079 ( .A1(n967), .A2(n966), .Y(n968) );
  AO22X1_RVT U1080 ( .A1(n1723), .A2(wrdata_d1[146]), .A3(n1759), .A4(n968), 
        .Y(n3474) );
  INVX1_RVT U1081 ( .A(n1598), .Y(n1489) );
  AO22X1_RVT U1082 ( .A1(n1740), .A2(\inq_ary[12][135] ), .A3(n1741), .A4(
        \inq_ary[7][135] ), .Y(n973) );
  AO22X1_RVT U1083 ( .A1(n1537), .A2(\inq_ary[15][135] ), .A3(n1748), .A4(
        \inq_ary[10][135] ), .Y(n972) );
  AO22X1_RVT U1084 ( .A1(n1747), .A2(\inq_ary[5][135] ), .A3(n1750), .A4(
        \inq_ary[11][135] ), .Y(n971) );
  AO22X1_RVT U1085 ( .A1(n1729), .A2(\inq_ary[4][135] ), .A3(n1751), .A4(
        \inq_ary[9][135] ), .Y(n970) );
  NOR4X1_RVT U1086 ( .A1(n973), .A2(n972), .A3(n971), .A4(n970), .Y(n979) );
  AO22X1_RVT U1087 ( .A1(n1742), .A2(\inq_ary[3][135] ), .A3(n1711), .A4(
        \inq_ary[13][135] ), .Y(n977) );
  AO22X1_RVT U1088 ( .A1(n1554), .A2(\inq_ary[14][135] ), .A3(n1686), .A4(
        \inq_ary[0][135] ), .Y(n976) );
  AO22X1_RVT U1089 ( .A1(n1612), .A2(\inq_ary[8][135] ), .A3(n1738), .A4(
        \inq_ary[6][135] ), .Y(n975) );
  AO22X1_RVT U1090 ( .A1(n1739), .A2(\inq_ary[2][135] ), .A3(n1749), .A4(
        \inq_ary[1][135] ), .Y(n974) );
  NOR4X1_RVT U1091 ( .A1(n977), .A2(n976), .A3(n975), .A4(n974), .Y(n978) );
  NAND2X0_RVT U1092 ( .A1(n979), .A2(n978), .Y(n980) );
  AO22X1_RVT U1093 ( .A1(n758), .A2(wrdata_d1[135]), .A3(n1489), .A4(n980), 
        .Y(n3462) );
  AO22X1_RVT U1094 ( .A1(n1742), .A2(\inq_ary[3][136] ), .A3(n1537), .A4(
        \inq_ary[15][136] ), .Y(n984) );
  AO22X1_RVT U1095 ( .A1(n1686), .A2(\inq_ary[0][136] ), .A3(n1612), .A4(
        \inq_ary[8][136] ), .Y(n983) );
  AO22X1_RVT U1096 ( .A1(n1554), .A2(\inq_ary[14][136] ), .A3(n1740), .A4(
        \inq_ary[12][136] ), .Y(n982) );
  AO22X1_RVT U1097 ( .A1(n1729), .A2(\inq_ary[4][136] ), .A3(n1749), .A4(
        \inq_ary[1][136] ), .Y(n981) );
  NOR4X1_RVT U1098 ( .A1(n984), .A2(n983), .A3(n982), .A4(n981), .Y(n990) );
  AO22X1_RVT U1099 ( .A1(n1738), .A2(\inq_ary[6][136] ), .A3(n1751), .A4(
        \inq_ary[9][136] ), .Y(n988) );
  AO22X1_RVT U1100 ( .A1(n1739), .A2(\inq_ary[2][136] ), .A3(n1750), .A4(
        \inq_ary[11][136] ), .Y(n987) );
  AO22X1_RVT U1101 ( .A1(n1741), .A2(\inq_ary[7][136] ), .A3(n1711), .A4(
        \inq_ary[13][136] ), .Y(n986) );
  AO22X1_RVT U1102 ( .A1(n1747), .A2(\inq_ary[5][136] ), .A3(n1748), .A4(
        \inq_ary[10][136] ), .Y(n985) );
  NOR4X1_RVT U1103 ( .A1(n988), .A2(n987), .A3(n986), .A4(n985), .Y(n989) );
  NAND2X0_RVT U1104 ( .A1(n990), .A2(n989), .Y(n991) );
  AO22X1_RVT U1105 ( .A1(n1025), .A2(wrdata_d1[136]), .A3(n2), .A4(n991), .Y(
        n3465) );
  AO22X1_RVT U1106 ( .A1(n1749), .A2(\inq_ary[1][8] ), .A3(n1741), .A4(
        \inq_ary[7][8] ), .Y(n995) );
  AO22X1_RVT U1107 ( .A1(n1740), .A2(\inq_ary[12][8] ), .A3(n1751), .A4(
        \inq_ary[9][8] ), .Y(n994) );
  AO22X1_RVT U1108 ( .A1(n1739), .A2(\inq_ary[2][8] ), .A3(n1686), .A4(
        \inq_ary[0][8] ), .Y(n993) );
  AO22X1_RVT U1109 ( .A1(n1742), .A2(\inq_ary[3][8] ), .A3(n1612), .A4(
        \inq_ary[8][8] ), .Y(n992) );
  NOR4X1_RVT U1110 ( .A1(n995), .A2(n994), .A3(n993), .A4(n992), .Y(n1001) );
  AO22X1_RVT U1111 ( .A1(n1729), .A2(\inq_ary[4][8] ), .A3(n1738), .A4(
        \inq_ary[6][8] ), .Y(n999) );
  AO22X1_RVT U1112 ( .A1(n1750), .A2(\inq_ary[11][8] ), .A3(n1711), .A4(
        \inq_ary[13][8] ), .Y(n998) );
  AO22X1_RVT U1113 ( .A1(n1554), .A2(\inq_ary[14][8] ), .A3(n1748), .A4(
        \inq_ary[10][8] ), .Y(n997) );
  AO22X1_RVT U1114 ( .A1(n1537), .A2(\inq_ary[15][8] ), .A3(n1747), .A4(
        \inq_ary[5][8] ), .Y(n996) );
  NOR4X1_RVT U1115 ( .A1(n999), .A2(n998), .A3(n997), .A4(n996), .Y(n1000) );
  NAND2X0_RVT U1116 ( .A1(n1001), .A2(n1000), .Y(n1002) );
  AO22X1_RVT U1117 ( .A1(n1760), .A2(wrdata_d1[8]), .A3(n2), .A4(n1002), .Y(
        n3344) );
  AO22X1_RVT U1118 ( .A1(n1537), .A2(\inq_ary[15][137] ), .A3(n1747), .A4(
        \inq_ary[5][137] ), .Y(n1006) );
  AO22X1_RVT U1119 ( .A1(n1729), .A2(\inq_ary[4][137] ), .A3(n1749), .A4(
        \inq_ary[1][137] ), .Y(n1005) );
  AO22X1_RVT U1120 ( .A1(n1742), .A2(\inq_ary[3][137] ), .A3(n1750), .A4(
        \inq_ary[11][137] ), .Y(n1004) );
  AO22X1_RVT U1121 ( .A1(n1740), .A2(\inq_ary[12][137] ), .A3(n1748), .A4(
        \inq_ary[10][137] ), .Y(n1003) );
  NOR4X1_RVT U1122 ( .A1(n1006), .A2(n1005), .A3(n1004), .A4(n1003), .Y(n1012)
         );
  AO22X1_RVT U1123 ( .A1(n1612), .A2(\inq_ary[8][137] ), .A3(n1738), .A4(
        \inq_ary[6][137] ), .Y(n1010) );
  AO22X1_RVT U1124 ( .A1(n1741), .A2(\inq_ary[7][137] ), .A3(n1711), .A4(
        \inq_ary[13][137] ), .Y(n1009) );
  AO22X1_RVT U1125 ( .A1(n1554), .A2(\inq_ary[14][137] ), .A3(n1686), .A4(
        \inq_ary[0][137] ), .Y(n1008) );
  AO22X1_RVT U1126 ( .A1(n1739), .A2(\inq_ary[2][137] ), .A3(n1751), .A4(
        \inq_ary[9][137] ), .Y(n1007) );
  NOR4X1_RVT U1127 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .Y(n1011)
         );
  NAND2X0_RVT U1128 ( .A1(n1012), .A2(n1011), .Y(n1013) );
  AO22X1_RVT U1129 ( .A1(n1025), .A2(wrdata_d1[137]), .A3(n2), .A4(n1013), .Y(
        n3467) );
  AO22X1_RVT U1130 ( .A1(n1739), .A2(\inq_ary[2][138] ), .A3(n1554), .A4(
        \inq_ary[14][138] ), .Y(n1017) );
  AO22X1_RVT U1131 ( .A1(n1612), .A2(\inq_ary[8][138] ), .A3(n1749), .A4(
        \inq_ary[1][138] ), .Y(n1016) );
  AO22X1_RVT U1132 ( .A1(n1740), .A2(\inq_ary[12][138] ), .A3(n1741), .A4(
        \inq_ary[7][138] ), .Y(n1015) );
  AO22X1_RVT U1133 ( .A1(n1711), .A2(\inq_ary[13][138] ), .A3(n1748), .A4(
        \inq_ary[10][138] ), .Y(n1014) );
  NOR4X1_RVT U1134 ( .A1(n1017), .A2(n1016), .A3(n1015), .A4(n1014), .Y(n1023)
         );
  AO22X1_RVT U1135 ( .A1(n1686), .A2(\inq_ary[0][138] ), .A3(n1537), .A4(
        \inq_ary[15][138] ), .Y(n1021) );
  AO22X1_RVT U1136 ( .A1(n1742), .A2(\inq_ary[3][138] ), .A3(n1747), .A4(
        \inq_ary[5][138] ), .Y(n1020) );
  AO22X1_RVT U1137 ( .A1(n1750), .A2(\inq_ary[11][138] ), .A3(n1738), .A4(
        \inq_ary[6][138] ), .Y(n1019) );
  AO22X1_RVT U1138 ( .A1(n1729), .A2(\inq_ary[4][138] ), .A3(n1751), .A4(
        \inq_ary[9][138] ), .Y(n1018) );
  NOR4X1_RVT U1139 ( .A1(n1021), .A2(n1020), .A3(n1019), .A4(n1018), .Y(n1022)
         );
  NAND2X0_RVT U1140 ( .A1(n1023), .A2(n1022), .Y(n1024) );
  AO22X1_RVT U1141 ( .A1(n1025), .A2(wrdata_d1[138]), .A3(n2), .A4(n1024), .Y(
        n3469) );
  AO22X1_RVT U1142 ( .A1(n1750), .A2(\inq_ary[11][9] ), .A3(n1751), .A4(
        \inq_ary[9][9] ), .Y(n1029) );
  AO22X1_RVT U1143 ( .A1(n1612), .A2(\inq_ary[8][9] ), .A3(n1738), .A4(
        \inq_ary[6][9] ), .Y(n1028) );
  AO22X1_RVT U1144 ( .A1(n1686), .A2(\inq_ary[0][9] ), .A3(n1747), .A4(
        \inq_ary[5][9] ), .Y(n1027) );
  AO22X1_RVT U1145 ( .A1(n1740), .A2(\inq_ary[12][9] ), .A3(n1749), .A4(
        \inq_ary[1][9] ), .Y(n1026) );
  NOR4X1_RVT U1146 ( .A1(n1029), .A2(n1028), .A3(n1027), .A4(n1026), .Y(n1035)
         );
  AO22X1_RVT U1147 ( .A1(n1739), .A2(\inq_ary[2][9] ), .A3(n1741), .A4(
        \inq_ary[7][9] ), .Y(n1033) );
  AO22X1_RVT U1148 ( .A1(n1742), .A2(\inq_ary[3][9] ), .A3(n1711), .A4(
        \inq_ary[13][9] ), .Y(n1032) );
  AO22X1_RVT U1149 ( .A1(n1729), .A2(\inq_ary[4][9] ), .A3(n1748), .A4(
        \inq_ary[10][9] ), .Y(n1031) );
  AO22X1_RVT U1150 ( .A1(n1554), .A2(\inq_ary[14][9] ), .A3(n1537), .A4(
        \inq_ary[15][9] ), .Y(n1030) );
  NOR4X1_RVT U1151 ( .A1(n1033), .A2(n1032), .A3(n1031), .A4(n1030), .Y(n1034)
         );
  NAND2X0_RVT U1152 ( .A1(n1035), .A2(n1034), .Y(n1036) );
  AO22X1_RVT U1153 ( .A1(n1477), .A2(wrdata_d1[9]), .A3(n2), .A4(n1036), .Y(
        n3346) );
  AO22X1_RVT U1154 ( .A1(n1739), .A2(\inq_ary[2][139] ), .A3(n1740), .A4(
        \inq_ary[12][139] ), .Y(n1040) );
  AO22X1_RVT U1155 ( .A1(n1537), .A2(\inq_ary[15][139] ), .A3(n1749), .A4(
        \inq_ary[1][139] ), .Y(n1039) );
  AO22X1_RVT U1156 ( .A1(n1612), .A2(\inq_ary[8][139] ), .A3(n1748), .A4(
        \inq_ary[10][139] ), .Y(n1038) );
  AO22X1_RVT U1157 ( .A1(n1554), .A2(\inq_ary[14][139] ), .A3(n1738), .A4(
        \inq_ary[6][139] ), .Y(n1037) );
  NOR4X1_RVT U1158 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), .Y(n1046)
         );
  AO22X1_RVT U1159 ( .A1(n1686), .A2(\inq_ary[0][139] ), .A3(n1741), .A4(
        \inq_ary[7][139] ), .Y(n1044) );
  AO22X1_RVT U1160 ( .A1(n1747), .A2(\inq_ary[5][139] ), .A3(n1750), .A4(
        \inq_ary[11][139] ), .Y(n1043) );
  AO22X1_RVT U1161 ( .A1(n1742), .A2(\inq_ary[3][139] ), .A3(n1711), .A4(
        \inq_ary[13][139] ), .Y(n1042) );
  AO22X1_RVT U1162 ( .A1(n1729), .A2(\inq_ary[4][139] ), .A3(n1751), .A4(
        \inq_ary[9][139] ), .Y(n1041) );
  NOR4X1_RVT U1163 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), .Y(n1045)
         );
  NAND2X0_RVT U1164 ( .A1(n1046), .A2(n1045), .Y(n1047) );
  AO22X1_RVT U1165 ( .A1(n1684), .A2(wrdata_d1[139]), .A3(n2), .A4(n1047), .Y(
        n3471) );
  AO22X1_RVT U1166 ( .A1(n1742), .A2(\inq_ary[3][25] ), .A3(n1711), .A4(
        \inq_ary[13][25] ), .Y(n1051) );
  AO22X1_RVT U1167 ( .A1(n1729), .A2(\inq_ary[4][25] ), .A3(n1749), .A4(
        \inq_ary[1][25] ), .Y(n1050) );
  AO22X1_RVT U1168 ( .A1(n1747), .A2(\inq_ary[5][25] ), .A3(n1748), .A4(
        \inq_ary[10][25] ), .Y(n1049) );
  AO22X1_RVT U1169 ( .A1(n1612), .A2(\inq_ary[8][25] ), .A3(n1751), .A4(
        \inq_ary[9][25] ), .Y(n1048) );
  NOR4X1_RVT U1170 ( .A1(n1051), .A2(n1050), .A3(n1049), .A4(n1048), .Y(n1057)
         );
  AO22X1_RVT U1171 ( .A1(n1686), .A2(\inq_ary[0][25] ), .A3(n1537), .A4(
        \inq_ary[15][25] ), .Y(n1055) );
  AO22X1_RVT U1172 ( .A1(n1554), .A2(\inq_ary[14][25] ), .A3(n1750), .A4(
        \inq_ary[11][25] ), .Y(n1054) );
  AO22X1_RVT U1173 ( .A1(n1739), .A2(\inq_ary[2][25] ), .A3(n1740), .A4(
        \inq_ary[12][25] ), .Y(n1053) );
  AO22X1_RVT U1174 ( .A1(n1741), .A2(\inq_ary[7][25] ), .A3(n1738), .A4(
        \inq_ary[6][25] ), .Y(n1052) );
  NOR4X1_RVT U1175 ( .A1(n1055), .A2(n1054), .A3(n1053), .A4(n1052), .Y(n1056)
         );
  NAND2X0_RVT U1176 ( .A1(n1057), .A2(n1056), .Y(n1058) );
  AO22X1_RVT U1177 ( .A1(n3), .A2(wrdata_d1[25]), .A3(n1489), .A4(n1058), .Y(
        n3362) );
  AO22X1_RVT U1178 ( .A1(n1741), .A2(\inq_ary[7][10] ), .A3(n1711), .A4(
        \inq_ary[13][10] ), .Y(n1062) );
  AO22X1_RVT U1179 ( .A1(n1537), .A2(\inq_ary[15][10] ), .A3(n1738), .A4(
        \inq_ary[6][10] ), .Y(n1061) );
  AO22X1_RVT U1180 ( .A1(n1686), .A2(\inq_ary[0][10] ), .A3(n1751), .A4(
        \inq_ary[9][10] ), .Y(n1060) );
  AO22X1_RVT U1181 ( .A1(n1554), .A2(\inq_ary[14][10] ), .A3(n1747), .A4(
        \inq_ary[5][10] ), .Y(n1059) );
  NOR4X1_RVT U1182 ( .A1(n1062), .A2(n1061), .A3(n1060), .A4(n1059), .Y(n1068)
         );
  AO22X1_RVT U1183 ( .A1(n1742), .A2(\inq_ary[3][10] ), .A3(n1748), .A4(
        \inq_ary[10][10] ), .Y(n1066) );
  AO22X1_RVT U1184 ( .A1(n1612), .A2(\inq_ary[8][10] ), .A3(n1750), .A4(
        \inq_ary[11][10] ), .Y(n1065) );
  AO22X1_RVT U1185 ( .A1(n1739), .A2(\inq_ary[2][10] ), .A3(n1740), .A4(
        \inq_ary[12][10] ), .Y(n1064) );
  AO22X1_RVT U1186 ( .A1(n1729), .A2(\inq_ary[4][10] ), .A3(n1749), .A4(
        \inq_ary[1][10] ), .Y(n1063) );
  NOR4X1_RVT U1187 ( .A1(n1066), .A2(n1065), .A3(n1064), .A4(n1063), .Y(n1067)
         );
  NAND2X0_RVT U1188 ( .A1(n1068), .A2(n1067), .Y(n1069) );
  AO22X1_RVT U1189 ( .A1(n758), .A2(wrdata_d1[10]), .A3(n1), .A4(n1069), .Y(
        n3348) );
  AO22X1_RVT U1190 ( .A1(n1686), .A2(\inq_ary[0][140] ), .A3(n1751), .A4(
        \inq_ary[9][140] ), .Y(n1073) );
  AO22X1_RVT U1191 ( .A1(n1742), .A2(\inq_ary[3][140] ), .A3(n1612), .A4(
        \inq_ary[8][140] ), .Y(n1072) );
  AO22X1_RVT U1192 ( .A1(n1554), .A2(\inq_ary[14][140] ), .A3(n1711), .A4(
        \inq_ary[13][140] ), .Y(n1071) );
  AO22X1_RVT U1193 ( .A1(n1747), .A2(\inq_ary[5][140] ), .A3(n1738), .A4(
        \inq_ary[6][140] ), .Y(n1070) );
  NOR4X1_RVT U1194 ( .A1(n1073), .A2(n1072), .A3(n1071), .A4(n1070), .Y(n1079)
         );
  AO22X1_RVT U1195 ( .A1(n1741), .A2(\inq_ary[7][140] ), .A3(n1750), .A4(
        \inq_ary[11][140] ), .Y(n1077) );
  AO22X1_RVT U1196 ( .A1(n1739), .A2(\inq_ary[2][140] ), .A3(n1740), .A4(
        \inq_ary[12][140] ), .Y(n1076) );
  AO22X1_RVT U1197 ( .A1(n1537), .A2(\inq_ary[15][140] ), .A3(n1749), .A4(
        \inq_ary[1][140] ), .Y(n1075) );
  AO22X1_RVT U1198 ( .A1(n1729), .A2(\inq_ary[4][140] ), .A3(n1748), .A4(
        \inq_ary[10][140] ), .Y(n1074) );
  NOR4X1_RVT U1199 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .Y(n1078)
         );
  NAND2X0_RVT U1200 ( .A1(n1079), .A2(n1078), .Y(n1080) );
  AO22X1_RVT U1201 ( .A1(n3), .A2(wrdata_d1[140]), .A3(n1489), .A4(n1080), .Y(
        n3464) );
  AO22X1_RVT U1202 ( .A1(n1686), .A2(\inq_ary[0][21] ), .A3(n1612), .A4(
        \inq_ary[8][21] ), .Y(n1084) );
  AO22X1_RVT U1203 ( .A1(n1739), .A2(\inq_ary[2][21] ), .A3(n1747), .A4(
        \inq_ary[5][21] ), .Y(n1083) );
  AO22X1_RVT U1204 ( .A1(n1537), .A2(\inq_ary[15][21] ), .A3(n1738), .A4(
        \inq_ary[6][21] ), .Y(n1082) );
  AO22X1_RVT U1205 ( .A1(n1750), .A2(\inq_ary[11][21] ), .A3(n1751), .A4(
        \inq_ary[9][21] ), .Y(n1081) );
  NOR4X1_RVT U1206 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .Y(n1090)
         );
  AO22X1_RVT U1207 ( .A1(n1554), .A2(\inq_ary[14][21] ), .A3(n1729), .A4(
        \inq_ary[4][21] ), .Y(n1088) );
  AO22X1_RVT U1208 ( .A1(n1740), .A2(\inq_ary[12][21] ), .A3(n1741), .A4(
        \inq_ary[7][21] ), .Y(n1087) );
  AO22X1_RVT U1209 ( .A1(n1749), .A2(\inq_ary[1][21] ), .A3(n1711), .A4(
        \inq_ary[13][21] ), .Y(n1086) );
  AO22X1_RVT U1210 ( .A1(n1742), .A2(\inq_ary[3][21] ), .A3(n1748), .A4(
        \inq_ary[10][21] ), .Y(n1085) );
  NOR4X1_RVT U1211 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .Y(n1089)
         );
  NAND2X0_RVT U1212 ( .A1(n1090), .A2(n1089), .Y(n1091) );
  AO22X1_RVT U1213 ( .A1(n1025), .A2(wrdata_d1[21]), .A3(n1489), .A4(n1091), 
        .Y(n3353) );
  AO22X1_RVT U1214 ( .A1(n1729), .A2(\inq_ary[4][18] ), .A3(n1738), .A4(
        \inq_ary[6][18] ), .Y(n1095) );
  AO22X1_RVT U1215 ( .A1(n1739), .A2(\inq_ary[2][18] ), .A3(n1711), .A4(
        \inq_ary[13][18] ), .Y(n1094) );
  AO22X1_RVT U1216 ( .A1(n1748), .A2(\inq_ary[10][18] ), .A3(n1751), .A4(
        \inq_ary[9][18] ), .Y(n1093) );
  AO22X1_RVT U1217 ( .A1(n1742), .A2(\inq_ary[3][18] ), .A3(n1747), .A4(
        \inq_ary[5][18] ), .Y(n1092) );
  NOR4X1_RVT U1218 ( .A1(n1095), .A2(n1094), .A3(n1093), .A4(n1092), .Y(n1101)
         );
  AO22X1_RVT U1219 ( .A1(n1686), .A2(\inq_ary[0][18] ), .A3(n1537), .A4(
        \inq_ary[15][18] ), .Y(n1099) );
  AO22X1_RVT U1220 ( .A1(n1740), .A2(\inq_ary[12][18] ), .A3(n1749), .A4(
        \inq_ary[1][18] ), .Y(n1098) );
  AO22X1_RVT U1221 ( .A1(n1612), .A2(\inq_ary[8][18] ), .A3(n1750), .A4(
        \inq_ary[11][18] ), .Y(n1097) );
  AO22X1_RVT U1222 ( .A1(n1554), .A2(\inq_ary[14][18] ), .A3(n1741), .A4(
        \inq_ary[7][18] ), .Y(n1096) );
  NOR4X1_RVT U1223 ( .A1(n1099), .A2(n1098), .A3(n1097), .A4(n1096), .Y(n1100)
         );
  NAND2X0_RVT U1224 ( .A1(n1101), .A2(n1100), .Y(n1102) );
  AO22X1_RVT U1225 ( .A1(n1477), .A2(wrdata_d1[18]), .A3(n1), .A4(n1102), .Y(
        n3356) );
  AO22X1_RVT U1226 ( .A1(n1686), .A2(\inq_ary[0][19] ), .A3(n1750), .A4(
        \inq_ary[11][19] ), .Y(n1106) );
  AO22X1_RVT U1227 ( .A1(n1742), .A2(\inq_ary[3][19] ), .A3(n1612), .A4(
        \inq_ary[8][19] ), .Y(n1105) );
  AO22X1_RVT U1228 ( .A1(n1739), .A2(\inq_ary[2][19] ), .A3(n1711), .A4(
        \inq_ary[13][19] ), .Y(n1104) );
  AO22X1_RVT U1229 ( .A1(n1740), .A2(\inq_ary[12][19] ), .A3(n1747), .A4(
        \inq_ary[5][19] ), .Y(n1103) );
  NOR4X1_RVT U1230 ( .A1(n1106), .A2(n1105), .A3(n1104), .A4(n1103), .Y(n1112)
         );
  AO22X1_RVT U1231 ( .A1(n1729), .A2(\inq_ary[4][19] ), .A3(n1741), .A4(
        \inq_ary[7][19] ), .Y(n1110) );
  AO22X1_RVT U1232 ( .A1(n1537), .A2(\inq_ary[15][19] ), .A3(n1751), .A4(
        \inq_ary[9][19] ), .Y(n1109) );
  AO22X1_RVT U1233 ( .A1(n1738), .A2(\inq_ary[6][19] ), .A3(n1748), .A4(
        \inq_ary[10][19] ), .Y(n1108) );
  AO22X1_RVT U1234 ( .A1(n1554), .A2(\inq_ary[14][19] ), .A3(n1749), .A4(
        \inq_ary[1][19] ), .Y(n1107) );
  NOR4X1_RVT U1235 ( .A1(n1110), .A2(n1109), .A3(n1108), .A4(n1107), .Y(n1111)
         );
  NAND2X0_RVT U1236 ( .A1(n1112), .A2(n1111), .Y(n1113) );
  AO22X1_RVT U1237 ( .A1(n3), .A2(wrdata_d1[19]), .A3(n1), .A4(n1113), .Y(
        n3358) );
  AO22X1_RVT U1238 ( .A1(n1686), .A2(\inq_ary[0][20] ), .A3(n1750), .A4(
        \inq_ary[11][20] ), .Y(n1117) );
  AO22X1_RVT U1239 ( .A1(n1749), .A2(\inq_ary[1][20] ), .A3(n1711), .A4(
        \inq_ary[13][20] ), .Y(n1116) );
  AO22X1_RVT U1240 ( .A1(n1739), .A2(\inq_ary[2][20] ), .A3(n1751), .A4(
        \inq_ary[9][20] ), .Y(n1115) );
  AO22X1_RVT U1241 ( .A1(n1554), .A2(\inq_ary[14][20] ), .A3(n1729), .A4(
        \inq_ary[4][20] ), .Y(n1114) );
  NOR4X1_RVT U1242 ( .A1(n1117), .A2(n1116), .A3(n1115), .A4(n1114), .Y(n1123)
         );
  AO22X1_RVT U1243 ( .A1(n1742), .A2(\inq_ary[3][20] ), .A3(n1748), .A4(
        \inq_ary[10][20] ), .Y(n1121) );
  AO22X1_RVT U1244 ( .A1(n1740), .A2(\inq_ary[12][20] ), .A3(n1747), .A4(
        \inq_ary[5][20] ), .Y(n1120) );
  AO22X1_RVT U1245 ( .A1(n1537), .A2(\inq_ary[15][20] ), .A3(n1741), .A4(
        \inq_ary[7][20] ), .Y(n1119) );
  AO22X1_RVT U1246 ( .A1(n1612), .A2(\inq_ary[8][20] ), .A3(n1738), .A4(
        \inq_ary[6][20] ), .Y(n1118) );
  NOR4X1_RVT U1247 ( .A1(n1121), .A2(n1120), .A3(n1119), .A4(n1118), .Y(n1122)
         );
  NAND2X0_RVT U1248 ( .A1(n1123), .A2(n1122), .Y(n1124) );
  AO22X1_RVT U1249 ( .A1(n3), .A2(wrdata_d1[20]), .A3(n1), .A4(n1124), .Y(
        n3351) );
  AO22X1_RVT U1250 ( .A1(n1686), .A2(\inq_ary[0][13] ), .A3(n1740), .A4(
        \inq_ary[12][13] ), .Y(n1128) );
  AO22X1_RVT U1251 ( .A1(n1747), .A2(\inq_ary[5][13] ), .A3(n1738), .A4(
        \inq_ary[6][13] ), .Y(n1127) );
  AO22X1_RVT U1252 ( .A1(n1612), .A2(\inq_ary[8][13] ), .A3(n1741), .A4(
        \inq_ary[7][13] ), .Y(n1126) );
  AO22X1_RVT U1253 ( .A1(n1750), .A2(\inq_ary[11][13] ), .A3(n1748), .A4(
        \inq_ary[10][13] ), .Y(n1125) );
  NOR4X1_RVT U1254 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), .Y(n1134)
         );
  AO22X1_RVT U1255 ( .A1(n1749), .A2(\inq_ary[1][13] ), .A3(n1711), .A4(
        \inq_ary[13][13] ), .Y(n1132) );
  AO22X1_RVT U1256 ( .A1(n1739), .A2(\inq_ary[2][13] ), .A3(n1729), .A4(
        \inq_ary[4][13] ), .Y(n1131) );
  AO22X1_RVT U1257 ( .A1(n1554), .A2(\inq_ary[14][13] ), .A3(n1537), .A4(
        \inq_ary[15][13] ), .Y(n1130) );
  AO22X1_RVT U1258 ( .A1(n1742), .A2(\inq_ary[3][13] ), .A3(n1751), .A4(
        \inq_ary[9][13] ), .Y(n1129) );
  NOR4X1_RVT U1259 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .Y(n1133)
         );
  NAND2X0_RVT U1260 ( .A1(n1134), .A2(n1133), .Y(n1135) );
  AO22X1_RVT U1261 ( .A1(n758), .A2(wrdata_d1[13]), .A3(n1759), .A4(n1135), 
        .Y(n3345) );
  AO22X1_RVT U1262 ( .A1(n1738), .A2(\inq_ary[6][23] ), .A3(n1751), .A4(
        \inq_ary[9][23] ), .Y(n1139) );
  AO22X1_RVT U1263 ( .A1(n1729), .A2(\inq_ary[4][23] ), .A3(n1741), .A4(
        \inq_ary[7][23] ), .Y(n1138) );
  AO22X1_RVT U1264 ( .A1(n1742), .A2(\inq_ary[3][23] ), .A3(n1537), .A4(
        \inq_ary[15][23] ), .Y(n1137) );
  AO22X1_RVT U1265 ( .A1(n1747), .A2(\inq_ary[5][23] ), .A3(n1711), .A4(
        \inq_ary[13][23] ), .Y(n1136) );
  NOR4X1_RVT U1266 ( .A1(n1139), .A2(n1138), .A3(n1137), .A4(n1136), .Y(n1145)
         );
  AO22X1_RVT U1267 ( .A1(n1739), .A2(\inq_ary[2][23] ), .A3(n1554), .A4(
        \inq_ary[14][23] ), .Y(n1143) );
  AO22X1_RVT U1268 ( .A1(n1740), .A2(\inq_ary[12][23] ), .A3(n1750), .A4(
        \inq_ary[11][23] ), .Y(n1142) );
  AO22X1_RVT U1269 ( .A1(n1686), .A2(\inq_ary[0][23] ), .A3(n1748), .A4(
        \inq_ary[10][23] ), .Y(n1141) );
  AO22X1_RVT U1270 ( .A1(n1612), .A2(\inq_ary[8][23] ), .A3(n1749), .A4(
        \inq_ary[1][23] ), .Y(n1140) );
  NOR4X1_RVT U1271 ( .A1(n1143), .A2(n1142), .A3(n1141), .A4(n1140), .Y(n1144)
         );
  NAND2X0_RVT U1272 ( .A1(n1145), .A2(n1144), .Y(n1146) );
  AO22X1_RVT U1273 ( .A1(n1723), .A2(wrdata_d1[23]), .A3(n1759), .A4(n1146), 
        .Y(n3357) );
  AO22X1_RVT U1274 ( .A1(n1748), .A2(\inq_ary[10][14] ), .A3(n1751), .A4(
        \inq_ary[9][14] ), .Y(n1150) );
  AO22X1_RVT U1275 ( .A1(n1742), .A2(\inq_ary[3][14] ), .A3(n1711), .A4(
        \inq_ary[13][14] ), .Y(n1149) );
  AO22X1_RVT U1276 ( .A1(n1554), .A2(\inq_ary[14][14] ), .A3(n1741), .A4(
        \inq_ary[7][14] ), .Y(n1148) );
  AO22X1_RVT U1277 ( .A1(n1740), .A2(\inq_ary[12][14] ), .A3(n1738), .A4(
        \inq_ary[6][14] ), .Y(n1147) );
  NOR4X1_RVT U1278 ( .A1(n1150), .A2(n1149), .A3(n1148), .A4(n1147), .Y(n1156)
         );
  AO22X1_RVT U1279 ( .A1(n1686), .A2(\inq_ary[0][14] ), .A3(n1749), .A4(
        \inq_ary[1][14] ), .Y(n1154) );
  AO22X1_RVT U1280 ( .A1(n1537), .A2(\inq_ary[15][14] ), .A3(n1747), .A4(
        \inq_ary[5][14] ), .Y(n1153) );
  AO22X1_RVT U1281 ( .A1(n1739), .A2(\inq_ary[2][14] ), .A3(n1750), .A4(
        \inq_ary[11][14] ), .Y(n1152) );
  AO22X1_RVT U1282 ( .A1(n1729), .A2(\inq_ary[4][14] ), .A3(n1612), .A4(
        \inq_ary[8][14] ), .Y(n1151) );
  NOR4X1_RVT U1283 ( .A1(n1154), .A2(n1153), .A3(n1152), .A4(n1151), .Y(n1155)
         );
  NAND2X0_RVT U1284 ( .A1(n1156), .A2(n1155), .Y(n1157) );
  AO22X1_RVT U1285 ( .A1(n1760), .A2(wrdata_d1[14]), .A3(n969), .A4(n1157), 
        .Y(n3347) );
  AO22X1_RVT U1286 ( .A1(n1749), .A2(\inq_ary[1][147] ), .A3(n1747), .A4(
        \inq_ary[5][147] ), .Y(n1161) );
  AO22X1_RVT U1287 ( .A1(n1686), .A2(\inq_ary[0][147] ), .A3(n1612), .A4(
        \inq_ary[8][147] ), .Y(n1160) );
  AO22X1_RVT U1288 ( .A1(n1742), .A2(\inq_ary[3][147] ), .A3(n1729), .A4(
        \inq_ary[4][147] ), .Y(n1159) );
  AO22X1_RVT U1289 ( .A1(n1739), .A2(\inq_ary[2][147] ), .A3(n1711), .A4(
        \inq_ary[13][147] ), .Y(n1158) );
  NOR4X1_RVT U1290 ( .A1(n1161), .A2(n1160), .A3(n1159), .A4(n1158), .Y(n1167)
         );
  AO22X1_RVT U1291 ( .A1(n1740), .A2(\inq_ary[12][147] ), .A3(n1738), .A4(
        \inq_ary[6][147] ), .Y(n1165) );
  AO22X1_RVT U1292 ( .A1(n1554), .A2(\inq_ary[14][147] ), .A3(n1741), .A4(
        \inq_ary[7][147] ), .Y(n1164) );
  AO22X1_RVT U1293 ( .A1(n1750), .A2(\inq_ary[11][147] ), .A3(n1748), .A4(
        \inq_ary[10][147] ), .Y(n1163) );
  AO22X1_RVT U1294 ( .A1(n1537), .A2(\inq_ary[15][147] ), .A3(n1751), .A4(
        \inq_ary[9][147] ), .Y(n1162) );
  NOR4X1_RVT U1295 ( .A1(n1165), .A2(n1164), .A3(n1163), .A4(n1162), .Y(n1166)
         );
  NAND2X0_RVT U1296 ( .A1(n1167), .A2(n1166), .Y(n1168) );
  AO22X1_RVT U1297 ( .A1(n1723), .A2(wrdata_d1[147]), .A3(n1759), .A4(n1168), 
        .Y(n3475) );
  AO22X1_RVT U1298 ( .A1(n1537), .A2(\inq_ary[15][15] ), .A3(n1747), .A4(
        \inq_ary[5][15] ), .Y(n1172) );
  AO22X1_RVT U1299 ( .A1(n1742), .A2(\inq_ary[3][15] ), .A3(n1749), .A4(
        \inq_ary[1][15] ), .Y(n1171) );
  AO22X1_RVT U1300 ( .A1(n1729), .A2(\inq_ary[4][15] ), .A3(n1741), .A4(
        \inq_ary[7][15] ), .Y(n1170) );
  AO22X1_RVT U1301 ( .A1(n1612), .A2(\inq_ary[8][15] ), .A3(n1740), .A4(
        \inq_ary[12][15] ), .Y(n1169) );
  NOR4X1_RVT U1302 ( .A1(n1172), .A2(n1171), .A3(n1170), .A4(n1169), .Y(n1178)
         );
  AO22X1_RVT U1303 ( .A1(n1739), .A2(\inq_ary[2][15] ), .A3(n1711), .A4(
        \inq_ary[13][15] ), .Y(n1176) );
  AO22X1_RVT U1304 ( .A1(n1686), .A2(\inq_ary[0][15] ), .A3(n1748), .A4(
        \inq_ary[10][15] ), .Y(n1175) );
  AO22X1_RVT U1305 ( .A1(n1554), .A2(\inq_ary[14][15] ), .A3(n1738), .A4(
        \inq_ary[6][15] ), .Y(n1174) );
  AO22X1_RVT U1306 ( .A1(n1750), .A2(\inq_ary[11][15] ), .A3(n1751), .A4(
        \inq_ary[9][15] ), .Y(n1173) );
  NOR4X1_RVT U1307 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), .Y(n1177)
         );
  NAND2X0_RVT U1308 ( .A1(n1178), .A2(n1177), .Y(n1179) );
  AO22X1_RVT U1309 ( .A1(n1684), .A2(wrdata_d1[15]), .A3(n2), .A4(n1179), .Y(
        n3349) );
  AO22X1_RVT U1310 ( .A1(n1749), .A2(\inq_ary[1][22] ), .A3(n1750), .A4(
        \inq_ary[11][22] ), .Y(n1183) );
  AO22X1_RVT U1311 ( .A1(n1747), .A2(\inq_ary[5][22] ), .A3(n1738), .A4(
        \inq_ary[6][22] ), .Y(n1182) );
  AO22X1_RVT U1312 ( .A1(n1742), .A2(\inq_ary[3][22] ), .A3(n1748), .A4(
        \inq_ary[10][22] ), .Y(n1181) );
  AO22X1_RVT U1313 ( .A1(n1537), .A2(\inq_ary[15][22] ), .A3(n1751), .A4(
        \inq_ary[9][22] ), .Y(n1180) );
  NOR4X1_RVT U1314 ( .A1(n1183), .A2(n1182), .A3(n1181), .A4(n1180), .Y(n1189)
         );
  AO22X1_RVT U1315 ( .A1(n1729), .A2(\inq_ary[4][22] ), .A3(n1711), .A4(
        \inq_ary[13][22] ), .Y(n1187) );
  AO22X1_RVT U1316 ( .A1(n1612), .A2(\inq_ary[8][22] ), .A3(n1740), .A4(
        \inq_ary[12][22] ), .Y(n1186) );
  AO22X1_RVT U1317 ( .A1(n1739), .A2(\inq_ary[2][22] ), .A3(n1554), .A4(
        \inq_ary[14][22] ), .Y(n1185) );
  AO22X1_RVT U1318 ( .A1(n1686), .A2(\inq_ary[0][22] ), .A3(n1741), .A4(
        \inq_ary[7][22] ), .Y(n1184) );
  NOR4X1_RVT U1319 ( .A1(n1187), .A2(n1186), .A3(n1185), .A4(n1184), .Y(n1188)
         );
  NAND2X0_RVT U1320 ( .A1(n1189), .A2(n1188), .Y(n1190) );
  AO22X1_RVT U1321 ( .A1(n1598), .A2(wrdata_d1[22]), .A3(n1759), .A4(n1190), 
        .Y(n3355) );
  AO22X1_RVT U1322 ( .A1(n1686), .A2(\inq_ary[0][16] ), .A3(n1741), .A4(
        \inq_ary[7][16] ), .Y(n1194) );
  AO22X1_RVT U1323 ( .A1(n1729), .A2(\inq_ary[4][16] ), .A3(n1738), .A4(
        \inq_ary[6][16] ), .Y(n1193) );
  AO22X1_RVT U1324 ( .A1(n1739), .A2(\inq_ary[2][16] ), .A3(n1747), .A4(
        \inq_ary[5][16] ), .Y(n1192) );
  AO22X1_RVT U1325 ( .A1(n1740), .A2(\inq_ary[12][16] ), .A3(n1749), .A4(
        \inq_ary[1][16] ), .Y(n1191) );
  NOR4X1_RVT U1326 ( .A1(n1194), .A2(n1193), .A3(n1192), .A4(n1191), .Y(n1200)
         );
  AO22X1_RVT U1327 ( .A1(n1554), .A2(\inq_ary[14][16] ), .A3(n1537), .A4(
        \inq_ary[15][16] ), .Y(n1198) );
  AO22X1_RVT U1328 ( .A1(n1742), .A2(\inq_ary[3][16] ), .A3(n1711), .A4(
        \inq_ary[13][16] ), .Y(n1197) );
  AO22X1_RVT U1329 ( .A1(n1612), .A2(\inq_ary[8][16] ), .A3(n1750), .A4(
        \inq_ary[11][16] ), .Y(n1196) );
  AO22X1_RVT U1330 ( .A1(n1748), .A2(\inq_ary[10][16] ), .A3(n1751), .A4(
        \inq_ary[9][16] ), .Y(n1195) );
  NOR4X1_RVT U1331 ( .A1(n1198), .A2(n1197), .A3(n1196), .A4(n1195), .Y(n1199)
         );
  NAND2X0_RVT U1332 ( .A1(n1200), .A2(n1199), .Y(n1201) );
  AO22X1_RVT U1333 ( .A1(n1684), .A2(wrdata_d1[16]), .A3(n946), .A4(n1201), 
        .Y(n3352) );
  AO22X1_RVT U1334 ( .A1(n1554), .A2(\inq_ary[14][17] ), .A3(n1537), .A4(
        \inq_ary[15][17] ), .Y(n1205) );
  AO22X1_RVT U1335 ( .A1(n1686), .A2(\inq_ary[0][17] ), .A3(n1748), .A4(
        \inq_ary[10][17] ), .Y(n1204) );
  AO22X1_RVT U1336 ( .A1(n1739), .A2(\inq_ary[2][17] ), .A3(n1711), .A4(
        \inq_ary[13][17] ), .Y(n1203) );
  AO22X1_RVT U1337 ( .A1(n1729), .A2(\inq_ary[4][17] ), .A3(n1750), .A4(
        \inq_ary[11][17] ), .Y(n1202) );
  NOR4X1_RVT U1338 ( .A1(n1205), .A2(n1204), .A3(n1203), .A4(n1202), .Y(n1211)
         );
  AO22X1_RVT U1339 ( .A1(n1740), .A2(\inq_ary[12][17] ), .A3(n1751), .A4(
        \inq_ary[9][17] ), .Y(n1209) );
  AO22X1_RVT U1340 ( .A1(n1749), .A2(\inq_ary[1][17] ), .A3(n1738), .A4(
        \inq_ary[6][17] ), .Y(n1208) );
  AO22X1_RVT U1341 ( .A1(n1742), .A2(\inq_ary[3][17] ), .A3(n1747), .A4(
        \inq_ary[5][17] ), .Y(n1207) );
  AO22X1_RVT U1342 ( .A1(n1612), .A2(\inq_ary[8][17] ), .A3(n1741), .A4(
        \inq_ary[7][17] ), .Y(n1206) );
  NOR4X1_RVT U1343 ( .A1(n1209), .A2(n1208), .A3(n1207), .A4(n1206), .Y(n1210)
         );
  NAND2X0_RVT U1344 ( .A1(n1211), .A2(n1210), .Y(n1212) );
  AO22X1_RVT U1345 ( .A1(n758), .A2(wrdata_d1[17]), .A3(n2), .A4(n1212), .Y(
        n3354) );
  AO22X1_RVT U1346 ( .A1(n1554), .A2(\inq_ary[14][129] ), .A3(n1612), .A4(
        \inq_ary[8][129] ), .Y(n1216) );
  AO22X1_RVT U1347 ( .A1(n1740), .A2(\inq_ary[12][129] ), .A3(n1750), .A4(
        \inq_ary[11][129] ), .Y(n1215) );
  AO22X1_RVT U1348 ( .A1(n1686), .A2(\inq_ary[0][129] ), .A3(n1738), .A4(
        \inq_ary[6][129] ), .Y(n1214) );
  AO22X1_RVT U1349 ( .A1(n1747), .A2(\inq_ary[5][129] ), .A3(n1748), .A4(
        \inq_ary[10][129] ), .Y(n1213) );
  NOR4X1_RVT U1350 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), .Y(n1222)
         );
  AO22X1_RVT U1351 ( .A1(n1742), .A2(\inq_ary[3][129] ), .A3(n1741), .A4(
        \inq_ary[7][129] ), .Y(n1220) );
  AO22X1_RVT U1352 ( .A1(n1729), .A2(\inq_ary[4][129] ), .A3(n1711), .A4(
        \inq_ary[13][129] ), .Y(n1219) );
  AO22X1_RVT U1353 ( .A1(n1739), .A2(\inq_ary[2][129] ), .A3(n1751), .A4(
        \inq_ary[9][129] ), .Y(n1218) );
  AO22X1_RVT U1354 ( .A1(n1537), .A2(\inq_ary[15][129] ), .A3(n1749), .A4(
        \inq_ary[1][129] ), .Y(n1217) );
  NOR4X1_RVT U1355 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), .Y(n1221)
         );
  NAND2X0_RVT U1356 ( .A1(n1222), .A2(n1221), .Y(n1223) );
  AO22X1_RVT U1357 ( .A1(n1025), .A2(wrdata_d1[129]), .A3(n1489), .A4(n1223), 
        .Y(n3459) );
  AO22X1_RVT U1358 ( .A1(n1686), .A2(\inq_ary[0][126] ), .A3(n1749), .A4(
        \inq_ary[1][126] ), .Y(n1227) );
  AO22X1_RVT U1359 ( .A1(n1612), .A2(\inq_ary[8][126] ), .A3(n1750), .A4(
        \inq_ary[11][126] ), .Y(n1226) );
  AO22X1_RVT U1360 ( .A1(n1740), .A2(\inq_ary[12][126] ), .A3(n1748), .A4(
        \inq_ary[10][126] ), .Y(n1225) );
  AO22X1_RVT U1361 ( .A1(n1742), .A2(\inq_ary[3][126] ), .A3(n1741), .A4(
        \inq_ary[7][126] ), .Y(n1224) );
  NOR4X1_RVT U1362 ( .A1(n1227), .A2(n1226), .A3(n1225), .A4(n1224), .Y(n1233)
         );
  AO22X1_RVT U1363 ( .A1(n1739), .A2(\inq_ary[2][126] ), .A3(n1711), .A4(
        \inq_ary[13][126] ), .Y(n1231) );
  AO22X1_RVT U1364 ( .A1(n1554), .A2(\inq_ary[14][126] ), .A3(n1729), .A4(
        \inq_ary[4][126] ), .Y(n1230) );
  AO22X1_RVT U1365 ( .A1(n1537), .A2(\inq_ary[15][126] ), .A3(n1751), .A4(
        \inq_ary[9][126] ), .Y(n1229) );
  AO22X1_RVT U1366 ( .A1(n1747), .A2(\inq_ary[5][126] ), .A3(n1738), .A4(
        \inq_ary[6][126] ), .Y(n1228) );
  NOR4X1_RVT U1367 ( .A1(n1231), .A2(n1230), .A3(n1229), .A4(n1228), .Y(n1232)
         );
  NAND2X0_RVT U1368 ( .A1(n1233), .A2(n1232), .Y(n1234) );
  AO22X1_RVT U1369 ( .A1(n1477), .A2(wrdata_d1[126]), .A3(n1), .A4(n1234), .Y(
        n3452) );
  AO22X1_RVT U1370 ( .A1(n1739), .A2(\inq_ary[2][121] ), .A3(n1750), .A4(
        \inq_ary[11][121] ), .Y(n1238) );
  AO22X1_RVT U1371 ( .A1(n1729), .A2(\inq_ary[4][121] ), .A3(n1749), .A4(
        \inq_ary[1][121] ), .Y(n1237) );
  AO22X1_RVT U1372 ( .A1(n1711), .A2(\inq_ary[13][121] ), .A3(n1748), .A4(
        \inq_ary[10][121] ), .Y(n1236) );
  AO22X1_RVT U1373 ( .A1(n1686), .A2(\inq_ary[0][121] ), .A3(n1751), .A4(
        \inq_ary[9][121] ), .Y(n1235) );
  NOR4X1_RVT U1374 ( .A1(n1238), .A2(n1237), .A3(n1236), .A4(n1235), .Y(n1244)
         );
  AO22X1_RVT U1375 ( .A1(n1554), .A2(\inq_ary[14][121] ), .A3(n1741), .A4(
        \inq_ary[7][121] ), .Y(n1242) );
  AO22X1_RVT U1376 ( .A1(n1612), .A2(\inq_ary[8][121] ), .A3(n1740), .A4(
        \inq_ary[12][121] ), .Y(n1241) );
  AO22X1_RVT U1377 ( .A1(n1537), .A2(\inq_ary[15][121] ), .A3(n1738), .A4(
        \inq_ary[6][121] ), .Y(n1240) );
  AO22X1_RVT U1378 ( .A1(n1742), .A2(\inq_ary[3][121] ), .A3(n1747), .A4(
        \inq_ary[5][121] ), .Y(n1239) );
  NOR4X1_RVT U1379 ( .A1(n1242), .A2(n1241), .A3(n1240), .A4(n1239), .Y(n1243)
         );
  NAND2X0_RVT U1380 ( .A1(n1244), .A2(n1243), .Y(n1245) );
  AO22X1_RVT U1381 ( .A1(n3), .A2(wrdata_d1[121]), .A3(n1), .A4(n1245), .Y(
        n3451) );
  AO22X1_RVT U1382 ( .A1(n1612), .A2(\inq_ary[8][127] ), .A3(n1748), .A4(
        \inq_ary[10][127] ), .Y(n1249) );
  AO22X1_RVT U1383 ( .A1(n1742), .A2(\inq_ary[3][127] ), .A3(n1741), .A4(
        \inq_ary[7][127] ), .Y(n1248) );
  AO22X1_RVT U1384 ( .A1(n1686), .A2(\inq_ary[0][127] ), .A3(n1749), .A4(
        \inq_ary[1][127] ), .Y(n1247) );
  AO22X1_RVT U1385 ( .A1(n1740), .A2(\inq_ary[12][127] ), .A3(n1747), .A4(
        \inq_ary[5][127] ), .Y(n1246) );
  NOR4X1_RVT U1386 ( .A1(n1249), .A2(n1248), .A3(n1247), .A4(n1246), .Y(n1255)
         );
  AO22X1_RVT U1387 ( .A1(n1739), .A2(\inq_ary[2][127] ), .A3(n1554), .A4(
        \inq_ary[14][127] ), .Y(n1253) );
  AO22X1_RVT U1388 ( .A1(n1537), .A2(\inq_ary[15][127] ), .A3(n1751), .A4(
        \inq_ary[9][127] ), .Y(n1252) );
  AO22X1_RVT U1389 ( .A1(n1729), .A2(\inq_ary[4][127] ), .A3(n1738), .A4(
        \inq_ary[6][127] ), .Y(n1251) );
  AO22X1_RVT U1390 ( .A1(n1750), .A2(\inq_ary[11][127] ), .A3(n1711), .A4(
        \inq_ary[13][127] ), .Y(n1250) );
  NOR4X1_RVT U1391 ( .A1(n1253), .A2(n1252), .A3(n1251), .A4(n1250), .Y(n1254)
         );
  NAND2X0_RVT U1392 ( .A1(n1255), .A2(n1254), .Y(n1256) );
  AO22X1_RVT U1393 ( .A1(n3), .A2(wrdata_d1[127]), .A3(n1489), .A4(n1256), .Y(
        n3454) );
  AO22X1_RVT U1394 ( .A1(n1554), .A2(\inq_ary[14][28] ), .A3(n1749), .A4(
        \inq_ary[1][28] ), .Y(n1260) );
  AO22X1_RVT U1395 ( .A1(n1747), .A2(\inq_ary[5][28] ), .A3(n1748), .A4(
        \inq_ary[10][28] ), .Y(n1259) );
  AO22X1_RVT U1396 ( .A1(n1686), .A2(\inq_ary[0][28] ), .A3(n1751), .A4(
        \inq_ary[9][28] ), .Y(n1258) );
  AO22X1_RVT U1397 ( .A1(n1739), .A2(\inq_ary[2][28] ), .A3(n1729), .A4(
        \inq_ary[4][28] ), .Y(n1257) );
  NOR4X1_RVT U1398 ( .A1(n1260), .A2(n1259), .A3(n1258), .A4(n1257), .Y(n1266)
         );
  AO22X1_RVT U1399 ( .A1(n1612), .A2(\inq_ary[8][28] ), .A3(n1750), .A4(
        \inq_ary[11][28] ), .Y(n1264) );
  AO22X1_RVT U1400 ( .A1(n1740), .A2(\inq_ary[12][28] ), .A3(n1741), .A4(
        \inq_ary[7][28] ), .Y(n1263) );
  AO22X1_RVT U1401 ( .A1(n1537), .A2(\inq_ary[15][28] ), .A3(n1738), .A4(
        \inq_ary[6][28] ), .Y(n1262) );
  AO22X1_RVT U1402 ( .A1(n1742), .A2(\inq_ary[3][28] ), .A3(n1711), .A4(
        \inq_ary[13][28] ), .Y(n1261) );
  NOR4X1_RVT U1403 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .Y(n1265)
         );
  NAND2X0_RVT U1404 ( .A1(n1266), .A2(n1265), .Y(n1267) );
  AO22X1_RVT U1405 ( .A1(n1723), .A2(wrdata_d1[28]), .A3(n969), .A4(n1267), 
        .Y(n3359) );
  AO22X1_RVT U1406 ( .A1(n1750), .A2(\inq_ary[11][125] ), .A3(n1711), .A4(
        \inq_ary[13][125] ), .Y(n1271) );
  AO22X1_RVT U1407 ( .A1(n1741), .A2(\inq_ary[7][125] ), .A3(n1751), .A4(
        \inq_ary[9][125] ), .Y(n1270) );
  AO22X1_RVT U1408 ( .A1(n1686), .A2(\inq_ary[0][125] ), .A3(n1738), .A4(
        \inq_ary[6][125] ), .Y(n1269) );
  AO22X1_RVT U1409 ( .A1(n1742), .A2(\inq_ary[3][125] ), .A3(n1748), .A4(
        \inq_ary[10][125] ), .Y(n1268) );
  NOR4X1_RVT U1410 ( .A1(n1271), .A2(n1270), .A3(n1269), .A4(n1268), .Y(n1277)
         );
  AO22X1_RVT U1411 ( .A1(n1612), .A2(\inq_ary[8][125] ), .A3(n1749), .A4(
        \inq_ary[1][125] ), .Y(n1275) );
  AO22X1_RVT U1412 ( .A1(n1739), .A2(\inq_ary[2][125] ), .A3(n1747), .A4(
        \inq_ary[5][125] ), .Y(n1274) );
  AO22X1_RVT U1413 ( .A1(n1537), .A2(\inq_ary[15][125] ), .A3(n1740), .A4(
        \inq_ary[12][125] ), .Y(n1273) );
  AO22X1_RVT U1414 ( .A1(n1554), .A2(\inq_ary[14][125] ), .A3(n1729), .A4(
        \inq_ary[4][125] ), .Y(n1272) );
  NOR4X1_RVT U1415 ( .A1(n1275), .A2(n1274), .A3(n1273), .A4(n1272), .Y(n1276)
         );
  NAND2X0_RVT U1416 ( .A1(n1277), .A2(n1276), .Y(n1278) );
  AO22X1_RVT U1417 ( .A1(n1760), .A2(wrdata_d1[125]), .A3(n1), .A4(n1278), .Y(
        n3450) );
  AO22X1_RVT U1418 ( .A1(n1554), .A2(\inq_ary[14][120] ), .A3(n1750), .A4(
        \inq_ary[11][120] ), .Y(n1282) );
  AO22X1_RVT U1419 ( .A1(n1537), .A2(\inq_ary[15][120] ), .A3(n1738), .A4(
        \inq_ary[6][120] ), .Y(n1281) );
  AO22X1_RVT U1420 ( .A1(n1740), .A2(\inq_ary[12][120] ), .A3(n1711), .A4(
        \inq_ary[13][120] ), .Y(n1280) );
  AO22X1_RVT U1421 ( .A1(n1739), .A2(\inq_ary[2][120] ), .A3(n1741), .A4(
        \inq_ary[7][120] ), .Y(n1279) );
  NOR4X1_RVT U1422 ( .A1(n1282), .A2(n1281), .A3(n1280), .A4(n1279), .Y(n1288)
         );
  AO22X1_RVT U1423 ( .A1(n1742), .A2(\inq_ary[3][120] ), .A3(n1749), .A4(
        \inq_ary[1][120] ), .Y(n1286) );
  AO22X1_RVT U1424 ( .A1(n1747), .A2(\inq_ary[5][120] ), .A3(n1748), .A4(
        \inq_ary[10][120] ), .Y(n1285) );
  AO22X1_RVT U1425 ( .A1(n1729), .A2(\inq_ary[4][120] ), .A3(n1751), .A4(
        \inq_ary[9][120] ), .Y(n1284) );
  AO22X1_RVT U1426 ( .A1(n1686), .A2(\inq_ary[0][120] ), .A3(n1612), .A4(
        \inq_ary[8][120] ), .Y(n1283) );
  NOR4X1_RVT U1427 ( .A1(n1286), .A2(n1285), .A3(n1284), .A4(n1283), .Y(n1287)
         );
  NAND2X0_RVT U1428 ( .A1(n1288), .A2(n1287), .Y(n1289) );
  AO22X1_RVT U1429 ( .A1(n1684), .A2(wrdata_d1[120]), .A3(n1), .A4(n1289), .Y(
        n3449) );
  AO22X1_RVT U1430 ( .A1(n1686), .A2(\inq_ary[0][128] ), .A3(n1749), .A4(
        \inq_ary[1][128] ), .Y(n1293) );
  AO22X1_RVT U1431 ( .A1(n1729), .A2(\inq_ary[4][128] ), .A3(n1740), .A4(
        \inq_ary[12][128] ), .Y(n1292) );
  AO22X1_RVT U1432 ( .A1(n1537), .A2(\inq_ary[15][128] ), .A3(n1748), .A4(
        \inq_ary[10][128] ), .Y(n1291) );
  AO22X1_RVT U1433 ( .A1(n1554), .A2(\inq_ary[14][128] ), .A3(n1751), .A4(
        \inq_ary[9][128] ), .Y(n1290) );
  NOR4X1_RVT U1434 ( .A1(n1293), .A2(n1292), .A3(n1291), .A4(n1290), .Y(n1299)
         );
  AO22X1_RVT U1435 ( .A1(n1747), .A2(\inq_ary[5][128] ), .A3(n1738), .A4(
        \inq_ary[6][128] ), .Y(n1297) );
  AO22X1_RVT U1436 ( .A1(n1739), .A2(\inq_ary[2][128] ), .A3(n1612), .A4(
        \inq_ary[8][128] ), .Y(n1296) );
  AO22X1_RVT U1437 ( .A1(n1742), .A2(\inq_ary[3][128] ), .A3(n1750), .A4(
        \inq_ary[11][128] ), .Y(n1295) );
  AO22X1_RVT U1438 ( .A1(n1741), .A2(\inq_ary[7][128] ), .A3(n1711), .A4(
        \inq_ary[13][128] ), .Y(n1294) );
  NOR4X1_RVT U1439 ( .A1(n1297), .A2(n1296), .A3(n1295), .A4(n1294), .Y(n1298)
         );
  NAND2X0_RVT U1440 ( .A1(n1299), .A2(n1298), .Y(n1300) );
  AO22X1_RVT U1441 ( .A1(n1598), .A2(wrdata_d1[128]), .A3(n1489), .A4(n1300), 
        .Y(n3457) );
  AO22X1_RVT U1442 ( .A1(n1537), .A2(\inq_ary[15][29] ), .A3(n1740), .A4(
        \inq_ary[12][29] ), .Y(n1304) );
  AO22X1_RVT U1443 ( .A1(n1729), .A2(\inq_ary[4][29] ), .A3(n1738), .A4(
        \inq_ary[6][29] ), .Y(n1303) );
  AO22X1_RVT U1444 ( .A1(n1742), .A2(\inq_ary[3][29] ), .A3(n1748), .A4(
        \inq_ary[10][29] ), .Y(n1302) );
  AO22X1_RVT U1445 ( .A1(n1739), .A2(\inq_ary[2][29] ), .A3(n1711), .A4(
        \inq_ary[13][29] ), .Y(n1301) );
  NOR4X1_RVT U1446 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .Y(n1310)
         );
  AO22X1_RVT U1447 ( .A1(n1686), .A2(\inq_ary[0][29] ), .A3(n1741), .A4(
        \inq_ary[7][29] ), .Y(n1308) );
  AO22X1_RVT U1448 ( .A1(n1554), .A2(\inq_ary[14][29] ), .A3(n1751), .A4(
        \inq_ary[9][29] ), .Y(n1307) );
  AO22X1_RVT U1449 ( .A1(n1749), .A2(\inq_ary[1][29] ), .A3(n1747), .A4(
        \inq_ary[5][29] ), .Y(n1306) );
  AO22X1_RVT U1450 ( .A1(n1612), .A2(\inq_ary[8][29] ), .A3(n1750), .A4(
        \inq_ary[11][29] ), .Y(n1305) );
  NOR4X1_RVT U1451 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .Y(n1309)
         );
  NAND2X0_RVT U1452 ( .A1(n1310), .A2(n1309), .Y(n1311) );
  AO22X1_RVT U1453 ( .A1(n758), .A2(wrdata_d1[29]), .A3(n2), .A4(n1311), .Y(
        n3361) );
  AO22X1_RVT U1454 ( .A1(n1729), .A2(\inq_ary[4][132] ), .A3(n1612), .A4(
        \inq_ary[8][132] ), .Y(n1315) );
  AO22X1_RVT U1455 ( .A1(n1742), .A2(\inq_ary[3][132] ), .A3(n1750), .A4(
        \inq_ary[11][132] ), .Y(n1314) );
  AO22X1_RVT U1456 ( .A1(n1554), .A2(\inq_ary[14][132] ), .A3(n1537), .A4(
        \inq_ary[15][132] ), .Y(n1313) );
  AO22X1_RVT U1457 ( .A1(n1747), .A2(\inq_ary[5][132] ), .A3(n1711), .A4(
        \inq_ary[13][132] ), .Y(n1312) );
  NOR4X1_RVT U1458 ( .A1(n1315), .A2(n1314), .A3(n1313), .A4(n1312), .Y(n1321)
         );
  AO22X1_RVT U1459 ( .A1(n1686), .A2(\inq_ary[0][132] ), .A3(n1738), .A4(
        \inq_ary[6][132] ), .Y(n1319) );
  AO22X1_RVT U1460 ( .A1(n1740), .A2(\inq_ary[12][132] ), .A3(n1749), .A4(
        \inq_ary[1][132] ), .Y(n1318) );
  AO22X1_RVT U1461 ( .A1(n1741), .A2(\inq_ary[7][132] ), .A3(n1751), .A4(
        \inq_ary[9][132] ), .Y(n1317) );
  AO22X1_RVT U1462 ( .A1(n1739), .A2(\inq_ary[2][132] ), .A3(n1748), .A4(
        \inq_ary[10][132] ), .Y(n1316) );
  NOR4X1_RVT U1463 ( .A1(n1319), .A2(n1318), .A3(n1317), .A4(n1316), .Y(n1320)
         );
  NAND2X0_RVT U1464 ( .A1(n1321), .A2(n1320), .Y(n1322) );
  AO22X1_RVT U1465 ( .A1(n758), .A2(wrdata_d1[132]), .A3(n1489), .A4(n1322), 
        .Y(n3456) );
  AO22X1_RVT U1466 ( .A1(n1729), .A2(\inq_ary[4][133] ), .A3(n1741), .A4(
        \inq_ary[7][133] ), .Y(n1326) );
  AO22X1_RVT U1467 ( .A1(n1554), .A2(\inq_ary[14][133] ), .A3(n1747), .A4(
        \inq_ary[5][133] ), .Y(n1325) );
  AO22X1_RVT U1468 ( .A1(n1742), .A2(\inq_ary[3][133] ), .A3(n1711), .A4(
        \inq_ary[13][133] ), .Y(n1324) );
  AO22X1_RVT U1469 ( .A1(n1739), .A2(\inq_ary[2][133] ), .A3(n1612), .A4(
        \inq_ary[8][133] ), .Y(n1323) );
  NOR4X1_RVT U1470 ( .A1(n1326), .A2(n1325), .A3(n1324), .A4(n1323), .Y(n1332)
         );
  AO22X1_RVT U1471 ( .A1(n1749), .A2(\inq_ary[1][133] ), .A3(n1738), .A4(
        \inq_ary[6][133] ), .Y(n1330) );
  AO22X1_RVT U1472 ( .A1(n1686), .A2(\inq_ary[0][133] ), .A3(n1740), .A4(
        \inq_ary[12][133] ), .Y(n1329) );
  AO22X1_RVT U1473 ( .A1(n1537), .A2(\inq_ary[15][133] ), .A3(n1751), .A4(
        \inq_ary[9][133] ), .Y(n1328) );
  AO22X1_RVT U1474 ( .A1(n1750), .A2(\inq_ary[11][133] ), .A3(n1748), .A4(
        \inq_ary[10][133] ), .Y(n1327) );
  NOR4X1_RVT U1475 ( .A1(n1330), .A2(n1329), .A3(n1328), .A4(n1327), .Y(n1331)
         );
  NAND2X0_RVT U1476 ( .A1(n1332), .A2(n1331), .Y(n1333) );
  AO22X1_RVT U1477 ( .A1(n1025), .A2(wrdata_d1[133]), .A3(n1489), .A4(n1333), 
        .Y(n3458) );
  AO22X1_RVT U1478 ( .A1(n1612), .A2(\inq_ary[8][123] ), .A3(n1738), .A4(
        \inq_ary[6][123] ), .Y(n1337) );
  AO22X1_RVT U1479 ( .A1(n1750), .A2(\inq_ary[11][123] ), .A3(n1748), .A4(
        \inq_ary[10][123] ), .Y(n1336) );
  AO22X1_RVT U1480 ( .A1(n1742), .A2(\inq_ary[3][123] ), .A3(n1711), .A4(
        \inq_ary[13][123] ), .Y(n1335) );
  AO22X1_RVT U1481 ( .A1(n1741), .A2(\inq_ary[7][123] ), .A3(n1751), .A4(
        \inq_ary[9][123] ), .Y(n1334) );
  NOR4X1_RVT U1482 ( .A1(n1337), .A2(n1336), .A3(n1335), .A4(n1334), .Y(n1343)
         );
  AO22X1_RVT U1483 ( .A1(n1729), .A2(\inq_ary[4][123] ), .A3(n1749), .A4(
        \inq_ary[1][123] ), .Y(n1341) );
  AO22X1_RVT U1484 ( .A1(n1739), .A2(\inq_ary[2][123] ), .A3(n1747), .A4(
        \inq_ary[5][123] ), .Y(n1340) );
  AO22X1_RVT U1485 ( .A1(n1554), .A2(\inq_ary[14][123] ), .A3(n1740), .A4(
        \inq_ary[12][123] ), .Y(n1339) );
  AO22X1_RVT U1486 ( .A1(n1686), .A2(\inq_ary[0][123] ), .A3(n1537), .A4(
        \inq_ary[15][123] ), .Y(n1338) );
  NOR4X1_RVT U1487 ( .A1(n1341), .A2(n1340), .A3(n1339), .A4(n1338), .Y(n1342)
         );
  NAND2X0_RVT U1488 ( .A1(n1343), .A2(n1342), .Y(n1344) );
  AO22X1_RVT U1489 ( .A1(n1477), .A2(wrdata_d1[123]), .A3(n1489), .A4(n1344), 
        .Y(n3455) );
  AO22X1_RVT U1490 ( .A1(n1612), .A2(\inq_ary[8][7] ), .A3(n1748), .A4(
        \inq_ary[10][7] ), .Y(n1348) );
  AO22X1_RVT U1491 ( .A1(n1739), .A2(\inq_ary[2][7] ), .A3(n1554), .A4(
        \inq_ary[14][7] ), .Y(n1347) );
  AO22X1_RVT U1492 ( .A1(n1742), .A2(\inq_ary[3][7] ), .A3(n1747), .A4(
        \inq_ary[5][7] ), .Y(n1346) );
  AO22X1_RVT U1493 ( .A1(n1729), .A2(\inq_ary[4][7] ), .A3(n1740), .A4(
        \inq_ary[12][7] ), .Y(n1345) );
  NOR4X1_RVT U1494 ( .A1(n1348), .A2(n1347), .A3(n1346), .A4(n1345), .Y(n1354)
         );
  AO22X1_RVT U1495 ( .A1(n1537), .A2(\inq_ary[15][7] ), .A3(n1711), .A4(
        \inq_ary[13][7] ), .Y(n1352) );
  AO22X1_RVT U1496 ( .A1(n1749), .A2(\inq_ary[1][7] ), .A3(n1750), .A4(
        \inq_ary[11][7] ), .Y(n1351) );
  AO22X1_RVT U1497 ( .A1(n1741), .A2(\inq_ary[7][7] ), .A3(n1738), .A4(
        \inq_ary[6][7] ), .Y(n1350) );
  AO22X1_RVT U1498 ( .A1(n1686), .A2(\inq_ary[0][7] ), .A3(n1751), .A4(
        \inq_ary[9][7] ), .Y(n1349) );
  NOR4X1_RVT U1499 ( .A1(n1352), .A2(n1351), .A3(n1350), .A4(n1349), .Y(n1353)
         );
  NAND2X0_RVT U1500 ( .A1(n1354), .A2(n1353), .Y(n1355) );
  AO22X1_RVT U1501 ( .A1(n3), .A2(wrdata_d1[7]), .A3(n1489), .A4(n1355), .Y(
        n3342) );
  AO22X1_RVT U1502 ( .A1(n1739), .A2(\inq_ary[2][117] ), .A3(n1747), .A4(
        \inq_ary[5][117] ), .Y(n1359) );
  AO22X1_RVT U1503 ( .A1(n1749), .A2(\inq_ary[1][117] ), .A3(n1748), .A4(
        \inq_ary[10][117] ), .Y(n1358) );
  AO22X1_RVT U1504 ( .A1(n1537), .A2(\inq_ary[15][117] ), .A3(n1738), .A4(
        \inq_ary[6][117] ), .Y(n1357) );
  AO22X1_RVT U1505 ( .A1(n1740), .A2(\inq_ary[12][117] ), .A3(n1751), .A4(
        \inq_ary[9][117] ), .Y(n1356) );
  NOR4X1_RVT U1506 ( .A1(n1359), .A2(n1358), .A3(n1357), .A4(n1356), .Y(n1365)
         );
  AO22X1_RVT U1507 ( .A1(n1729), .A2(\inq_ary[4][117] ), .A3(n1686), .A4(
        \inq_ary[0][117] ), .Y(n1363) );
  AO22X1_RVT U1508 ( .A1(n1612), .A2(\inq_ary[8][117] ), .A3(n1741), .A4(
        \inq_ary[7][117] ), .Y(n1362) );
  AO22X1_RVT U1509 ( .A1(n1742), .A2(\inq_ary[3][117] ), .A3(n1711), .A4(
        \inq_ary[13][117] ), .Y(n1361) );
  AO22X1_RVT U1510 ( .A1(n1554), .A2(\inq_ary[14][117] ), .A3(n1750), .A4(
        \inq_ary[11][117] ), .Y(n1360) );
  NOR4X1_RVT U1511 ( .A1(n1363), .A2(n1362), .A3(n1361), .A4(n1360), .Y(n1364)
         );
  NAND2X0_RVT U1512 ( .A1(n1365), .A2(n1364), .Y(n1366) );
  AO22X1_RVT U1513 ( .A1(n1477), .A2(wrdata_d1[117]), .A3(n1), .A4(n1366), .Y(
        n3442) );
  AO22X1_RVT U1514 ( .A1(n1750), .A2(\inq_ary[11][134] ), .A3(n1738), .A4(
        \inq_ary[6][134] ), .Y(n1370) );
  AO22X1_RVT U1515 ( .A1(n1554), .A2(\inq_ary[14][134] ), .A3(n1748), .A4(
        \inq_ary[10][134] ), .Y(n1369) );
  AO22X1_RVT U1516 ( .A1(n1612), .A2(\inq_ary[8][134] ), .A3(n1711), .A4(
        \inq_ary[13][134] ), .Y(n1368) );
  AO22X1_RVT U1517 ( .A1(n1742), .A2(\inq_ary[3][134] ), .A3(n1741), .A4(
        \inq_ary[7][134] ), .Y(n1367) );
  NOR4X1_RVT U1518 ( .A1(n1370), .A2(n1369), .A3(n1368), .A4(n1367), .Y(n1376)
         );
  AO22X1_RVT U1519 ( .A1(n1739), .A2(\inq_ary[2][134] ), .A3(n1751), .A4(
        \inq_ary[9][134] ), .Y(n1374) );
  AO22X1_RVT U1520 ( .A1(n1729), .A2(\inq_ary[4][134] ), .A3(n1749), .A4(
        \inq_ary[1][134] ), .Y(n1373) );
  AO22X1_RVT U1521 ( .A1(n1537), .A2(\inq_ary[15][134] ), .A3(n1740), .A4(
        \inq_ary[12][134] ), .Y(n1372) );
  AO22X1_RVT U1522 ( .A1(n1686), .A2(\inq_ary[0][134] ), .A3(n1747), .A4(
        \inq_ary[5][134] ), .Y(n1371) );
  NOR4X1_RVT U1523 ( .A1(n1374), .A2(n1373), .A3(n1372), .A4(n1371), .Y(n1375)
         );
  NAND2X0_RVT U1524 ( .A1(n1376), .A2(n1375), .Y(n1377) );
  AO22X1_RVT U1525 ( .A1(n1025), .A2(wrdata_d1[134]), .A3(n1489), .A4(n1377), 
        .Y(n3460) );
  AO22X1_RVT U1526 ( .A1(n1729), .A2(\inq_ary[4][26] ), .A3(n1749), .A4(
        \inq_ary[1][26] ), .Y(n1381) );
  AO22X1_RVT U1527 ( .A1(n1739), .A2(\inq_ary[2][26] ), .A3(n1747), .A4(
        \inq_ary[5][26] ), .Y(n1380) );
  AO22X1_RVT U1528 ( .A1(n1612), .A2(\inq_ary[8][26] ), .A3(n1751), .A4(
        \inq_ary[9][26] ), .Y(n1379) );
  AO22X1_RVT U1529 ( .A1(n1686), .A2(\inq_ary[0][26] ), .A3(n1748), .A4(
        \inq_ary[10][26] ), .Y(n1378) );
  NOR4X1_RVT U1530 ( .A1(n1381), .A2(n1380), .A3(n1379), .A4(n1378), .Y(n1387)
         );
  AO22X1_RVT U1531 ( .A1(n1750), .A2(\inq_ary[11][26] ), .A3(n1711), .A4(
        \inq_ary[13][26] ), .Y(n1385) );
  AO22X1_RVT U1532 ( .A1(n1742), .A2(\inq_ary[3][26] ), .A3(n1740), .A4(
        \inq_ary[12][26] ), .Y(n1384) );
  AO22X1_RVT U1533 ( .A1(n1537), .A2(\inq_ary[15][26] ), .A3(n1738), .A4(
        \inq_ary[6][26] ), .Y(n1383) );
  AO22X1_RVT U1534 ( .A1(n1554), .A2(\inq_ary[14][26] ), .A3(n1741), .A4(
        \inq_ary[7][26] ), .Y(n1382) );
  NOR4X1_RVT U1535 ( .A1(n1385), .A2(n1384), .A3(n1383), .A4(n1382), .Y(n1386)
         );
  NAND2X0_RVT U1536 ( .A1(n1387), .A2(n1386), .Y(n1388) );
  AO22X1_RVT U1537 ( .A1(n3), .A2(wrdata_d1[26]), .A3(n2), .A4(n1388), .Y(
        n3364) );
  AO22X1_RVT U1538 ( .A1(n1740), .A2(\inq_ary[12][119] ), .A3(n1741), .A4(
        \inq_ary[7][119] ), .Y(n1392) );
  AO22X1_RVT U1539 ( .A1(n1537), .A2(\inq_ary[15][119] ), .A3(n1612), .A4(
        \inq_ary[8][119] ), .Y(n1391) );
  AO22X1_RVT U1540 ( .A1(n1739), .A2(\inq_ary[2][119] ), .A3(n1711), .A4(
        \inq_ary[13][119] ), .Y(n1390) );
  AO22X1_RVT U1541 ( .A1(n1729), .A2(\inq_ary[4][119] ), .A3(n1750), .A4(
        \inq_ary[11][119] ), .Y(n1389) );
  NOR4X1_RVT U1542 ( .A1(n1392), .A2(n1391), .A3(n1390), .A4(n1389), .Y(n1398)
         );
  AO22X1_RVT U1543 ( .A1(n1749), .A2(\inq_ary[1][119] ), .A3(n1747), .A4(
        \inq_ary[5][119] ), .Y(n1396) );
  AO22X1_RVT U1544 ( .A1(n1742), .A2(\inq_ary[3][119] ), .A3(n1686), .A4(
        \inq_ary[0][119] ), .Y(n1395) );
  AO22X1_RVT U1545 ( .A1(n1738), .A2(\inq_ary[6][119] ), .A3(n1748), .A4(
        \inq_ary[10][119] ), .Y(n1394) );
  AO22X1_RVT U1546 ( .A1(n1554), .A2(\inq_ary[14][119] ), .A3(n1751), .A4(
        \inq_ary[9][119] ), .Y(n1393) );
  NOR4X1_RVT U1547 ( .A1(n1396), .A2(n1395), .A3(n1394), .A4(n1393), .Y(n1397)
         );
  NAND2X0_RVT U1548 ( .A1(n1398), .A2(n1397), .Y(n1399) );
  AO22X1_RVT U1549 ( .A1(n1684), .A2(wrdata_d1[119]), .A3(n1), .A4(n1399), .Y(
        n3446) );
  AO22X1_RVT U1550 ( .A1(n1747), .A2(\inq_ary[5][31] ), .A3(n1711), .A4(
        \inq_ary[13][31] ), .Y(n1403) );
  AO22X1_RVT U1551 ( .A1(n1729), .A2(\inq_ary[4][31] ), .A3(n1738), .A4(
        \inq_ary[6][31] ), .Y(n1402) );
  AO22X1_RVT U1552 ( .A1(n1612), .A2(\inq_ary[8][31] ), .A3(n1750), .A4(
        \inq_ary[11][31] ), .Y(n1401) );
  AO22X1_RVT U1553 ( .A1(n1537), .A2(\inq_ary[15][31] ), .A3(n1741), .A4(
        \inq_ary[7][31] ), .Y(n1400) );
  NOR4X1_RVT U1554 ( .A1(n1403), .A2(n1402), .A3(n1401), .A4(n1400), .Y(n1409)
         );
  AO22X1_RVT U1555 ( .A1(n1686), .A2(\inq_ary[0][31] ), .A3(n1748), .A4(
        \inq_ary[10][31] ), .Y(n1407) );
  AO22X1_RVT U1556 ( .A1(n1554), .A2(\inq_ary[14][31] ), .A3(n1751), .A4(
        \inq_ary[9][31] ), .Y(n1406) );
  AO22X1_RVT U1557 ( .A1(n1742), .A2(\inq_ary[3][31] ), .A3(n1749), .A4(
        \inq_ary[1][31] ), .Y(n1405) );
  AO22X1_RVT U1558 ( .A1(n1739), .A2(\inq_ary[2][31] ), .A3(n1740), .A4(
        \inq_ary[12][31] ), .Y(n1404) );
  NOR4X1_RVT U1559 ( .A1(n1407), .A2(n1406), .A3(n1405), .A4(n1404), .Y(n1408)
         );
  NAND2X0_RVT U1560 ( .A1(n1409), .A2(n1408), .Y(n1410) );
  AO22X1_RVT U1561 ( .A1(n1723), .A2(wrdata_d1[31]), .A3(n2), .A4(n1410), .Y(
        n3365) );
  AO22X1_RVT U1562 ( .A1(n1739), .A2(\inq_ary[2][130] ), .A3(n1741), .A4(
        \inq_ary[7][130] ), .Y(n1414) );
  AO22X1_RVT U1563 ( .A1(n1537), .A2(\inq_ary[15][130] ), .A3(n1612), .A4(
        \inq_ary[8][130] ), .Y(n1413) );
  AO22X1_RVT U1564 ( .A1(n1554), .A2(\inq_ary[14][130] ), .A3(n1749), .A4(
        \inq_ary[1][130] ), .Y(n1412) );
  AO22X1_RVT U1565 ( .A1(n1750), .A2(\inq_ary[11][130] ), .A3(n1711), .A4(
        \inq_ary[13][130] ), .Y(n1411) );
  NOR4X1_RVT U1566 ( .A1(n1414), .A2(n1413), .A3(n1412), .A4(n1411), .Y(n1420)
         );
  AO22X1_RVT U1567 ( .A1(n1748), .A2(\inq_ary[10][130] ), .A3(n1751), .A4(
        \inq_ary[9][130] ), .Y(n1418) );
  AO22X1_RVT U1568 ( .A1(n1686), .A2(\inq_ary[0][130] ), .A3(n1740), .A4(
        \inq_ary[12][130] ), .Y(n1417) );
  AO22X1_RVT U1569 ( .A1(n1742), .A2(\inq_ary[3][130] ), .A3(n1729), .A4(
        \inq_ary[4][130] ), .Y(n1416) );
  AO22X1_RVT U1570 ( .A1(n1747), .A2(\inq_ary[5][130] ), .A3(n1738), .A4(
        \inq_ary[6][130] ), .Y(n1415) );
  NOR4X1_RVT U1571 ( .A1(n1418), .A2(n1417), .A3(n1416), .A4(n1415), .Y(n1419)
         );
  NAND2X0_RVT U1572 ( .A1(n1420), .A2(n1419), .Y(n1421) );
  AO22X1_RVT U1573 ( .A1(n1477), .A2(wrdata_d1[130]), .A3(n1489), .A4(n1421), 
        .Y(n3461) );
  AO22X1_RVT U1574 ( .A1(\inq_ary[5][5] ), .A2(n1747), .A3(\inq_ary[11][5] ), 
        .A4(n1750), .Y(n1425) );
  AO22X1_RVT U1575 ( .A1(\inq_ary[1][5] ), .A2(n1749), .A3(\inq_ary[7][5] ), 
        .A4(n1741), .Y(n1424) );
  AO22X1_RVT U1576 ( .A1(\inq_ary[10][5] ), .A2(n1748), .A3(\inq_ary[9][5] ), 
        .A4(n1751), .Y(n1423) );
  AO22X1_RVT U1577 ( .A1(\inq_ary[6][5] ), .A2(n1738), .A3(\inq_ary[13][5] ), 
        .A4(n1711), .Y(n1422) );
  NOR4X1_RVT U1578 ( .A1(n1425), .A2(n1424), .A3(n1423), .A4(n1422), .Y(n1431)
         );
  AO22X1_RVT U1579 ( .A1(\inq_ary[3][5] ), .A2(n1742), .A3(\inq_ary[4][5] ), 
        .A4(n1729), .Y(n1429) );
  AO22X1_RVT U1580 ( .A1(\inq_ary[2][5] ), .A2(n1739), .A3(\inq_ary[14][5] ), 
        .A4(n1554), .Y(n1428) );
  AO22X1_RVT U1581 ( .A1(\inq_ary[8][5] ), .A2(n1612), .A3(\inq_ary[12][5] ), 
        .A4(n1740), .Y(n1427) );
  AO22X1_RVT U1582 ( .A1(\inq_ary[0][5] ), .A2(n1686), .A3(\inq_ary[15][5] ), 
        .A4(n1537), .Y(n1426) );
  NOR4X1_RVT U1583 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .Y(n1430)
         );
  NAND2X0_RVT U1584 ( .A1(n1431), .A2(n1430), .Y(n1432) );
  AO22X1_RVT U1585 ( .A1(n3), .A2(wrdata_d1[5]), .A3(n1), .A4(n1432), .Y(n3340) );
  AO22X1_RVT U1586 ( .A1(n1750), .A2(\inq_ary[11][27] ), .A3(n1751), .A4(
        \inq_ary[9][27] ), .Y(n1436) );
  AO22X1_RVT U1587 ( .A1(n1537), .A2(\inq_ary[15][27] ), .A3(n1711), .A4(
        \inq_ary[13][27] ), .Y(n1435) );
  AO22X1_RVT U1588 ( .A1(n1729), .A2(\inq_ary[4][27] ), .A3(n1741), .A4(
        \inq_ary[7][27] ), .Y(n1434) );
  AO22X1_RVT U1589 ( .A1(n1686), .A2(\inq_ary[0][27] ), .A3(n1747), .A4(
        \inq_ary[5][27] ), .Y(n1433) );
  NOR4X1_RVT U1590 ( .A1(n1436), .A2(n1435), .A3(n1434), .A4(n1433), .Y(n1442)
         );
  AO22X1_RVT U1591 ( .A1(n1742), .A2(\inq_ary[3][27] ), .A3(n1740), .A4(
        \inq_ary[12][27] ), .Y(n1440) );
  AO22X1_RVT U1592 ( .A1(n1554), .A2(\inq_ary[14][27] ), .A3(n1738), .A4(
        \inq_ary[6][27] ), .Y(n1439) );
  AO22X1_RVT U1593 ( .A1(n1612), .A2(\inq_ary[8][27] ), .A3(n1748), .A4(
        \inq_ary[10][27] ), .Y(n1438) );
  AO22X1_RVT U1594 ( .A1(n1739), .A2(\inq_ary[2][27] ), .A3(n1749), .A4(
        \inq_ary[1][27] ), .Y(n1437) );
  NOR4X1_RVT U1595 ( .A1(n1440), .A2(n1439), .A3(n1438), .A4(n1437), .Y(n1441)
         );
  NAND2X0_RVT U1596 ( .A1(n1442), .A2(n1441), .Y(n1443) );
  AO22X1_RVT U1597 ( .A1(n1760), .A2(wrdata_d1[27]), .A3(n2), .A4(n1443), .Y(
        n3366) );
  AO22X1_RVT U1598 ( .A1(n1739), .A2(\inq_ary[2][124] ), .A3(n1742), .A4(
        \inq_ary[3][124] ), .Y(n1447) );
  AO22X1_RVT U1599 ( .A1(n1686), .A2(\inq_ary[0][124] ), .A3(n1749), .A4(
        \inq_ary[1][124] ), .Y(n1446) );
  AO22X1_RVT U1600 ( .A1(n1537), .A2(\inq_ary[15][124] ), .A3(n1612), .A4(
        \inq_ary[8][124] ), .Y(n1445) );
  AO22X1_RVT U1601 ( .A1(n1747), .A2(\inq_ary[5][124] ), .A3(n1750), .A4(
        \inq_ary[11][124] ), .Y(n1444) );
  NOR4X1_RVT U1602 ( .A1(n1447), .A2(n1446), .A3(n1445), .A4(n1444), .Y(n1453)
         );
  AO22X1_RVT U1603 ( .A1(n1738), .A2(\inq_ary[6][124] ), .A3(n1751), .A4(
        \inq_ary[9][124] ), .Y(n1451) );
  AO22X1_RVT U1604 ( .A1(n1740), .A2(\inq_ary[12][124] ), .A3(n1741), .A4(
        \inq_ary[7][124] ), .Y(n1450) );
  AO22X1_RVT U1605 ( .A1(n1554), .A2(\inq_ary[14][124] ), .A3(n1711), .A4(
        \inq_ary[13][124] ), .Y(n1449) );
  AO22X1_RVT U1606 ( .A1(n1729), .A2(\inq_ary[4][124] ), .A3(n1748), .A4(
        \inq_ary[10][124] ), .Y(n1448) );
  NOR4X1_RVT U1607 ( .A1(n1451), .A2(n1450), .A3(n1449), .A4(n1448), .Y(n1452)
         );
  NAND2X0_RVT U1608 ( .A1(n1453), .A2(n1452), .Y(n1454) );
  AO22X1_RVT U1609 ( .A1(n1723), .A2(wrdata_d1[124]), .A3(n1), .A4(n1454), .Y(
        n3448) );
  AO22X1_RVT U1610 ( .A1(n1740), .A2(\inq_ary[12][122] ), .A3(n1711), .A4(
        \inq_ary[13][122] ), .Y(n1458) );
  AO22X1_RVT U1611 ( .A1(n1742), .A2(\inq_ary[3][122] ), .A3(n1537), .A4(
        \inq_ary[15][122] ), .Y(n1457) );
  AO22X1_RVT U1612 ( .A1(n1729), .A2(\inq_ary[4][122] ), .A3(n1738), .A4(
        \inq_ary[6][122] ), .Y(n1456) );
  AO22X1_RVT U1613 ( .A1(n1741), .A2(\inq_ary[7][122] ), .A3(n1751), .A4(
        \inq_ary[9][122] ), .Y(n1455) );
  NOR4X1_RVT U1614 ( .A1(n1458), .A2(n1457), .A3(n1456), .A4(n1455), .Y(n1464)
         );
  AO22X1_RVT U1615 ( .A1(n1739), .A2(\inq_ary[2][122] ), .A3(n1612), .A4(
        \inq_ary[8][122] ), .Y(n1462) );
  AO22X1_RVT U1616 ( .A1(n1554), .A2(\inq_ary[14][122] ), .A3(n1748), .A4(
        \inq_ary[10][122] ), .Y(n1461) );
  AO22X1_RVT U1617 ( .A1(n1686), .A2(\inq_ary[0][122] ), .A3(n1750), .A4(
        \inq_ary[11][122] ), .Y(n1460) );
  AO22X1_RVT U1618 ( .A1(n1749), .A2(\inq_ary[1][122] ), .A3(n1747), .A4(
        \inq_ary[5][122] ), .Y(n1459) );
  NOR4X1_RVT U1619 ( .A1(n1462), .A2(n1461), .A3(n1460), .A4(n1459), .Y(n1463)
         );
  NAND2X0_RVT U1620 ( .A1(n1464), .A2(n1463), .Y(n1465) );
  AO22X1_RVT U1621 ( .A1(n1760), .A2(wrdata_d1[122]), .A3(n1489), .A4(n1465), 
        .Y(n3453) );
  AO22X1_RVT U1622 ( .A1(n1554), .A2(\inq_ary[14][118] ), .A3(n1711), .A4(
        \inq_ary[13][118] ), .Y(n1469) );
  AO22X1_RVT U1623 ( .A1(n1747), .A2(\inq_ary[5][118] ), .A3(n1751), .A4(
        \inq_ary[9][118] ), .Y(n1468) );
  AO22X1_RVT U1624 ( .A1(n1742), .A2(\inq_ary[3][118] ), .A3(n1729), .A4(
        \inq_ary[4][118] ), .Y(n1467) );
  AO22X1_RVT U1625 ( .A1(n1686), .A2(\inq_ary[0][118] ), .A3(n1740), .A4(
        \inq_ary[12][118] ), .Y(n1466) );
  NOR4X1_RVT U1626 ( .A1(n1469), .A2(n1468), .A3(n1467), .A4(n1466), .Y(n1475)
         );
  AO22X1_RVT U1627 ( .A1(n1612), .A2(\inq_ary[8][118] ), .A3(n1750), .A4(
        \inq_ary[11][118] ), .Y(n1473) );
  AO22X1_RVT U1628 ( .A1(n1738), .A2(\inq_ary[6][118] ), .A3(n1748), .A4(
        \inq_ary[10][118] ), .Y(n1472) );
  AO22X1_RVT U1629 ( .A1(n1739), .A2(\inq_ary[2][118] ), .A3(n1741), .A4(
        \inq_ary[7][118] ), .Y(n1471) );
  AO22X1_RVT U1630 ( .A1(n1537), .A2(\inq_ary[15][118] ), .A3(n1749), .A4(
        \inq_ary[1][118] ), .Y(n1470) );
  NOR4X1_RVT U1631 ( .A1(n1473), .A2(n1472), .A3(n1471), .A4(n1470), .Y(n1474)
         );
  NAND2X0_RVT U1632 ( .A1(n1475), .A2(n1474), .Y(n1476) );
  AO22X1_RVT U1633 ( .A1(n1477), .A2(wrdata_d1[118]), .A3(n1), .A4(n1476), .Y(
        n3444) );
  AO22X1_RVT U1634 ( .A1(n1686), .A2(\inq_ary[0][131] ), .A3(n1750), .A4(
        \inq_ary[11][131] ), .Y(n1481) );
  AO22X1_RVT U1635 ( .A1(n1741), .A2(\inq_ary[7][131] ), .A3(n1748), .A4(
        \inq_ary[10][131] ), .Y(n1480) );
  AO22X1_RVT U1636 ( .A1(n1729), .A2(\inq_ary[4][131] ), .A3(n1612), .A4(
        \inq_ary[8][131] ), .Y(n1479) );
  AO22X1_RVT U1637 ( .A1(n1742), .A2(\inq_ary[3][131] ), .A3(n1747), .A4(
        \inq_ary[5][131] ), .Y(n1478) );
  NOR4X1_RVT U1638 ( .A1(n1481), .A2(n1480), .A3(n1479), .A4(n1478), .Y(n1487)
         );
  AO22X1_RVT U1639 ( .A1(n1537), .A2(\inq_ary[15][131] ), .A3(n1751), .A4(
        \inq_ary[9][131] ), .Y(n1485) );
  AO22X1_RVT U1640 ( .A1(n1749), .A2(\inq_ary[1][131] ), .A3(n1711), .A4(
        \inq_ary[13][131] ), .Y(n1484) );
  AO22X1_RVT U1641 ( .A1(n1740), .A2(\inq_ary[12][131] ), .A3(n1738), .A4(
        \inq_ary[6][131] ), .Y(n1483) );
  AO22X1_RVT U1642 ( .A1(n1739), .A2(\inq_ary[2][131] ), .A3(n1554), .A4(
        \inq_ary[14][131] ), .Y(n1482) );
  NOR4X1_RVT U1643 ( .A1(n1485), .A2(n1484), .A3(n1483), .A4(n1482), .Y(n1486)
         );
  NAND2X0_RVT U1644 ( .A1(n1487), .A2(n1486), .Y(n1488) );
  AO22X1_RVT U1645 ( .A1(n1684), .A2(wrdata_d1[131]), .A3(n1489), .A4(n1488), 
        .Y(n3463) );
  AO22X1_RVT U1646 ( .A1(n1739), .A2(\inq_ary[2][6] ), .A3(n1751), .A4(
        \inq_ary[9][6] ), .Y(n1493) );
  AO22X1_RVT U1647 ( .A1(n1612), .A2(\inq_ary[8][6] ), .A3(n1738), .A4(
        \inq_ary[6][6] ), .Y(n1492) );
  AO22X1_RVT U1648 ( .A1(n1554), .A2(\inq_ary[14][6] ), .A3(n1748), .A4(
        \inq_ary[10][6] ), .Y(n1491) );
  AO22X1_RVT U1649 ( .A1(n1686), .A2(\inq_ary[0][6] ), .A3(n1747), .A4(
        \inq_ary[5][6] ), .Y(n1490) );
  NOR4X1_RVT U1650 ( .A1(n1493), .A2(n1492), .A3(n1491), .A4(n1490), .Y(n1499)
         );
  AO22X1_RVT U1651 ( .A1(n1729), .A2(\inq_ary[4][6] ), .A3(n1537), .A4(
        \inq_ary[15][6] ), .Y(n1497) );
  AO22X1_RVT U1652 ( .A1(n1740), .A2(\inq_ary[12][6] ), .A3(n1741), .A4(
        \inq_ary[7][6] ), .Y(n1496) );
  AO22X1_RVT U1653 ( .A1(n1749), .A2(\inq_ary[1][6] ), .A3(n1750), .A4(
        \inq_ary[11][6] ), .Y(n1495) );
  AO22X1_RVT U1654 ( .A1(n1742), .A2(\inq_ary[3][6] ), .A3(n1711), .A4(
        \inq_ary[13][6] ), .Y(n1494) );
  NOR4X1_RVT U1655 ( .A1(n1497), .A2(n1496), .A3(n1495), .A4(n1494), .Y(n1498)
         );
  NAND2X0_RVT U1656 ( .A1(n1499), .A2(n1498), .Y(n1500) );
  AO22X1_RVT U1657 ( .A1(n1684), .A2(wrdata_d1[6]), .A3(n1489), .A4(n1500), 
        .Y(n3341) );
  AO22X1_RVT U1658 ( .A1(n1554), .A2(\inq_ary[14][30] ), .A3(n1729), .A4(
        \inq_ary[4][30] ), .Y(n1504) );
  AO22X1_RVT U1659 ( .A1(n1612), .A2(\inq_ary[8][30] ), .A3(n1747), .A4(
        \inq_ary[5][30] ), .Y(n1503) );
  AO22X1_RVT U1660 ( .A1(n1739), .A2(\inq_ary[2][30] ), .A3(n1537), .A4(
        \inq_ary[15][30] ), .Y(n1502) );
  AO22X1_RVT U1661 ( .A1(n1686), .A2(\inq_ary[0][30] ), .A3(n1738), .A4(
        \inq_ary[6][30] ), .Y(n1501) );
  NOR4X1_RVT U1662 ( .A1(n1504), .A2(n1503), .A3(n1502), .A4(n1501), .Y(n1510)
         );
  AO22X1_RVT U1663 ( .A1(n1750), .A2(\inq_ary[11][30] ), .A3(n1751), .A4(
        \inq_ary[9][30] ), .Y(n1508) );
  AO22X1_RVT U1664 ( .A1(n1740), .A2(\inq_ary[12][30] ), .A3(n1748), .A4(
        \inq_ary[10][30] ), .Y(n1507) );
  AO22X1_RVT U1665 ( .A1(n1749), .A2(\inq_ary[1][30] ), .A3(n1711), .A4(
        \inq_ary[13][30] ), .Y(n1506) );
  AO22X1_RVT U1666 ( .A1(n1742), .A2(\inq_ary[3][30] ), .A3(n1741), .A4(
        \inq_ary[7][30] ), .Y(n1505) );
  NOR4X1_RVT U1667 ( .A1(n1508), .A2(n1507), .A3(n1506), .A4(n1505), .Y(n1509)
         );
  NAND2X0_RVT U1668 ( .A1(n1510), .A2(n1509), .Y(n1511) );
  AO22X1_RVT U1669 ( .A1(n1598), .A2(wrdata_d1[30]), .A3(n946), .A4(n1511), 
        .Y(n3363) );
  AND2X1_RVT U1670 ( .A1(n1760), .A2(reset_l), .Y(n1512) );
  AND2X1_RVT U1671 ( .A1(n1747), .A2(n1512), .Y(n3486) );
  AND2X1_RVT U1672 ( .A1(n1738), .A2(n1512), .Y(n3485) );
  AND2X1_RVT U1673 ( .A1(n1741), .A2(n1512), .Y(n3484) );
  AND2X1_RVT U1674 ( .A1(n1612), .A2(n1512), .Y(n3483) );
  AND2X1_RVT U1675 ( .A1(n1751), .A2(n1512), .Y(n3482) );
  AND2X1_RVT U1676 ( .A1(n1748), .A2(n1512), .Y(n3481) );
  AND2X1_RVT U1677 ( .A1(n1750), .A2(n1512), .Y(n3480) );
  AND2X1_RVT U1678 ( .A1(n1740), .A2(n1512), .Y(n3479) );
  AND2X1_RVT U1679 ( .A1(n1711), .A2(n1512), .Y(n3478) );
  AND2X1_RVT U1680 ( .A1(n1554), .A2(n1512), .Y(n3477) );
  AND2X1_RVT U1681 ( .A1(n1537), .A2(n1512), .Y(n3476) );
  AND2X1_RVT U1682 ( .A1(n1686), .A2(n1512), .Y(n3491) );
  AND2X1_RVT U1683 ( .A1(n1749), .A2(n1512), .Y(n3490) );
  AND2X1_RVT U1684 ( .A1(n1739), .A2(n1512), .Y(n3489) );
  AND2X1_RVT U1685 ( .A1(n1742), .A2(n1512), .Y(n3488) );
  AND2X1_RVT U1686 ( .A1(n1729), .A2(n1512), .Y(n3487) );
  INVX1_RVT U1687 ( .A(sehold), .Y(n3574) );
  AO22X1_RVT U1688 ( .A1(n1612), .A2(\inq_ary[8][59] ), .A3(n1740), .A4(
        \inq_ary[12][59] ), .Y(n1516) );
  AO22X1_RVT U1689 ( .A1(n1739), .A2(\inq_ary[2][59] ), .A3(n1537), .A4(
        \inq_ary[15][59] ), .Y(n1515) );
  AO22X1_RVT U1690 ( .A1(n1686), .A2(\inq_ary[0][59] ), .A3(n1741), .A4(
        \inq_ary[7][59] ), .Y(n1514) );
  AO22X1_RVT U1691 ( .A1(n1711), .A2(\inq_ary[13][59] ), .A3(n1751), .A4(
        \inq_ary[9][59] ), .Y(n1513) );
  NOR4X1_RVT U1692 ( .A1(n1516), .A2(n1515), .A3(n1514), .A4(n1513), .Y(n1522)
         );
  AO22X1_RVT U1693 ( .A1(n1729), .A2(\inq_ary[4][59] ), .A3(n1738), .A4(
        \inq_ary[6][59] ), .Y(n1520) );
  AO22X1_RVT U1694 ( .A1(n1554), .A2(\inq_ary[14][59] ), .A3(n1749), .A4(
        \inq_ary[1][59] ), .Y(n1519) );
  AO22X1_RVT U1695 ( .A1(n1750), .A2(\inq_ary[11][59] ), .A3(n1748), .A4(
        \inq_ary[10][59] ), .Y(n1518) );
  AO22X1_RVT U1696 ( .A1(n1742), .A2(\inq_ary[3][59] ), .A3(n1747), .A4(
        \inq_ary[5][59] ), .Y(n1517) );
  NOR4X1_RVT U1697 ( .A1(n1520), .A2(n1519), .A3(n1518), .A4(n1517), .Y(n1521)
         );
  NAND2X0_RVT U1698 ( .A1(n1522), .A2(n1521), .Y(n1523) );
  AO22X1_RVT U1699 ( .A1(n3), .A2(wrdata_d1[59]), .A3(n969), .A4(n1523), .Y(
        n1524) );
  AO22X1_RVT U1700 ( .A1(n1740), .A2(\inq_ary[12][62] ), .A3(n1751), .A4(
        \inq_ary[9][62] ), .Y(n1528) );
  AO22X1_RVT U1701 ( .A1(n1749), .A2(\inq_ary[1][62] ), .A3(n1711), .A4(
        \inq_ary[13][62] ), .Y(n1527) );
  AO22X1_RVT U1702 ( .A1(n1612), .A2(\inq_ary[8][62] ), .A3(n1738), .A4(
        \inq_ary[6][62] ), .Y(n1526) );
  AO22X1_RVT U1703 ( .A1(n1537), .A2(\inq_ary[15][62] ), .A3(n1750), .A4(
        \inq_ary[11][62] ), .Y(n1525) );
  NOR4X1_RVT U1704 ( .A1(n1528), .A2(n1527), .A3(n1526), .A4(n1525), .Y(n1534)
         );
  AO22X1_RVT U1705 ( .A1(n1739), .A2(\inq_ary[2][62] ), .A3(n1686), .A4(
        \inq_ary[0][62] ), .Y(n1532) );
  AO22X1_RVT U1706 ( .A1(n1554), .A2(\inq_ary[14][62] ), .A3(n1742), .A4(
        \inq_ary[3][62] ), .Y(n1531) );
  AO22X1_RVT U1707 ( .A1(n1729), .A2(\inq_ary[4][62] ), .A3(n1741), .A4(
        \inq_ary[7][62] ), .Y(n1530) );
  AO22X1_RVT U1708 ( .A1(n1747), .A2(\inq_ary[5][62] ), .A3(n1748), .A4(
        \inq_ary[10][62] ), .Y(n1529) );
  NOR4X1_RVT U1709 ( .A1(n1532), .A2(n1531), .A3(n1530), .A4(n1529), .Y(n1533)
         );
  NAND2X0_RVT U1710 ( .A1(n1534), .A2(n1533), .Y(n1535) );
  AO22X1_RVT U1711 ( .A1(n3), .A2(wrdata_d1[62]), .A3(n2), .A4(n1535), .Y(
        n1536) );
  AO22X1_RVT U1712 ( .A1(n1739), .A2(\inq_ary[2][63] ), .A3(n1749), .A4(
        \inq_ary[1][63] ), .Y(n1541) );
  AO22X1_RVT U1713 ( .A1(n1686), .A2(\inq_ary[0][63] ), .A3(n1738), .A4(
        \inq_ary[6][63] ), .Y(n1540) );
  AO22X1_RVT U1714 ( .A1(n1537), .A2(\inq_ary[15][63] ), .A3(n1612), .A4(
        \inq_ary[8][63] ), .Y(n1539) );
  AO22X1_RVT U1715 ( .A1(n1750), .A2(\inq_ary[11][63] ), .A3(n1748), .A4(
        \inq_ary[10][63] ), .Y(n1538) );
  NOR4X1_RVT U1716 ( .A1(n1541), .A2(n1540), .A3(n1539), .A4(n1538), .Y(n1547)
         );
  AO22X1_RVT U1717 ( .A1(n1729), .A2(\inq_ary[4][63] ), .A3(n1711), .A4(
        \inq_ary[13][63] ), .Y(n1545) );
  AO22X1_RVT U1718 ( .A1(n1740), .A2(\inq_ary[12][63] ), .A3(n1741), .A4(
        \inq_ary[7][63] ), .Y(n1544) );
  AO22X1_RVT U1719 ( .A1(n1747), .A2(\inq_ary[5][63] ), .A3(n1751), .A4(
        \inq_ary[9][63] ), .Y(n1543) );
  AO22X1_RVT U1720 ( .A1(n1554), .A2(\inq_ary[14][63] ), .A3(n1742), .A4(
        \inq_ary[3][63] ), .Y(n1542) );
  NOR4X1_RVT U1721 ( .A1(n1545), .A2(n1544), .A3(n1543), .A4(n1542), .Y(n1546)
         );
  NAND2X0_RVT U1722 ( .A1(n1547), .A2(n1546), .Y(n1548) );
  AO22X1_RVT U1723 ( .A1(n3), .A2(wrdata_d1[63]), .A3(n1489), .A4(n1548), .Y(
        n1549) );
  AO22X1_RVT U1724 ( .A1(n1739), .A2(\inq_ary[2][58] ), .A3(n1749), .A4(
        \inq_ary[1][58] ), .Y(n1553) );
  AO22X1_RVT U1725 ( .A1(n1740), .A2(\inq_ary[12][58] ), .A3(n1738), .A4(
        \inq_ary[6][58] ), .Y(n1552) );
  AO22X1_RVT U1726 ( .A1(n1729), .A2(\inq_ary[4][58] ), .A3(n1750), .A4(
        \inq_ary[11][58] ), .Y(n1551) );
  AO22X1_RVT U1727 ( .A1(n1686), .A2(\inq_ary[0][58] ), .A3(n1741), .A4(
        \inq_ary[7][58] ), .Y(n1550) );
  NOR4X1_RVT U1728 ( .A1(n1553), .A2(n1552), .A3(n1551), .A4(n1550), .Y(n1560)
         );
  AO22X1_RVT U1729 ( .A1(n1742), .A2(\inq_ary[3][58] ), .A3(n1748), .A4(
        \inq_ary[10][58] ), .Y(n1558) );
  AO22X1_RVT U1730 ( .A1(n1554), .A2(\inq_ary[14][58] ), .A3(n1747), .A4(
        \inq_ary[5][58] ), .Y(n1557) );
  AO22X1_RVT U1731 ( .A1(n1537), .A2(\inq_ary[15][58] ), .A3(n1612), .A4(
        \inq_ary[8][58] ), .Y(n1556) );
  AO22X1_RVT U1732 ( .A1(n1711), .A2(\inq_ary[13][58] ), .A3(n1751), .A4(
        \inq_ary[9][58] ), .Y(n1555) );
  NOR4X1_RVT U1733 ( .A1(n1558), .A2(n1557), .A3(n1556), .A4(n1555), .Y(n1559)
         );
  NAND2X0_RVT U1734 ( .A1(n1560), .A2(n1559), .Y(n1561) );
  AO22X1_RVT U1735 ( .A1(n3), .A2(wrdata_d1[58]), .A3(n1), .A4(n1561), .Y(
        n1562) );
  AO22X1_RVT U1736 ( .A1(n1742), .A2(\inq_ary[3][57] ), .A3(n1612), .A4(
        \inq_ary[8][57] ), .Y(n1566) );
  AO22X1_RVT U1737 ( .A1(n1750), .A2(\inq_ary[11][57] ), .A3(n1711), .A4(
        \inq_ary[13][57] ), .Y(n1565) );
  AO22X1_RVT U1738 ( .A1(n1747), .A2(\inq_ary[5][57] ), .A3(n1738), .A4(
        \inq_ary[6][57] ), .Y(n1564) );
  AO22X1_RVT U1739 ( .A1(n1554), .A2(\inq_ary[14][57] ), .A3(n1741), .A4(
        \inq_ary[7][57] ), .Y(n1563) );
  NOR4X1_RVT U1740 ( .A1(n1566), .A2(n1565), .A3(n1564), .A4(n1563), .Y(n1572)
         );
  AO22X1_RVT U1741 ( .A1(n1686), .A2(\inq_ary[0][57] ), .A3(n1537), .A4(
        \inq_ary[15][57] ), .Y(n1570) );
  AO22X1_RVT U1742 ( .A1(n1740), .A2(\inq_ary[12][57] ), .A3(n1748), .A4(
        \inq_ary[10][57] ), .Y(n1569) );
  AO22X1_RVT U1743 ( .A1(n1739), .A2(\inq_ary[2][57] ), .A3(n1751), .A4(
        \inq_ary[9][57] ), .Y(n1568) );
  AO22X1_RVT U1744 ( .A1(n1729), .A2(\inq_ary[4][57] ), .A3(n1749), .A4(
        \inq_ary[1][57] ), .Y(n1567) );
  NOR4X1_RVT U1745 ( .A1(n1570), .A2(n1569), .A3(n1568), .A4(n1567), .Y(n1571)
         );
  NAND2X0_RVT U1746 ( .A1(n1572), .A2(n1571), .Y(n1573) );
  AO22X1_RVT U1747 ( .A1(n3), .A2(wrdata_d1[57]), .A3(n1), .A4(n1573), .Y(
        n1574) );
  AO22X1_RVT U1748 ( .A1(n1740), .A2(\inq_ary[12][56] ), .A3(n1741), .A4(
        \inq_ary[7][56] ), .Y(n1578) );
  AO22X1_RVT U1749 ( .A1(n1739), .A2(\inq_ary[2][56] ), .A3(n1751), .A4(
        \inq_ary[9][56] ), .Y(n1577) );
  AO22X1_RVT U1750 ( .A1(n1686), .A2(\inq_ary[0][56] ), .A3(n1750), .A4(
        \inq_ary[11][56] ), .Y(n1576) );
  AO22X1_RVT U1751 ( .A1(n1747), .A2(\inq_ary[5][56] ), .A3(n1748), .A4(
        \inq_ary[10][56] ), .Y(n1575) );
  NOR4X1_RVT U1752 ( .A1(n1578), .A2(n1577), .A3(n1576), .A4(n1575), .Y(n1584)
         );
  AO22X1_RVT U1753 ( .A1(n1554), .A2(\inq_ary[14][56] ), .A3(n1738), .A4(
        \inq_ary[6][56] ), .Y(n1582) );
  AO22X1_RVT U1754 ( .A1(n1749), .A2(\inq_ary[1][56] ), .A3(n1711), .A4(
        \inq_ary[13][56] ), .Y(n1581) );
  AO22X1_RVT U1755 ( .A1(n1742), .A2(\inq_ary[3][56] ), .A3(n1537), .A4(
        \inq_ary[15][56] ), .Y(n1580) );
  AO22X1_RVT U1756 ( .A1(n1729), .A2(\inq_ary[4][56] ), .A3(n1612), .A4(
        \inq_ary[8][56] ), .Y(n1579) );
  NOR4X1_RVT U1757 ( .A1(n1582), .A2(n1581), .A3(n1580), .A4(n1579), .Y(n1583)
         );
  NAND2X0_RVT U1758 ( .A1(n1584), .A2(n1583), .Y(n1585) );
  AO22X1_RVT U1759 ( .A1(n1760), .A2(wrdata_d1[56]), .A3(n1759), .A4(n1585), 
        .Y(n1586) );
  AO22X1_RVT U1760 ( .A1(n1554), .A2(\inq_ary[14][52] ), .A3(n1740), .A4(
        \inq_ary[12][52] ), .Y(n1590) );
  AO22X1_RVT U1761 ( .A1(n1739), .A2(\inq_ary[2][52] ), .A3(n1686), .A4(
        \inq_ary[0][52] ), .Y(n1589) );
  AO22X1_RVT U1762 ( .A1(n1742), .A2(\inq_ary[3][52] ), .A3(n1751), .A4(
        \inq_ary[9][52] ), .Y(n1588) );
  AO22X1_RVT U1763 ( .A1(n1612), .A2(\inq_ary[8][52] ), .A3(n1749), .A4(
        \inq_ary[1][52] ), .Y(n1587) );
  NOR4X1_RVT U1764 ( .A1(n1590), .A2(n1589), .A3(n1588), .A4(n1587), .Y(n1596)
         );
  AO22X1_RVT U1765 ( .A1(n1750), .A2(\inq_ary[11][52] ), .A3(n1748), .A4(
        \inq_ary[10][52] ), .Y(n1594) );
  AO22X1_RVT U1766 ( .A1(n1537), .A2(\inq_ary[15][52] ), .A3(n1741), .A4(
        \inq_ary[7][52] ), .Y(n1593) );
  AO22X1_RVT U1767 ( .A1(n1747), .A2(\inq_ary[5][52] ), .A3(n1711), .A4(
        \inq_ary[13][52] ), .Y(n1592) );
  AO22X1_RVT U1768 ( .A1(n1729), .A2(\inq_ary[4][52] ), .A3(n1738), .A4(
        \inq_ary[6][52] ), .Y(n1591) );
  NOR4X1_RVT U1769 ( .A1(n1594), .A2(n1593), .A3(n1592), .A4(n1591), .Y(n1595)
         );
  NAND2X0_RVT U1770 ( .A1(n1596), .A2(n1595), .Y(n1597) );
  AO22X1_RVT U1771 ( .A1(n1598), .A2(wrdata_d1[52]), .A3(n969), .A4(n1597), 
        .Y(n1599) );
  AO22X1_RVT U1772 ( .A1(n1740), .A2(\inq_ary[12][154] ), .A3(n1749), .A4(
        \inq_ary[1][154] ), .Y(n1603) );
  AO22X1_RVT U1773 ( .A1(n1554), .A2(\inq_ary[14][154] ), .A3(n1686), .A4(
        \inq_ary[0][154] ), .Y(n1602) );
  AO22X1_RVT U1774 ( .A1(n1729), .A2(\inq_ary[4][154] ), .A3(n1537), .A4(
        \inq_ary[15][154] ), .Y(n1601) );
  AO22X1_RVT U1775 ( .A1(n1738), .A2(\inq_ary[6][154] ), .A3(n1751), .A4(
        \inq_ary[9][154] ), .Y(n1600) );
  NOR4X1_RVT U1776 ( .A1(n1603), .A2(n1602), .A3(n1601), .A4(n1600), .Y(n1609)
         );
  AO22X1_RVT U1777 ( .A1(n1747), .A2(\inq_ary[5][154] ), .A3(n1711), .A4(
        \inq_ary[13][154] ), .Y(n1607) );
  AO22X1_RVT U1778 ( .A1(n1750), .A2(\inq_ary[11][154] ), .A3(n1748), .A4(
        \inq_ary[10][154] ), .Y(n1606) );
  AO22X1_RVT U1779 ( .A1(n1739), .A2(\inq_ary[2][154] ), .A3(n1741), .A4(
        \inq_ary[7][154] ), .Y(n1605) );
  AO22X1_RVT U1780 ( .A1(n1742), .A2(\inq_ary[3][154] ), .A3(n1612), .A4(
        \inq_ary[8][154] ), .Y(n1604) );
  NOR4X1_RVT U1781 ( .A1(n1607), .A2(n1606), .A3(n1605), .A4(n1604), .Y(n1608)
         );
  NAND2X0_RVT U1782 ( .A1(n1609), .A2(n1608), .Y(n1610) );
  AO22X1_RVT U1783 ( .A1(n1760), .A2(wrdata_d1[154]), .A3(n1759), .A4(n1610), 
        .Y(n1611) );
  AO22X1_RVT U1784 ( .A1(n1750), .A2(\inq_ary[11][155] ), .A3(n1711), .A4(
        \inq_ary[13][155] ), .Y(n1616) );
  AO22X1_RVT U1785 ( .A1(n1739), .A2(\inq_ary[2][155] ), .A3(n1554), .A4(
        \inq_ary[14][155] ), .Y(n1615) );
  AO22X1_RVT U1786 ( .A1(n1729), .A2(\inq_ary[4][155] ), .A3(n1738), .A4(
        \inq_ary[6][155] ), .Y(n1614) );
  AO22X1_RVT U1787 ( .A1(n1537), .A2(\inq_ary[15][155] ), .A3(n1612), .A4(
        \inq_ary[8][155] ), .Y(n1613) );
  NOR4X1_RVT U1788 ( .A1(n1616), .A2(n1615), .A3(n1614), .A4(n1613), .Y(n1622)
         );
  AO22X1_RVT U1789 ( .A1(n1742), .A2(\inq_ary[3][155] ), .A3(n1747), .A4(
        \inq_ary[5][155] ), .Y(n1620) );
  AO22X1_RVT U1790 ( .A1(n1749), .A2(\inq_ary[1][155] ), .A3(n1751), .A4(
        \inq_ary[9][155] ), .Y(n1619) );
  AO22X1_RVT U1791 ( .A1(n1741), .A2(\inq_ary[7][155] ), .A3(n1748), .A4(
        \inq_ary[10][155] ), .Y(n1618) );
  AO22X1_RVT U1792 ( .A1(n1686), .A2(\inq_ary[0][155] ), .A3(n1740), .A4(
        \inq_ary[12][155] ), .Y(n1617) );
  NOR4X1_RVT U1793 ( .A1(n1620), .A2(n1619), .A3(n1618), .A4(n1617), .Y(n1621)
         );
  NAND2X0_RVT U1794 ( .A1(n1622), .A2(n1621), .Y(n1623) );
  AO22X1_RVT U1795 ( .A1(n1760), .A2(wrdata_d1[155]), .A3(n1759), .A4(n1623), 
        .Y(n1624) );
  AO22X1_RVT U1796 ( .A1(n1748), .A2(\inq_ary[10][156] ), .A3(n1751), .A4(
        \inq_ary[9][156] ), .Y(n1628) );
  AO22X1_RVT U1797 ( .A1(n1740), .A2(\inq_ary[12][156] ), .A3(n1738), .A4(
        \inq_ary[6][156] ), .Y(n1627) );
  AO22X1_RVT U1798 ( .A1(n1686), .A2(\inq_ary[0][156] ), .A3(n1612), .A4(
        \inq_ary[8][156] ), .Y(n1626) );
  AO22X1_RVT U1799 ( .A1(n1749), .A2(\inq_ary[1][156] ), .A3(n1750), .A4(
        \inq_ary[11][156] ), .Y(n1625) );
  NOR4X1_RVT U1800 ( .A1(n1628), .A2(n1627), .A3(n1626), .A4(n1625), .Y(n1634)
         );
  AO22X1_RVT U1801 ( .A1(n1537), .A2(\inq_ary[15][156] ), .A3(n1747), .A4(
        \inq_ary[5][156] ), .Y(n1632) );
  AO22X1_RVT U1802 ( .A1(n1554), .A2(\inq_ary[14][156] ), .A3(n1742), .A4(
        \inq_ary[3][156] ), .Y(n1631) );
  AO22X1_RVT U1803 ( .A1(n1729), .A2(\inq_ary[4][156] ), .A3(n1741), .A4(
        \inq_ary[7][156] ), .Y(n1630) );
  AO22X1_RVT U1804 ( .A1(n1739), .A2(\inq_ary[2][156] ), .A3(n1711), .A4(
        \inq_ary[13][156] ), .Y(n1629) );
  NOR4X1_RVT U1805 ( .A1(n1632), .A2(n1631), .A3(n1630), .A4(n1629), .Y(n1633)
         );
  NAND2X0_RVT U1806 ( .A1(n1634), .A2(n1633), .Y(n1635) );
  AO22X1_RVT U1807 ( .A1(n1723), .A2(wrdata_d1[156]), .A3(n1759), .A4(n1635), 
        .Y(n1636) );
  AO22X1_RVT U1808 ( .A1(n1750), .A2(\inq_ary[11][157] ), .A3(n1738), .A4(
        \inq_ary[6][157] ), .Y(n1640) );
  AO22X1_RVT U1809 ( .A1(n1554), .A2(\inq_ary[14][157] ), .A3(n1748), .A4(
        \inq_ary[10][157] ), .Y(n1639) );
  AO22X1_RVT U1810 ( .A1(n1740), .A2(\inq_ary[12][157] ), .A3(n1747), .A4(
        \inq_ary[5][157] ), .Y(n1638) );
  AO22X1_RVT U1811 ( .A1(n1686), .A2(\inq_ary[0][157] ), .A3(n1741), .A4(
        \inq_ary[7][157] ), .Y(n1637) );
  NOR4X1_RVT U1812 ( .A1(n1640), .A2(n1639), .A3(n1638), .A4(n1637), .Y(n1646)
         );
  AO22X1_RVT U1813 ( .A1(n1739), .A2(\inq_ary[2][157] ), .A3(n1742), .A4(
        \inq_ary[3][157] ), .Y(n1644) );
  AO22X1_RVT U1814 ( .A1(n1711), .A2(\inq_ary[13][157] ), .A3(n1751), .A4(
        \inq_ary[9][157] ), .Y(n1643) );
  AO22X1_RVT U1815 ( .A1(n1729), .A2(\inq_ary[4][157] ), .A3(n1749), .A4(
        \inq_ary[1][157] ), .Y(n1642) );
  AO22X1_RVT U1816 ( .A1(n1537), .A2(\inq_ary[15][157] ), .A3(n1612), .A4(
        \inq_ary[8][157] ), .Y(n1641) );
  NOR4X1_RVT U1817 ( .A1(n1644), .A2(n1643), .A3(n1642), .A4(n1641), .Y(n1645)
         );
  NAND2X0_RVT U1818 ( .A1(n1646), .A2(n1645), .Y(n1647) );
  AO22X1_RVT U1819 ( .A1(n1760), .A2(wrdata_d1[157]), .A3(n1759), .A4(n1647), 
        .Y(n1648) );
  AO22X1_RVT U1820 ( .A1(n1741), .A2(\inq_ary[7][158] ), .A3(n1738), .A4(
        \inq_ary[6][158] ), .Y(n1652) );
  AO22X1_RVT U1821 ( .A1(n1537), .A2(\inq_ary[15][158] ), .A3(n1740), .A4(
        \inq_ary[12][158] ), .Y(n1651) );
  AO22X1_RVT U1822 ( .A1(n1554), .A2(\inq_ary[14][158] ), .A3(n1711), .A4(
        \inq_ary[13][158] ), .Y(n1650) );
  AO22X1_RVT U1823 ( .A1(n1739), .A2(\inq_ary[2][158] ), .A3(n1612), .A4(
        \inq_ary[8][158] ), .Y(n1649) );
  NOR4X1_RVT U1824 ( .A1(n1652), .A2(n1651), .A3(n1650), .A4(n1649), .Y(n1658)
         );
  AO22X1_RVT U1825 ( .A1(n1750), .A2(\inq_ary[11][158] ), .A3(n1751), .A4(
        \inq_ary[9][158] ), .Y(n1656) );
  AO22X1_RVT U1826 ( .A1(n1686), .A2(\inq_ary[0][158] ), .A3(n1747), .A4(
        \inq_ary[5][158] ), .Y(n1655) );
  AO22X1_RVT U1827 ( .A1(n1742), .A2(\inq_ary[3][158] ), .A3(n1748), .A4(
        \inq_ary[10][158] ), .Y(n1654) );
  AO22X1_RVT U1828 ( .A1(n1729), .A2(\inq_ary[4][158] ), .A3(n1749), .A4(
        \inq_ary[1][158] ), .Y(n1653) );
  NOR4X1_RVT U1829 ( .A1(n1656), .A2(n1655), .A3(n1654), .A4(n1653), .Y(n1657)
         );
  NAND2X0_RVT U1830 ( .A1(n1658), .A2(n1657), .Y(n1659) );
  AO22X1_RVT U1831 ( .A1(n1760), .A2(wrdata_d1[158]), .A3(n1759), .A4(n1659), 
        .Y(n1660) );
  AO22X1_RVT U1832 ( .A1(n1739), .A2(\inq_ary[2][148] ), .A3(n1747), .A4(
        \inq_ary[5][148] ), .Y(n1664) );
  AO22X1_RVT U1833 ( .A1(n1749), .A2(\inq_ary[1][148] ), .A3(n1738), .A4(
        \inq_ary[6][148] ), .Y(n1663) );
  AO22X1_RVT U1834 ( .A1(n1554), .A2(\inq_ary[14][148] ), .A3(n1741), .A4(
        \inq_ary[7][148] ), .Y(n1662) );
  AO22X1_RVT U1835 ( .A1(n1537), .A2(\inq_ary[15][148] ), .A3(n1751), .A4(
        \inq_ary[9][148] ), .Y(n1661) );
  NOR4X1_RVT U1836 ( .A1(n1664), .A2(n1663), .A3(n1662), .A4(n1661), .Y(n1670)
         );
  AO22X1_RVT U1837 ( .A1(n1750), .A2(\inq_ary[11][148] ), .A3(n1748), .A4(
        \inq_ary[10][148] ), .Y(n1668) );
  AO22X1_RVT U1838 ( .A1(n1686), .A2(\inq_ary[0][148] ), .A3(n1740), .A4(
        \inq_ary[12][148] ), .Y(n1667) );
  AO22X1_RVT U1839 ( .A1(n1612), .A2(\inq_ary[8][148] ), .A3(n1711), .A4(
        \inq_ary[13][148] ), .Y(n1666) );
  AO22X1_RVT U1840 ( .A1(n1742), .A2(\inq_ary[3][148] ), .A3(n1729), .A4(
        \inq_ary[4][148] ), .Y(n1665) );
  NOR4X1_RVT U1841 ( .A1(n1668), .A2(n1667), .A3(n1666), .A4(n1665), .Y(n1669)
         );
  NAND2X0_RVT U1842 ( .A1(n1670), .A2(n1669), .Y(n1671) );
  AO22X1_RVT U1843 ( .A1(n1684), .A2(wrdata_d1[148]), .A3(n2), .A4(n1671), .Y(
        n1672) );
  AO22X1_RVT U1844 ( .A1(n1612), .A2(\inq_ary[8][149] ), .A3(n1750), .A4(
        \inq_ary[11][149] ), .Y(n1676) );
  AO22X1_RVT U1845 ( .A1(n1741), .A2(\inq_ary[7][149] ), .A3(n1751), .A4(
        \inq_ary[9][149] ), .Y(n1675) );
  AO22X1_RVT U1846 ( .A1(n1729), .A2(\inq_ary[4][149] ), .A3(n1711), .A4(
        \inq_ary[13][149] ), .Y(n1674) );
  AO22X1_RVT U1847 ( .A1(n1749), .A2(\inq_ary[1][149] ), .A3(n1747), .A4(
        \inq_ary[5][149] ), .Y(n1673) );
  NOR4X1_RVT U1848 ( .A1(n1676), .A2(n1675), .A3(n1674), .A4(n1673), .Y(n1682)
         );
  AO22X1_RVT U1849 ( .A1(n1686), .A2(\inq_ary[0][149] ), .A3(n1748), .A4(
        \inq_ary[10][149] ), .Y(n1680) );
  AO22X1_RVT U1850 ( .A1(n1742), .A2(\inq_ary[3][149] ), .A3(n1740), .A4(
        \inq_ary[12][149] ), .Y(n1679) );
  AO22X1_RVT U1851 ( .A1(n1739), .A2(\inq_ary[2][149] ), .A3(n1554), .A4(
        \inq_ary[14][149] ), .Y(n1678) );
  AO22X1_RVT U1852 ( .A1(n1537), .A2(\inq_ary[15][149] ), .A3(n1738), .A4(
        \inq_ary[6][149] ), .Y(n1677) );
  NOR4X1_RVT U1853 ( .A1(n1680), .A2(n1679), .A3(n1678), .A4(n1677), .Y(n1681)
         );
  NAND2X0_RVT U1854 ( .A1(n1682), .A2(n1681), .Y(n1683) );
  AO22X1_RVT U1855 ( .A1(n1684), .A2(wrdata_d1[149]), .A3(n2), .A4(n1683), .Y(
        n1685) );
  AO22X1_RVT U1856 ( .A1(n1554), .A2(\inq_ary[14][150] ), .A3(n1749), .A4(
        \inq_ary[1][150] ), .Y(n1690) );
  AO22X1_RVT U1857 ( .A1(n1742), .A2(\inq_ary[3][150] ), .A3(n1740), .A4(
        \inq_ary[12][150] ), .Y(n1689) );
  AO22X1_RVT U1858 ( .A1(n1748), .A2(\inq_ary[10][150] ), .A3(n1751), .A4(
        \inq_ary[9][150] ), .Y(n1688) );
  AO22X1_RVT U1859 ( .A1(n1739), .A2(\inq_ary[2][150] ), .A3(n1686), .A4(
        \inq_ary[0][150] ), .Y(n1687) );
  NOR4X1_RVT U1860 ( .A1(n1690), .A2(n1689), .A3(n1688), .A4(n1687), .Y(n1696)
         );
  AO22X1_RVT U1861 ( .A1(n1747), .A2(\inq_ary[5][150] ), .A3(n1711), .A4(
        \inq_ary[13][150] ), .Y(n1694) );
  AO22X1_RVT U1862 ( .A1(n1750), .A2(\inq_ary[11][150] ), .A3(n1738), .A4(
        \inq_ary[6][150] ), .Y(n1693) );
  AO22X1_RVT U1863 ( .A1(n1537), .A2(\inq_ary[15][150] ), .A3(n1741), .A4(
        \inq_ary[7][150] ), .Y(n1692) );
  AO22X1_RVT U1864 ( .A1(n1729), .A2(\inq_ary[4][150] ), .A3(n1612), .A4(
        \inq_ary[8][150] ), .Y(n1691) );
  NOR4X1_RVT U1865 ( .A1(n1694), .A2(n1693), .A3(n1692), .A4(n1691), .Y(n1695)
         );
  NAND2X0_RVT U1866 ( .A1(n1696), .A2(n1695), .Y(n1697) );
  AO22X1_RVT U1867 ( .A1(n1723), .A2(wrdata_d1[150]), .A3(n2), .A4(n1697), .Y(
        n1698) );
  AO22X1_RVT U1868 ( .A1(n1739), .A2(\inq_ary[2][151] ), .A3(n1747), .A4(
        \inq_ary[5][151] ), .Y(n1702) );
  AO22X1_RVT U1869 ( .A1(n1750), .A2(\inq_ary[11][151] ), .A3(n1738), .A4(
        \inq_ary[6][151] ), .Y(n1701) );
  AO22X1_RVT U1870 ( .A1(n1612), .A2(\inq_ary[8][151] ), .A3(n1749), .A4(
        \inq_ary[1][151] ), .Y(n1700) );
  AO22X1_RVT U1871 ( .A1(n1742), .A2(\inq_ary[3][151] ), .A3(n1686), .A4(
        \inq_ary[0][151] ), .Y(n1699) );
  NOR4X1_RVT U1872 ( .A1(n1702), .A2(n1701), .A3(n1700), .A4(n1699), .Y(n1708)
         );
  AO22X1_RVT U1873 ( .A1(n1740), .A2(\inq_ary[12][151] ), .A3(n1711), .A4(
        \inq_ary[13][151] ), .Y(n1706) );
  AO22X1_RVT U1874 ( .A1(n1537), .A2(\inq_ary[15][151] ), .A3(n1748), .A4(
        \inq_ary[10][151] ), .Y(n1705) );
  AO22X1_RVT U1875 ( .A1(n1741), .A2(\inq_ary[7][151] ), .A3(n1751), .A4(
        \inq_ary[9][151] ), .Y(n1704) );
  AO22X1_RVT U1876 ( .A1(n1554), .A2(\inq_ary[14][151] ), .A3(n1729), .A4(
        \inq_ary[4][151] ), .Y(n1703) );
  NOR4X1_RVT U1877 ( .A1(n1706), .A2(n1705), .A3(n1704), .A4(n1703), .Y(n1707)
         );
  NAND2X0_RVT U1878 ( .A1(n1708), .A2(n1707), .Y(n1709) );
  AO22X1_RVT U1879 ( .A1(n1723), .A2(wrdata_d1[151]), .A3(n1759), .A4(n1709), 
        .Y(n1710) );
  AO22X1_RVT U1880 ( .A1(n1738), .A2(\inq_ary[6][152] ), .A3(n1751), .A4(
        \inq_ary[9][152] ), .Y(n1715) );
  AO22X1_RVT U1881 ( .A1(n1740), .A2(\inq_ary[12][152] ), .A3(n1750), .A4(
        \inq_ary[11][152] ), .Y(n1714) );
  AO22X1_RVT U1882 ( .A1(n1747), .A2(\inq_ary[5][152] ), .A3(n1711), .A4(
        \inq_ary[13][152] ), .Y(n1713) );
  AO22X1_RVT U1883 ( .A1(n1741), .A2(\inq_ary[7][152] ), .A3(n1748), .A4(
        \inq_ary[10][152] ), .Y(n1712) );
  NOR4X1_RVT U1884 ( .A1(n1715), .A2(n1714), .A3(n1713), .A4(n1712), .Y(n1721)
         );
  AO22X1_RVT U1885 ( .A1(n1739), .A2(\inq_ary[2][152] ), .A3(n1729), .A4(
        \inq_ary[4][152] ), .Y(n1719) );
  AO22X1_RVT U1886 ( .A1(n1537), .A2(\inq_ary[15][152] ), .A3(n1749), .A4(
        \inq_ary[1][152] ), .Y(n1718) );
  AO22X1_RVT U1887 ( .A1(n1742), .A2(\inq_ary[3][152] ), .A3(n1686), .A4(
        \inq_ary[0][152] ), .Y(n1717) );
  AO22X1_RVT U1888 ( .A1(n1554), .A2(\inq_ary[14][152] ), .A3(n1612), .A4(
        \inq_ary[8][152] ), .Y(n1716) );
  NOR4X1_RVT U1889 ( .A1(n1719), .A2(n1718), .A3(n1717), .A4(n1716), .Y(n1720)
         );
  NAND2X0_RVT U1890 ( .A1(n1721), .A2(n1720), .Y(n1722) );
  AO22X1_RVT U1891 ( .A1(n1723), .A2(wrdata_d1[152]), .A3(n1759), .A4(n1722), 
        .Y(n1724) );
  AO22X1_RVT U1892 ( .A1(n1612), .A2(\inq_ary[8][153] ), .A3(n1747), .A4(
        \inq_ary[5][153] ), .Y(n1728) );
  AO22X1_RVT U1893 ( .A1(n1739), .A2(\inq_ary[2][153] ), .A3(n1554), .A4(
        \inq_ary[14][153] ), .Y(n1727) );
  AO22X1_RVT U1894 ( .A1(n1749), .A2(\inq_ary[1][153] ), .A3(n1751), .A4(
        \inq_ary[9][153] ), .Y(n1726) );
  AO22X1_RVT U1895 ( .A1(n1740), .A2(\inq_ary[12][153] ), .A3(n1738), .A4(
        \inq_ary[6][153] ), .Y(n1725) );
  NOR4X1_RVT U1896 ( .A1(n1728), .A2(n1727), .A3(n1726), .A4(n1725), .Y(n1735)
         );
  AO22X1_RVT U1897 ( .A1(n1742), .A2(\inq_ary[3][153] ), .A3(n1741), .A4(
        \inq_ary[7][153] ), .Y(n1733) );
  AO22X1_RVT U1898 ( .A1(n1537), .A2(\inq_ary[15][153] ), .A3(n1748), .A4(
        \inq_ary[10][153] ), .Y(n1732) );
  AO22X1_RVT U1899 ( .A1(n1686), .A2(\inq_ary[0][153] ), .A3(n1711), .A4(
        \inq_ary[13][153] ), .Y(n1731) );
  AO22X1_RVT U1900 ( .A1(n1729), .A2(\inq_ary[4][153] ), .A3(n1750), .A4(
        \inq_ary[11][153] ), .Y(n1730) );
  NOR4X1_RVT U1901 ( .A1(n1733), .A2(n1732), .A3(n1731), .A4(n1730), .Y(n1734)
         );
  NAND2X0_RVT U1902 ( .A1(n1735), .A2(n1734), .Y(n1736) );
  AO22X1_RVT U1903 ( .A1(n1760), .A2(wrdata_d1[153]), .A3(n1759), .A4(n1736), 
        .Y(n1737) );
  AO22X1_RVT U1904 ( .A1(n1739), .A2(\inq_ary[2][159] ), .A3(n1738), .A4(
        \inq_ary[6][159] ), .Y(n1746) );
  AO22X1_RVT U1905 ( .A1(n1612), .A2(\inq_ary[8][159] ), .A3(n1740), .A4(
        \inq_ary[12][159] ), .Y(n1745) );
  AO22X1_RVT U1906 ( .A1(n1729), .A2(\inq_ary[4][159] ), .A3(n1711), .A4(
        \inq_ary[13][159] ), .Y(n1744) );
  AO22X1_RVT U1907 ( .A1(n1742), .A2(\inq_ary[3][159] ), .A3(n1741), .A4(
        \inq_ary[7][159] ), .Y(n1743) );
  NOR4X1_RVT U1908 ( .A1(n1746), .A2(n1745), .A3(n1744), .A4(n1743), .Y(n1757)
         );
  AO22X1_RVT U1909 ( .A1(n1537), .A2(\inq_ary[15][159] ), .A3(n1747), .A4(
        \inq_ary[5][159] ), .Y(n1755) );
  AO22X1_RVT U1910 ( .A1(n1749), .A2(\inq_ary[1][159] ), .A3(n1748), .A4(
        \inq_ary[10][159] ), .Y(n1754) );
  AO22X1_RVT U1911 ( .A1(n1686), .A2(\inq_ary[0][159] ), .A3(n1750), .A4(
        \inq_ary[11][159] ), .Y(n1753) );
  AO22X1_RVT U1912 ( .A1(n1554), .A2(\inq_ary[14][159] ), .A3(n1751), .A4(
        \inq_ary[9][159] ), .Y(n1752) );
  NOR4X1_RVT U1913 ( .A1(n1755), .A2(n1754), .A3(n1753), .A4(n1752), .Y(n1756)
         );
  NAND2X0_RVT U1914 ( .A1(n1757), .A2(n1756), .Y(n1758) );
  AO22X1_RVT U1915 ( .A1(n1760), .A2(wrdata_d1[159]), .A3(n1759), .A4(n1758), 
        .Y(n1761) );
  AND2X1_RVT U1917 ( .A1(reset_l), .A2(rdptr_d1[2]), .Y(n1762) );
  AND4X1_RVT U1918 ( .A1(rdptr_d1[1]), .A2(n1762), .A3(rdptr_d1[3]), .A4(
        rdptr_d1[0]), .Y(n3312) );
  AND3X1_RVT U1919 ( .A1(reset_l), .A2(rdptr_d1[2]), .A3(n3337), .Y(n1768) );
  AND3X1_RVT U1920 ( .A1(rdptr_d1[3]), .A2(n1768), .A3(n3334), .Y(n3303) );
  AO22X1_RVT U1921 ( .A1(\inq_ary[15][5] ), .A2(n3312), .A3(\inq_ary[12][5] ), 
        .A4(n3303), .Y(n1766) );
  AND3X1_RVT U1922 ( .A1(n5), .A2(n3334), .A3(n1768), .Y(n3321) );
  AND2X1_RVT U1923 ( .A1(reset_l), .A2(n3338), .Y(n1770) );
  AND2X1_RVT U1924 ( .A1(n1770), .A2(n3337), .Y(n1767) );
  AND3X1_RVT U1925 ( .A1(rdptr_d1[3]), .A2(n1767), .A3(n3334), .Y(n3313) );
  AO22X1_RVT U1926 ( .A1(\inq_ary[4][5] ), .A2(n3321), .A3(\inq_ary[8][5] ), 
        .A4(n3313), .Y(n1765) );
  AND4X1_RVT U1927 ( .A1(n1762), .A2(rdptr_d1[1]), .A3(rdptr_d1[3]), .A4(n3334), .Y(n3325) );
  AND3X1_RVT U1928 ( .A1(rdptr_d1[0]), .A2(n1767), .A3(n5), .Y(n3324) );
  AO22X1_RVT U1929 ( .A1(\inq_ary[14][5] ), .A2(n3325), .A3(\inq_ary[1][5] ), 
        .A4(n3324), .Y(n1764) );
  AND4X1_RVT U1930 ( .A1(n1762), .A2(rdptr_d1[1]), .A3(rdptr_d1[0]), .A4(n5), 
        .Y(n3322) );
  AND4X1_RVT U1931 ( .A1(rdptr_d1[3]), .A2(rdptr_d1[1]), .A3(n1770), .A4(n3334), .Y(n3326) );
  AO22X1_RVT U1932 ( .A1(\inq_ary[7][5] ), .A2(n3322), .A3(\inq_ary[10][5] ), 
        .A4(n3326), .Y(n1763) );
  NOR4X1_RVT U1933 ( .A1(n1766), .A2(n1765), .A3(n1764), .A4(n1763), .Y(n1776)
         );
  AND3X1_RVT U1934 ( .A1(n5), .A2(n3334), .A3(n1767), .Y(n3315) );
  AND3X1_RVT U1935 ( .A1(rdptr_d1[3]), .A2(rdptr_d1[0]), .A3(n1767), .Y(n3314)
         );
  AO22X1_RVT U1936 ( .A1(\inq_ary[0][5] ), .A2(n3315), .A3(\inq_ary[9][5] ), 
        .A4(n3314), .Y(n1774) );
  AND3X1_RVT U1937 ( .A1(n1768), .A2(rdptr_d1[0]), .A3(n5), .Y(n3298) );
  AND3X1_RVT U1938 ( .A1(n1768), .A2(rdptr_d1[3]), .A3(rdptr_d1[0]), .Y(n3323)
         );
  AO22X1_RVT U1939 ( .A1(\inq_ary[5][5] ), .A2(n3298), .A3(\inq_ary[13][5] ), 
        .A4(n3323), .Y(n1773) );
  AND4X1_RVT U1940 ( .A1(rdptr_d1[1]), .A2(rdptr_d1[0]), .A3(n1770), .A4(n5), 
        .Y(n3310) );
  AND2X1_RVT U1941 ( .A1(n5), .A2(n3334), .Y(n1769) );
  AND4X1_RVT U1942 ( .A1(rdptr_d1[1]), .A2(reset_l), .A3(rdptr_d1[2]), .A4(
        n1769), .Y(n3311) );
  AO22X1_RVT U1943 ( .A1(\inq_ary[3][5] ), .A2(n3310), .A3(\inq_ary[6][5] ), 
        .A4(n3311), .Y(n1772) );
  AND4X1_RVT U1944 ( .A1(rdptr_d1[1]), .A2(n1770), .A3(n3334), .A4(n5), .Y(
        n3271) );
  AND4X1_RVT U1945 ( .A1(rdptr_d1[1]), .A2(rdptr_d1[3]), .A3(rdptr_d1[0]), 
        .A4(n1770), .Y(n3316) );
  AO22X1_RVT U1946 ( .A1(\inq_ary[2][5] ), .A2(n3271), .A3(\inq_ary[11][5] ), 
        .A4(n3316), .Y(n1771) );
  NOR4X1_RVT U1947 ( .A1(n1774), .A2(n1773), .A3(n1772), .A4(n1771), .Y(n1775)
         );
  NAND2X0_RVT U1948 ( .A1(n1776), .A2(n1775), .Y(N266) );
  AO22X1_RVT U1949 ( .A1(\inq_ary[11][6] ), .A2(n3316), .A3(\inq_ary[10][6] ), 
        .A4(n3326), .Y(n1780) );
  AO22X1_RVT U1950 ( .A1(\inq_ary[3][6] ), .A2(n3310), .A3(\inq_ary[5][6] ), 
        .A4(n3298), .Y(n1779) );
  AO22X1_RVT U1951 ( .A1(\inq_ary[8][6] ), .A2(n3313), .A3(\inq_ary[9][6] ), 
        .A4(n3314), .Y(n1778) );
  AO22X1_RVT U1952 ( .A1(\inq_ary[15][6] ), .A2(n3312), .A3(\inq_ary[2][6] ), 
        .A4(n3271), .Y(n1777) );
  NOR4X1_RVT U1953 ( .A1(n1780), .A2(n1779), .A3(n1778), .A4(n1777), .Y(n1786)
         );
  AO22X1_RVT U1954 ( .A1(\inq_ary[12][6] ), .A2(n3303), .A3(\inq_ary[1][6] ), 
        .A4(n3324), .Y(n1784) );
  AO22X1_RVT U1955 ( .A1(\inq_ary[4][6] ), .A2(n3321), .A3(\inq_ary[6][6] ), 
        .A4(n3311), .Y(n1783) );
  AO22X1_RVT U1956 ( .A1(\inq_ary[13][6] ), .A2(n3323), .A3(\inq_ary[0][6] ), 
        .A4(n3315), .Y(n1782) );
  AO22X1_RVT U1957 ( .A1(\inq_ary[7][6] ), .A2(n3322), .A3(\inq_ary[14][6] ), 
        .A4(n3325), .Y(n1781) );
  NOR4X1_RVT U1958 ( .A1(n1784), .A2(n1783), .A3(n1782), .A4(n1781), .Y(n1785)
         );
  NAND2X0_RVT U1959 ( .A1(n1786), .A2(n1785), .Y(N267) );
  AO22X1_RVT U1960 ( .A1(\inq_ary[11][7] ), .A2(n3316), .A3(\inq_ary[3][7] ), 
        .A4(n3310), .Y(n1790) );
  AO22X1_RVT U1961 ( .A1(\inq_ary[0][7] ), .A2(n3315), .A3(\inq_ary[10][7] ), 
        .A4(n3326), .Y(n1789) );
  AO22X1_RVT U1962 ( .A1(\inq_ary[13][7] ), .A2(n3323), .A3(\inq_ary[14][7] ), 
        .A4(n3325), .Y(n1788) );
  AO22X1_RVT U1963 ( .A1(\inq_ary[9][7] ), .A2(n3314), .A3(\inq_ary[4][7] ), 
        .A4(n3321), .Y(n1787) );
  NOR4X1_RVT U1964 ( .A1(n1790), .A2(n1789), .A3(n1788), .A4(n1787), .Y(n1796)
         );
  AO22X1_RVT U1965 ( .A1(\inq_ary[7][7] ), .A2(n3322), .A3(\inq_ary[8][7] ), 
        .A4(n3313), .Y(n1794) );
  AO22X1_RVT U1966 ( .A1(\inq_ary[15][7] ), .A2(n3312), .A3(\inq_ary[5][7] ), 
        .A4(n3298), .Y(n1793) );
  AO22X1_RVT U1967 ( .A1(\inq_ary[6][7] ), .A2(n3311), .A3(\inq_ary[2][7] ), 
        .A4(n3271), .Y(n1792) );
  AO22X1_RVT U1968 ( .A1(\inq_ary[1][7] ), .A2(n3324), .A3(\inq_ary[12][7] ), 
        .A4(n3303), .Y(n1791) );
  NOR4X1_RVT U1969 ( .A1(n1794), .A2(n1793), .A3(n1792), .A4(n1791), .Y(n1795)
         );
  NAND2X0_RVT U1970 ( .A1(n1796), .A2(n1795), .Y(N268) );
  AO22X1_RVT U1971 ( .A1(\inq_ary[8][8] ), .A2(n3313), .A3(\inq_ary[2][8] ), 
        .A4(n3271), .Y(n1800) );
  AO22X1_RVT U1972 ( .A1(\inq_ary[6][8] ), .A2(n3311), .A3(\inq_ary[5][8] ), 
        .A4(n3298), .Y(n1799) );
  AO22X1_RVT U1973 ( .A1(\inq_ary[11][8] ), .A2(n3316), .A3(\inq_ary[12][8] ), 
        .A4(n3303), .Y(n1798) );
  AO22X1_RVT U1974 ( .A1(\inq_ary[13][8] ), .A2(n3323), .A3(\inq_ary[1][8] ), 
        .A4(n3324), .Y(n1797) );
  NOR4X1_RVT U1975 ( .A1(n1800), .A2(n1799), .A3(n1798), .A4(n1797), .Y(n1806)
         );
  AO22X1_RVT U1976 ( .A1(\inq_ary[4][8] ), .A2(n3321), .A3(\inq_ary[10][8] ), 
        .A4(n3326), .Y(n1804) );
  AO22X1_RVT U1977 ( .A1(\inq_ary[15][8] ), .A2(n3312), .A3(\inq_ary[0][8] ), 
        .A4(n3315), .Y(n1803) );
  AO22X1_RVT U1978 ( .A1(\inq_ary[14][8] ), .A2(n3325), .A3(\inq_ary[7][8] ), 
        .A4(n3322), .Y(n1802) );
  AO22X1_RVT U1979 ( .A1(\inq_ary[9][8] ), .A2(n3314), .A3(\inq_ary[3][8] ), 
        .A4(n3310), .Y(n1801) );
  NOR4X1_RVT U1980 ( .A1(n1804), .A2(n1803), .A3(n1802), .A4(n1801), .Y(n1805)
         );
  NAND2X0_RVT U1981 ( .A1(n1806), .A2(n1805), .Y(N269) );
  AO22X1_RVT U1982 ( .A1(\inq_ary[13][9] ), .A2(n3323), .A3(\inq_ary[10][9] ), 
        .A4(n3326), .Y(n1810) );
  AO22X1_RVT U1983 ( .A1(\inq_ary[4][9] ), .A2(n3321), .A3(\inq_ary[6][9] ), 
        .A4(n3311), .Y(n1809) );
  AO22X1_RVT U1984 ( .A1(\inq_ary[7][9] ), .A2(n3322), .A3(\inq_ary[2][9] ), 
        .A4(n3271), .Y(n1808) );
  AO22X1_RVT U1985 ( .A1(\inq_ary[9][9] ), .A2(n3314), .A3(\inq_ary[5][9] ), 
        .A4(n3298), .Y(n1807) );
  NOR4X1_RVT U1986 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .Y(n1816)
         );
  AO22X1_RVT U1987 ( .A1(\inq_ary[1][9] ), .A2(n3324), .A3(\inq_ary[12][9] ), 
        .A4(n3303), .Y(n1814) );
  AO22X1_RVT U1988 ( .A1(\inq_ary[14][9] ), .A2(n3325), .A3(\inq_ary[15][9] ), 
        .A4(n3312), .Y(n1813) );
  AO22X1_RVT U1989 ( .A1(\inq_ary[3][9] ), .A2(n3310), .A3(\inq_ary[0][9] ), 
        .A4(n3315), .Y(n1812) );
  AO22X1_RVT U1990 ( .A1(\inq_ary[8][9] ), .A2(n3313), .A3(\inq_ary[11][9] ), 
        .A4(n3316), .Y(n1811) );
  NOR4X1_RVT U1991 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .Y(n1815)
         );
  NAND2X0_RVT U1992 ( .A1(n1816), .A2(n1815), .Y(N270) );
  AO22X1_RVT U1993 ( .A1(\inq_ary[10][10] ), .A2(n3326), .A3(\inq_ary[12][10] ), .A4(n3303), .Y(n1820) );
  AO22X1_RVT U1994 ( .A1(\inq_ary[7][10] ), .A2(n3322), .A3(\inq_ary[9][10] ), 
        .A4(n3314), .Y(n1819) );
  AO22X1_RVT U1995 ( .A1(\inq_ary[11][10] ), .A2(n3316), .A3(\inq_ary[5][10] ), 
        .A4(n3298), .Y(n1818) );
  AO22X1_RVT U1996 ( .A1(\inq_ary[2][10] ), .A2(n3271), .A3(\inq_ary[14][10] ), 
        .A4(n3325), .Y(n1817) );
  NOR4X1_RVT U1997 ( .A1(n1820), .A2(n1819), .A3(n1818), .A4(n1817), .Y(n1826)
         );
  AO22X1_RVT U1998 ( .A1(\inq_ary[3][10] ), .A2(n3310), .A3(\inq_ary[4][10] ), 
        .A4(n3321), .Y(n1824) );
  AO22X1_RVT U1999 ( .A1(\inq_ary[1][10] ), .A2(n3324), .A3(\inq_ary[15][10] ), 
        .A4(n3312), .Y(n1823) );
  AO22X1_RVT U2000 ( .A1(\inq_ary[6][10] ), .A2(n3311), .A3(\inq_ary[0][10] ), 
        .A4(n3315), .Y(n1822) );
  AO22X1_RVT U2001 ( .A1(\inq_ary[8][10] ), .A2(n3313), .A3(\inq_ary[13][10] ), 
        .A4(n3323), .Y(n1821) );
  NOR4X1_RVT U2002 ( .A1(n1824), .A2(n1823), .A3(n1822), .A4(n1821), .Y(n1825)
         );
  NAND2X0_RVT U2003 ( .A1(n1826), .A2(n1825), .Y(N271) );
  AO22X1_RVT U2004 ( .A1(\inq_ary[9][11] ), .A2(n3314), .A3(\inq_ary[6][11] ), 
        .A4(n3311), .Y(n1830) );
  AO22X1_RVT U2005 ( .A1(\inq_ary[13][11] ), .A2(n3323), .A3(\inq_ary[11][11] ), .A4(n3316), .Y(n1829) );
  AO22X1_RVT U2006 ( .A1(\inq_ary[4][11] ), .A2(n3321), .A3(\inq_ary[0][11] ), 
        .A4(n3315), .Y(n1828) );
  AO22X1_RVT U2007 ( .A1(\inq_ary[5][11] ), .A2(n3298), .A3(\inq_ary[10][11] ), 
        .A4(n3326), .Y(n1827) );
  NOR4X1_RVT U2008 ( .A1(n1830), .A2(n1829), .A3(n1828), .A4(n1827), .Y(n1836)
         );
  AO22X1_RVT U2009 ( .A1(\inq_ary[14][11] ), .A2(n3325), .A3(\inq_ary[8][11] ), 
        .A4(n3313), .Y(n1834) );
  AO22X1_RVT U2010 ( .A1(\inq_ary[2][11] ), .A2(n3271), .A3(\inq_ary[3][11] ), 
        .A4(n3310), .Y(n1833) );
  AO22X1_RVT U2011 ( .A1(\inq_ary[7][11] ), .A2(n3322), .A3(\inq_ary[12][11] ), 
        .A4(n3303), .Y(n1832) );
  AO22X1_RVT U2012 ( .A1(\inq_ary[1][11] ), .A2(n3324), .A3(\inq_ary[15][11] ), 
        .A4(n3312), .Y(n1831) );
  NOR4X1_RVT U2013 ( .A1(n1834), .A2(n1833), .A3(n1832), .A4(n1831), .Y(n1835)
         );
  NAND2X0_RVT U2014 ( .A1(n1836), .A2(n1835), .Y(N272) );
  AO22X1_RVT U2015 ( .A1(\inq_ary[3][12] ), .A2(n3310), .A3(\inq_ary[14][12] ), 
        .A4(n3325), .Y(n1840) );
  AO22X1_RVT U2016 ( .A1(\inq_ary[15][12] ), .A2(n3312), .A3(\inq_ary[4][12] ), 
        .A4(n3321), .Y(n1839) );
  AO22X1_RVT U2017 ( .A1(\inq_ary[9][12] ), .A2(n3314), .A3(\inq_ary[5][12] ), 
        .A4(n3298), .Y(n1838) );
  AO22X1_RVT U2018 ( .A1(\inq_ary[12][12] ), .A2(n3303), .A3(\inq_ary[2][12] ), 
        .A4(n3271), .Y(n1837) );
  NOR4X1_RVT U2019 ( .A1(n1840), .A2(n1839), .A3(n1838), .A4(n1837), .Y(n1846)
         );
  AO22X1_RVT U2020 ( .A1(\inq_ary[10][12] ), .A2(n3326), .A3(\inq_ary[1][12] ), 
        .A4(n3324), .Y(n1844) );
  AO22X1_RVT U2021 ( .A1(\inq_ary[11][12] ), .A2(n3316), .A3(\inq_ary[8][12] ), 
        .A4(n3313), .Y(n1843) );
  AO22X1_RVT U2022 ( .A1(\inq_ary[0][12] ), .A2(n3315), .A3(\inq_ary[6][12] ), 
        .A4(n3311), .Y(n1842) );
  AO22X1_RVT U2023 ( .A1(\inq_ary[13][12] ), .A2(n3323), .A3(\inq_ary[7][12] ), 
        .A4(n3322), .Y(n1841) );
  NOR4X1_RVT U2024 ( .A1(n1844), .A2(n1843), .A3(n1842), .A4(n1841), .Y(n1845)
         );
  NAND2X0_RVT U2025 ( .A1(n1846), .A2(n1845), .Y(N273) );
  AO22X1_RVT U2026 ( .A1(\inq_ary[9][13] ), .A2(n3314), .A3(\inq_ary[12][13] ), 
        .A4(n3303), .Y(n1850) );
  AO22X1_RVT U2027 ( .A1(\inq_ary[4][13] ), .A2(n3321), .A3(\inq_ary[0][13] ), 
        .A4(n3315), .Y(n1849) );
  AO22X1_RVT U2028 ( .A1(\inq_ary[15][13] ), .A2(n3312), .A3(\inq_ary[10][13] ), .A4(n3326), .Y(n1848) );
  AO22X1_RVT U2029 ( .A1(\inq_ary[3][13] ), .A2(n3310), .A3(\inq_ary[11][13] ), 
        .A4(n3316), .Y(n1847) );
  NOR4X1_RVT U2030 ( .A1(n1850), .A2(n1849), .A3(n1848), .A4(n1847), .Y(n1856)
         );
  AO22X1_RVT U2031 ( .A1(\inq_ary[2][13] ), .A2(n3271), .A3(\inq_ary[1][13] ), 
        .A4(n3324), .Y(n1854) );
  AO22X1_RVT U2032 ( .A1(\inq_ary[14][13] ), .A2(n3325), .A3(\inq_ary[8][13] ), 
        .A4(n3313), .Y(n1853) );
  AO22X1_RVT U2033 ( .A1(\inq_ary[5][13] ), .A2(n3298), .A3(\inq_ary[7][13] ), 
        .A4(n3322), .Y(n1852) );
  AO22X1_RVT U2034 ( .A1(\inq_ary[13][13] ), .A2(n3323), .A3(\inq_ary[6][13] ), 
        .A4(n3311), .Y(n1851) );
  NOR4X1_RVT U2035 ( .A1(n1854), .A2(n1853), .A3(n1852), .A4(n1851), .Y(n1855)
         );
  NAND2X0_RVT U2036 ( .A1(n1856), .A2(n1855), .Y(N274) );
  AO22X1_RVT U2037 ( .A1(\inq_ary[0][14] ), .A2(n3315), .A3(\inq_ary[3][14] ), 
        .A4(n3310), .Y(n1860) );
  AO22X1_RVT U2038 ( .A1(\inq_ary[4][14] ), .A2(n3321), .A3(\inq_ary[11][14] ), 
        .A4(n3316), .Y(n1859) );
  AO22X1_RVT U2039 ( .A1(\inq_ary[2][14] ), .A2(n3271), .A3(\inq_ary[6][14] ), 
        .A4(n3311), .Y(n1858) );
  AO22X1_RVT U2040 ( .A1(\inq_ary[15][14] ), .A2(n3312), .A3(\inq_ary[7][14] ), 
        .A4(n3322), .Y(n1857) );
  NOR4X1_RVT U2041 ( .A1(n1860), .A2(n1859), .A3(n1858), .A4(n1857), .Y(n1866)
         );
  AO22X1_RVT U2042 ( .A1(\inq_ary[13][14] ), .A2(n3323), .A3(\inq_ary[10][14] ), .A4(n3326), .Y(n1864) );
  AO22X1_RVT U2043 ( .A1(\inq_ary[8][14] ), .A2(n3313), .A3(\inq_ary[12][14] ), 
        .A4(n3303), .Y(n1863) );
  AO22X1_RVT U2044 ( .A1(\inq_ary[1][14] ), .A2(n3324), .A3(\inq_ary[14][14] ), 
        .A4(n3325), .Y(n1862) );
  AO22X1_RVT U2045 ( .A1(\inq_ary[5][14] ), .A2(n3298), .A3(\inq_ary[9][14] ), 
        .A4(n3314), .Y(n1861) );
  NOR4X1_RVT U2046 ( .A1(n1864), .A2(n1863), .A3(n1862), .A4(n1861), .Y(n1865)
         );
  NAND2X0_RVT U2047 ( .A1(n1866), .A2(n1865), .Y(N275) );
  AO22X1_RVT U2048 ( .A1(\inq_ary[10][15] ), .A2(n3326), .A3(\inq_ary[7][15] ), 
        .A4(n3322), .Y(n1870) );
  AO22X1_RVT U2049 ( .A1(\inq_ary[2][15] ), .A2(n3271), .A3(\inq_ary[1][15] ), 
        .A4(n3324), .Y(n1869) );
  AO22X1_RVT U2050 ( .A1(\inq_ary[0][15] ), .A2(n3315), .A3(\inq_ary[3][15] ), 
        .A4(n3310), .Y(n1868) );
  AO22X1_RVT U2051 ( .A1(\inq_ary[13][15] ), .A2(n3323), .A3(\inq_ary[6][15] ), 
        .A4(n3311), .Y(n1867) );
  NOR4X1_RVT U2052 ( .A1(n1870), .A2(n1869), .A3(n1868), .A4(n1867), .Y(n1876)
         );
  AO22X1_RVT U2053 ( .A1(\inq_ary[9][15] ), .A2(n3314), .A3(\inq_ary[4][15] ), 
        .A4(n3321), .Y(n1874) );
  AO22X1_RVT U2054 ( .A1(\inq_ary[11][15] ), .A2(n3316), .A3(\inq_ary[15][15] ), .A4(n3312), .Y(n1873) );
  AO22X1_RVT U2055 ( .A1(\inq_ary[12][15] ), .A2(n3303), .A3(\inq_ary[8][15] ), 
        .A4(n3313), .Y(n1872) );
  AO22X1_RVT U2056 ( .A1(\inq_ary[14][15] ), .A2(n3325), .A3(\inq_ary[5][15] ), 
        .A4(n3298), .Y(n1871) );
  NOR4X1_RVT U2057 ( .A1(n1874), .A2(n1873), .A3(n1872), .A4(n1871), .Y(n1875)
         );
  NAND2X0_RVT U2058 ( .A1(n1876), .A2(n1875), .Y(N276) );
  AO22X1_RVT U2059 ( .A1(\inq_ary[11][16] ), .A2(n3316), .A3(\inq_ary[4][16] ), 
        .A4(n3321), .Y(n1880) );
  AO22X1_RVT U2060 ( .A1(\inq_ary[14][16] ), .A2(n3325), .A3(\inq_ary[9][16] ), 
        .A4(n3314), .Y(n1879) );
  AO22X1_RVT U2061 ( .A1(\inq_ary[13][16] ), .A2(n3323), .A3(\inq_ary[12][16] ), .A4(n3303), .Y(n1878) );
  AO22X1_RVT U2062 ( .A1(\inq_ary[3][16] ), .A2(n3310), .A3(\inq_ary[5][16] ), 
        .A4(n3298), .Y(n1877) );
  NOR4X1_RVT U2063 ( .A1(n1880), .A2(n1879), .A3(n1878), .A4(n1877), .Y(n1886)
         );
  AO22X1_RVT U2064 ( .A1(\inq_ary[15][16] ), .A2(n3312), .A3(\inq_ary[0][16] ), 
        .A4(n3315), .Y(n1884) );
  AO22X1_RVT U2065 ( .A1(\inq_ary[10][16] ), .A2(n3326), .A3(\inq_ary[2][16] ), 
        .A4(n3271), .Y(n1883) );
  AO22X1_RVT U2066 ( .A1(\inq_ary[8][16] ), .A2(n3313), .A3(\inq_ary[6][16] ), 
        .A4(n3311), .Y(n1882) );
  AO22X1_RVT U2067 ( .A1(\inq_ary[7][16] ), .A2(n3322), .A3(\inq_ary[1][16] ), 
        .A4(n3324), .Y(n1881) );
  NOR4X1_RVT U2068 ( .A1(n1884), .A2(n1883), .A3(n1882), .A4(n1881), .Y(n1885)
         );
  NAND2X0_RVT U2069 ( .A1(n1886), .A2(n1885), .Y(N277) );
  AO22X1_RVT U2070 ( .A1(\inq_ary[8][17] ), .A2(n3313), .A3(\inq_ary[4][17] ), 
        .A4(n3321), .Y(n1890) );
  AO22X1_RVT U2071 ( .A1(\inq_ary[10][17] ), .A2(n3326), .A3(\inq_ary[2][17] ), 
        .A4(n3271), .Y(n1889) );
  AO22X1_RVT U2072 ( .A1(\inq_ary[3][17] ), .A2(n3310), .A3(\inq_ary[0][17] ), 
        .A4(n3315), .Y(n1888) );
  AO22X1_RVT U2073 ( .A1(\inq_ary[6][17] ), .A2(n3311), .A3(\inq_ary[9][17] ), 
        .A4(n3314), .Y(n1887) );
  NOR4X1_RVT U2074 ( .A1(n1890), .A2(n1889), .A3(n1888), .A4(n1887), .Y(n1896)
         );
  AO22X1_RVT U2075 ( .A1(\inq_ary[11][17] ), .A2(n3316), .A3(\inq_ary[13][17] ), .A4(n3323), .Y(n1894) );
  AO22X1_RVT U2076 ( .A1(\inq_ary[1][17] ), .A2(n3324), .A3(\inq_ary[12][17] ), 
        .A4(n3303), .Y(n1893) );
  AO22X1_RVT U2077 ( .A1(\inq_ary[15][17] ), .A2(n3312), .A3(\inq_ary[14][17] ), .A4(n3325), .Y(n1892) );
  AO22X1_RVT U2078 ( .A1(\inq_ary[7][17] ), .A2(n3322), .A3(\inq_ary[5][17] ), 
        .A4(n3298), .Y(n1891) );
  NOR4X1_RVT U2079 ( .A1(n1894), .A2(n1893), .A3(n1892), .A4(n1891), .Y(n1895)
         );
  NAND2X0_RVT U2080 ( .A1(n1896), .A2(n1895), .Y(N278) );
  AO22X1_RVT U2081 ( .A1(\inq_ary[8][18] ), .A2(n3313), .A3(\inq_ary[13][18] ), 
        .A4(n3323), .Y(n1900) );
  AO22X1_RVT U2082 ( .A1(\inq_ary[14][18] ), .A2(n3325), .A3(\inq_ary[10][18] ), .A4(n3326), .Y(n1899) );
  AO22X1_RVT U2083 ( .A1(\inq_ary[1][18] ), .A2(n3324), .A3(\inq_ary[15][18] ), 
        .A4(n3312), .Y(n1898) );
  AO22X1_RVT U2084 ( .A1(\inq_ary[7][18] ), .A2(n3322), .A3(\inq_ary[2][18] ), 
        .A4(n3271), .Y(n1897) );
  NOR4X1_RVT U2085 ( .A1(n1900), .A2(n1899), .A3(n1898), .A4(n1897), .Y(n1906)
         );
  AO22X1_RVT U2086 ( .A1(\inq_ary[3][18] ), .A2(n3310), .A3(\inq_ary[5][18] ), 
        .A4(n3298), .Y(n1904) );
  AO22X1_RVT U2087 ( .A1(\inq_ary[12][18] ), .A2(n3303), .A3(\inq_ary[4][18] ), 
        .A4(n3321), .Y(n1903) );
  AO22X1_RVT U2088 ( .A1(\inq_ary[0][18] ), .A2(n3315), .A3(\inq_ary[6][18] ), 
        .A4(n3311), .Y(n1902) );
  AO22X1_RVT U2089 ( .A1(\inq_ary[11][18] ), .A2(n3316), .A3(\inq_ary[9][18] ), 
        .A4(n3314), .Y(n1901) );
  NOR4X1_RVT U2090 ( .A1(n1904), .A2(n1903), .A3(n1902), .A4(n1901), .Y(n1905)
         );
  NAND2X0_RVT U2091 ( .A1(n1906), .A2(n1905), .Y(N279) );
  AO22X1_RVT U2092 ( .A1(\inq_ary[6][19] ), .A2(n3311), .A3(\inq_ary[5][19] ), 
        .A4(n3298), .Y(n1910) );
  AO22X1_RVT U2093 ( .A1(\inq_ary[9][19] ), .A2(n3314), .A3(\inq_ary[0][19] ), 
        .A4(n3315), .Y(n1909) );
  AO22X1_RVT U2094 ( .A1(\inq_ary[4][19] ), .A2(n3321), .A3(\inq_ary[8][19] ), 
        .A4(n3313), .Y(n1908) );
  AO22X1_RVT U2095 ( .A1(\inq_ary[11][19] ), .A2(n3316), .A3(\inq_ary[13][19] ), .A4(n3323), .Y(n1907) );
  NOR4X1_RVT U2096 ( .A1(n1910), .A2(n1909), .A3(n1908), .A4(n1907), .Y(n1916)
         );
  AO22X1_RVT U2097 ( .A1(\inq_ary[7][19] ), .A2(n3322), .A3(\inq_ary[3][19] ), 
        .A4(n3310), .Y(n1914) );
  AO22X1_RVT U2098 ( .A1(\inq_ary[14][19] ), .A2(n3325), .A3(\inq_ary[2][19] ), 
        .A4(n3271), .Y(n1913) );
  AO22X1_RVT U2099 ( .A1(\inq_ary[15][19] ), .A2(n3312), .A3(\inq_ary[10][19] ), .A4(n3326), .Y(n1912) );
  AO22X1_RVT U2100 ( .A1(\inq_ary[1][19] ), .A2(n3324), .A3(\inq_ary[12][19] ), 
        .A4(n3303), .Y(n1911) );
  NOR4X1_RVT U2101 ( .A1(n1914), .A2(n1913), .A3(n1912), .A4(n1911), .Y(n1915)
         );
  NAND2X0_RVT U2102 ( .A1(n1916), .A2(n1915), .Y(N280) );
  AO22X1_RVT U2103 ( .A1(\inq_ary[0][20] ), .A2(n3315), .A3(\inq_ary[14][20] ), 
        .A4(n3325), .Y(n1920) );
  AO22X1_RVT U2104 ( .A1(\inq_ary[7][20] ), .A2(n3322), .A3(\inq_ary[4][20] ), 
        .A4(n3321), .Y(n1919) );
  AO22X1_RVT U2105 ( .A1(\inq_ary[15][20] ), .A2(n3312), .A3(\inq_ary[1][20] ), 
        .A4(n3324), .Y(n1918) );
  AO22X1_RVT U2106 ( .A1(\inq_ary[12][20] ), .A2(n3303), .A3(\inq_ary[10][20] ), .A4(n3326), .Y(n1917) );
  NOR4X1_RVT U2107 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), .Y(n1926)
         );
  AO22X1_RVT U2108 ( .A1(\inq_ary[3][20] ), .A2(n3310), .A3(\inq_ary[13][20] ), 
        .A4(n3323), .Y(n1924) );
  AO22X1_RVT U2109 ( .A1(\inq_ary[5][20] ), .A2(n3298), .A3(\inq_ary[9][20] ), 
        .A4(n3314), .Y(n1923) );
  AO22X1_RVT U2110 ( .A1(\inq_ary[6][20] ), .A2(n3311), .A3(\inq_ary[2][20] ), 
        .A4(n3271), .Y(n1922) );
  AO22X1_RVT U2111 ( .A1(\inq_ary[8][20] ), .A2(n3313), .A3(\inq_ary[11][20] ), 
        .A4(n3316), .Y(n1921) );
  NOR4X1_RVT U2112 ( .A1(n1924), .A2(n1923), .A3(n1922), .A4(n1921), .Y(n1925)
         );
  NAND2X0_RVT U2113 ( .A1(n1926), .A2(n1925), .Y(N281) );
  AO22X1_RVT U2114 ( .A1(\inq_ary[3][21] ), .A2(n3310), .A3(\inq_ary[11][21] ), 
        .A4(n3316), .Y(n1930) );
  AO22X1_RVT U2115 ( .A1(\inq_ary[12][21] ), .A2(n3303), .A3(\inq_ary[7][21] ), 
        .A4(n3322), .Y(n1929) );
  AO22X1_RVT U2116 ( .A1(\inq_ary[10][21] ), .A2(n3326), .A3(\inq_ary[9][21] ), 
        .A4(n3314), .Y(n1928) );
  AO22X1_RVT U2117 ( .A1(\inq_ary[1][21] ), .A2(n3324), .A3(\inq_ary[5][21] ), 
        .A4(n3298), .Y(n1927) );
  NOR4X1_RVT U2118 ( .A1(n1930), .A2(n1929), .A3(n1928), .A4(n1927), .Y(n1936)
         );
  AO22X1_RVT U2119 ( .A1(\inq_ary[13][21] ), .A2(n3323), .A3(\inq_ary[2][21] ), 
        .A4(n3271), .Y(n1934) );
  AO22X1_RVT U2120 ( .A1(\inq_ary[14][21] ), .A2(n3325), .A3(\inq_ary[6][21] ), 
        .A4(n3311), .Y(n1933) );
  AO22X1_RVT U2121 ( .A1(\inq_ary[8][21] ), .A2(n3313), .A3(\inq_ary[15][21] ), 
        .A4(n3312), .Y(n1932) );
  AO22X1_RVT U2122 ( .A1(\inq_ary[4][21] ), .A2(n3321), .A3(\inq_ary[0][21] ), 
        .A4(n3315), .Y(n1931) );
  NOR4X1_RVT U2123 ( .A1(n1934), .A2(n1933), .A3(n1932), .A4(n1931), .Y(n1935)
         );
  NAND2X0_RVT U2124 ( .A1(n1936), .A2(n1935), .Y(N282) );
  AO22X1_RVT U2125 ( .A1(\inq_ary[14][22] ), .A2(n3325), .A3(\inq_ary[10][22] ), .A4(n3326), .Y(n1940) );
  AO22X1_RVT U2126 ( .A1(\inq_ary[13][22] ), .A2(n3323), .A3(\inq_ary[7][22] ), 
        .A4(n3322), .Y(n1939) );
  AO22X1_RVT U2127 ( .A1(\inq_ary[12][22] ), .A2(n3303), .A3(\inq_ary[1][22] ), 
        .A4(n3324), .Y(n1938) );
  AO22X1_RVT U2128 ( .A1(\inq_ary[5][22] ), .A2(n3298), .A3(\inq_ary[3][22] ), 
        .A4(n3310), .Y(n1937) );
  NOR4X1_RVT U2129 ( .A1(n1940), .A2(n1939), .A3(n1938), .A4(n1937), .Y(n1946)
         );
  AO22X1_RVT U2130 ( .A1(\inq_ary[8][22] ), .A2(n3313), .A3(\inq_ary[15][22] ), 
        .A4(n3312), .Y(n1944) );
  AO22X1_RVT U2131 ( .A1(\inq_ary[0][22] ), .A2(n3315), .A3(\inq_ary[6][22] ), 
        .A4(n3311), .Y(n1943) );
  AO22X1_RVT U2132 ( .A1(\inq_ary[2][22] ), .A2(n3271), .A3(\inq_ary[9][22] ), 
        .A4(n3314), .Y(n1942) );
  AO22X1_RVT U2133 ( .A1(\inq_ary[4][22] ), .A2(n3321), .A3(\inq_ary[11][22] ), 
        .A4(n3316), .Y(n1941) );
  NOR4X1_RVT U2134 ( .A1(n1944), .A2(n1943), .A3(n1942), .A4(n1941), .Y(n1945)
         );
  NAND2X0_RVT U2135 ( .A1(n1946), .A2(n1945), .Y(N283) );
  AO22X1_RVT U2136 ( .A1(\inq_ary[4][23] ), .A2(n3321), .A3(\inq_ary[9][23] ), 
        .A4(n3314), .Y(n1950) );
  AO22X1_RVT U2137 ( .A1(\inq_ary[2][23] ), .A2(n3271), .A3(\inq_ary[13][23] ), 
        .A4(n3323), .Y(n1949) );
  AO22X1_RVT U2138 ( .A1(\inq_ary[8][23] ), .A2(n3313), .A3(\inq_ary[6][23] ), 
        .A4(n3311), .Y(n1948) );
  AO22X1_RVT U2139 ( .A1(\inq_ary[14][23] ), .A2(n3325), .A3(\inq_ary[5][23] ), 
        .A4(n3298), .Y(n1947) );
  NOR4X1_RVT U2140 ( .A1(n1950), .A2(n1949), .A3(n1948), .A4(n1947), .Y(n1956)
         );
  AO22X1_RVT U2141 ( .A1(\inq_ary[12][23] ), .A2(n3303), .A3(\inq_ary[7][23] ), 
        .A4(n3322), .Y(n1954) );
  AO22X1_RVT U2142 ( .A1(\inq_ary[11][23] ), .A2(n3316), .A3(\inq_ary[0][23] ), 
        .A4(n3315), .Y(n1953) );
  AO22X1_RVT U2143 ( .A1(\inq_ary[1][23] ), .A2(n3324), .A3(\inq_ary[10][23] ), 
        .A4(n3326), .Y(n1952) );
  AO22X1_RVT U2144 ( .A1(\inq_ary[3][23] ), .A2(n3310), .A3(\inq_ary[15][23] ), 
        .A4(n3312), .Y(n1951) );
  NOR4X1_RVT U2145 ( .A1(n1954), .A2(n1953), .A3(n1952), .A4(n1951), .Y(n1955)
         );
  NAND2X0_RVT U2146 ( .A1(n1956), .A2(n1955), .Y(N284) );
  AO22X1_RVT U2147 ( .A1(\inq_ary[14][24] ), .A2(n3325), .A3(\inq_ary[9][24] ), 
        .A4(n3314), .Y(n1960) );
  AO22X1_RVT U2148 ( .A1(\inq_ary[12][24] ), .A2(n3303), .A3(\inq_ary[5][24] ), 
        .A4(n3298), .Y(n1959) );
  AO22X1_RVT U2149 ( .A1(\inq_ary[13][24] ), .A2(n3323), .A3(\inq_ary[8][24] ), 
        .A4(n3313), .Y(n1958) );
  AO22X1_RVT U2150 ( .A1(\inq_ary[2][24] ), .A2(n3271), .A3(\inq_ary[1][24] ), 
        .A4(n3324), .Y(n1957) );
  NOR4X1_RVT U2151 ( .A1(n1960), .A2(n1959), .A3(n1958), .A4(n1957), .Y(n1966)
         );
  AO22X1_RVT U2152 ( .A1(\inq_ary[15][24] ), .A2(n3312), .A3(\inq_ary[6][24] ), 
        .A4(n3311), .Y(n1964) );
  AO22X1_RVT U2153 ( .A1(\inq_ary[4][24] ), .A2(n3321), .A3(\inq_ary[7][24] ), 
        .A4(n3322), .Y(n1963) );
  AO22X1_RVT U2154 ( .A1(\inq_ary[11][24] ), .A2(n3316), .A3(\inq_ary[3][24] ), 
        .A4(n3310), .Y(n1962) );
  AO22X1_RVT U2155 ( .A1(\inq_ary[10][24] ), .A2(n3326), .A3(\inq_ary[0][24] ), 
        .A4(n3315), .Y(n1961) );
  NOR4X1_RVT U2156 ( .A1(n1964), .A2(n1963), .A3(n1962), .A4(n1961), .Y(n1965)
         );
  NAND2X0_RVT U2157 ( .A1(n1966), .A2(n1965), .Y(N285) );
  AO22X1_RVT U2158 ( .A1(\inq_ary[0][25] ), .A2(n3315), .A3(\inq_ary[8][25] ), 
        .A4(n3313), .Y(n1970) );
  AO22X1_RVT U2159 ( .A1(\inq_ary[12][25] ), .A2(n3303), .A3(\inq_ary[9][25] ), 
        .A4(n3314), .Y(n1969) );
  AO22X1_RVT U2160 ( .A1(\inq_ary[14][25] ), .A2(n3325), .A3(\inq_ary[10][25] ), .A4(n3326), .Y(n1968) );
  AO22X1_RVT U2161 ( .A1(\inq_ary[15][25] ), .A2(n3312), .A3(\inq_ary[3][25] ), 
        .A4(n3310), .Y(n1967) );
  NOR4X1_RVT U2162 ( .A1(n1970), .A2(n1969), .A3(n1968), .A4(n1967), .Y(n1976)
         );
  AO22X1_RVT U2163 ( .A1(\inq_ary[2][25] ), .A2(n3271), .A3(\inq_ary[13][25] ), 
        .A4(n3323), .Y(n1974) );
  AO22X1_RVT U2164 ( .A1(\inq_ary[7][25] ), .A2(n3322), .A3(\inq_ary[4][25] ), 
        .A4(n3321), .Y(n1973) );
  AO22X1_RVT U2165 ( .A1(\inq_ary[11][25] ), .A2(n3316), .A3(\inq_ary[1][25] ), 
        .A4(n3324), .Y(n1972) );
  AO22X1_RVT U2166 ( .A1(\inq_ary[6][25] ), .A2(n3311), .A3(\inq_ary[5][25] ), 
        .A4(n3298), .Y(n1971) );
  NOR4X1_RVT U2167 ( .A1(n1974), .A2(n1973), .A3(n1972), .A4(n1971), .Y(n1975)
         );
  NAND2X0_RVT U2168 ( .A1(n1976), .A2(n1975), .Y(N286) );
  AO22X1_RVT U2169 ( .A1(\inq_ary[0][26] ), .A2(n3315), .A3(\inq_ary[8][26] ), 
        .A4(n3313), .Y(n1980) );
  AO22X1_RVT U2170 ( .A1(\inq_ary[11][26] ), .A2(n3316), .A3(\inq_ary[1][26] ), 
        .A4(n3324), .Y(n1979) );
  AO22X1_RVT U2171 ( .A1(\inq_ary[14][26] ), .A2(n3325), .A3(\inq_ary[5][26] ), 
        .A4(n3298), .Y(n1978) );
  AO22X1_RVT U2172 ( .A1(\inq_ary[3][26] ), .A2(n3310), .A3(\inq_ary[6][26] ), 
        .A4(n3311), .Y(n1977) );
  NOR4X1_RVT U2173 ( .A1(n1980), .A2(n1979), .A3(n1978), .A4(n1977), .Y(n1986)
         );
  AO22X1_RVT U2174 ( .A1(\inq_ary[13][26] ), .A2(n3323), .A3(\inq_ary[2][26] ), 
        .A4(n3271), .Y(n1984) );
  AO22X1_RVT U2175 ( .A1(\inq_ary[15][26] ), .A2(n3312), .A3(\inq_ary[10][26] ), .A4(n3326), .Y(n1983) );
  AO22X1_RVT U2176 ( .A1(\inq_ary[7][26] ), .A2(n3322), .A3(\inq_ary[4][26] ), 
        .A4(n3321), .Y(n1982) );
  AO22X1_RVT U2177 ( .A1(\inq_ary[12][26] ), .A2(n3303), .A3(\inq_ary[9][26] ), 
        .A4(n3314), .Y(n1981) );
  NOR4X1_RVT U2178 ( .A1(n1984), .A2(n1983), .A3(n1982), .A4(n1981), .Y(n1985)
         );
  NAND2X0_RVT U2179 ( .A1(n1986), .A2(n1985), .Y(N287) );
  AO22X1_RVT U2180 ( .A1(\inq_ary[6][27] ), .A2(n3311), .A3(\inq_ary[5][27] ), 
        .A4(n3298), .Y(n1990) );
  AO22X1_RVT U2181 ( .A1(\inq_ary[2][27] ), .A2(n3271), .A3(\inq_ary[9][27] ), 
        .A4(n3314), .Y(n1989) );
  AO22X1_RVT U2182 ( .A1(\inq_ary[3][27] ), .A2(n3310), .A3(\inq_ary[7][27] ), 
        .A4(n3322), .Y(n1988) );
  AO22X1_RVT U2183 ( .A1(\inq_ary[11][27] ), .A2(n3316), .A3(\inq_ary[0][27] ), 
        .A4(n3315), .Y(n1987) );
  NOR4X1_RVT U2184 ( .A1(n1990), .A2(n1989), .A3(n1988), .A4(n1987), .Y(n1996)
         );
  AO22X1_RVT U2185 ( .A1(\inq_ary[12][27] ), .A2(n3303), .A3(\inq_ary[1][27] ), 
        .A4(n3324), .Y(n1994) );
  AO22X1_RVT U2186 ( .A1(\inq_ary[15][27] ), .A2(n3312), .A3(\inq_ary[4][27] ), 
        .A4(n3321), .Y(n1993) );
  AO22X1_RVT U2187 ( .A1(\inq_ary[10][27] ), .A2(n3326), .A3(\inq_ary[13][27] ), .A4(n3323), .Y(n1992) );
  AO22X1_RVT U2188 ( .A1(\inq_ary[14][27] ), .A2(n3325), .A3(\inq_ary[8][27] ), 
        .A4(n3313), .Y(n1991) );
  NOR4X1_RVT U2189 ( .A1(n1994), .A2(n1993), .A3(n1992), .A4(n1991), .Y(n1995)
         );
  NAND2X0_RVT U2190 ( .A1(n1996), .A2(n1995), .Y(N288) );
  AO22X1_RVT U2191 ( .A1(\inq_ary[8][28] ), .A2(n3313), .A3(\inq_ary[2][28] ), 
        .A4(n3271), .Y(n2000) );
  AO22X1_RVT U2192 ( .A1(\inq_ary[6][28] ), .A2(n3311), .A3(\inq_ary[14][28] ), 
        .A4(n3325), .Y(n1999) );
  AO22X1_RVT U2193 ( .A1(\inq_ary[7][28] ), .A2(n3322), .A3(\inq_ary[5][28] ), 
        .A4(n3298), .Y(n1998) );
  AO22X1_RVT U2194 ( .A1(\inq_ary[12][28] ), .A2(n3303), .A3(\inq_ary[0][28] ), 
        .A4(n3315), .Y(n1997) );
  NOR4X1_RVT U2195 ( .A1(n2000), .A2(n1999), .A3(n1998), .A4(n1997), .Y(n2006)
         );
  AO22X1_RVT U2196 ( .A1(\inq_ary[1][28] ), .A2(n3324), .A3(\inq_ary[4][28] ), 
        .A4(n3321), .Y(n2004) );
  AO22X1_RVT U2197 ( .A1(\inq_ary[3][28] ), .A2(n3310), .A3(\inq_ary[10][28] ), 
        .A4(n3326), .Y(n2003) );
  AO22X1_RVT U2198 ( .A1(\inq_ary[11][28] ), .A2(n3316), .A3(\inq_ary[9][28] ), 
        .A4(n3314), .Y(n2002) );
  AO22X1_RVT U2199 ( .A1(\inq_ary[13][28] ), .A2(n3323), .A3(\inq_ary[15][28] ), .A4(n3312), .Y(n2001) );
  NOR4X1_RVT U2200 ( .A1(n2004), .A2(n2003), .A3(n2002), .A4(n2001), .Y(n2005)
         );
  NAND2X0_RVT U2201 ( .A1(n2006), .A2(n2005), .Y(N289) );
  AO22X1_RVT U2202 ( .A1(\inq_ary[14][29] ), .A2(n3325), .A3(\inq_ary[8][29] ), 
        .A4(n3313), .Y(n2010) );
  AO22X1_RVT U2203 ( .A1(\inq_ary[11][29] ), .A2(n3316), .A3(\inq_ary[6][29] ), 
        .A4(n3311), .Y(n2009) );
  AO22X1_RVT U2204 ( .A1(\inq_ary[4][29] ), .A2(n3321), .A3(\inq_ary[13][29] ), 
        .A4(n3323), .Y(n2008) );
  AO22X1_RVT U2205 ( .A1(\inq_ary[0][29] ), .A2(n3315), .A3(\inq_ary[1][29] ), 
        .A4(n3324), .Y(n2007) );
  NOR4X1_RVT U2206 ( .A1(n2010), .A2(n2009), .A3(n2008), .A4(n2007), .Y(n2016)
         );
  AO22X1_RVT U2207 ( .A1(\inq_ary[12][29] ), .A2(n3303), .A3(\inq_ary[15][29] ), .A4(n3312), .Y(n2014) );
  AO22X1_RVT U2208 ( .A1(\inq_ary[9][29] ), .A2(n3314), .A3(\inq_ary[3][29] ), 
        .A4(n3310), .Y(n2013) );
  AO22X1_RVT U2209 ( .A1(\inq_ary[7][29] ), .A2(n3322), .A3(\inq_ary[2][29] ), 
        .A4(n3271), .Y(n2012) );
  AO22X1_RVT U2210 ( .A1(\inq_ary[5][29] ), .A2(n3298), .A3(\inq_ary[10][29] ), 
        .A4(n3326), .Y(n2011) );
  NOR4X1_RVT U2211 ( .A1(n2014), .A2(n2013), .A3(n2012), .A4(n2011), .Y(n2015)
         );
  NAND2X0_RVT U2212 ( .A1(n2016), .A2(n2015), .Y(N290) );
  AO22X1_RVT U2213 ( .A1(\inq_ary[9][30] ), .A2(n3314), .A3(\inq_ary[1][30] ), 
        .A4(n3324), .Y(n2020) );
  AO22X1_RVT U2214 ( .A1(\inq_ary[5][30] ), .A2(n3298), .A3(\inq_ary[0][30] ), 
        .A4(n3315), .Y(n2019) );
  AO22X1_RVT U2215 ( .A1(\inq_ary[4][30] ), .A2(n3321), .A3(\inq_ary[14][30] ), 
        .A4(n3325), .Y(n2018) );
  AO22X1_RVT U2216 ( .A1(\inq_ary[3][30] ), .A2(n3310), .A3(\inq_ary[13][30] ), 
        .A4(n3323), .Y(n2017) );
  NOR4X1_RVT U2217 ( .A1(n2020), .A2(n2019), .A3(n2018), .A4(n2017), .Y(n2026)
         );
  AO22X1_RVT U2218 ( .A1(\inq_ary[10][30] ), .A2(n3326), .A3(\inq_ary[11][30] ), .A4(n3316), .Y(n2024) );
  AO22X1_RVT U2219 ( .A1(\inq_ary[8][30] ), .A2(n3313), .A3(\inq_ary[2][30] ), 
        .A4(n3271), .Y(n2023) );
  AO22X1_RVT U2220 ( .A1(\inq_ary[7][30] ), .A2(n3322), .A3(\inq_ary[15][30] ), 
        .A4(n3312), .Y(n2022) );
  AO22X1_RVT U2221 ( .A1(\inq_ary[12][30] ), .A2(n3303), .A3(\inq_ary[6][30] ), 
        .A4(n3311), .Y(n2021) );
  NOR4X1_RVT U2222 ( .A1(n2024), .A2(n2023), .A3(n2022), .A4(n2021), .Y(n2025)
         );
  NAND2X0_RVT U2223 ( .A1(n2026), .A2(n2025), .Y(N291) );
  AO22X1_RVT U2224 ( .A1(\inq_ary[3][31] ), .A2(n3310), .A3(\inq_ary[8][31] ), 
        .A4(n3313), .Y(n2030) );
  AO22X1_RVT U2225 ( .A1(\inq_ary[12][31] ), .A2(n3303), .A3(\inq_ary[1][31] ), 
        .A4(n3324), .Y(n2029) );
  AO22X1_RVT U2226 ( .A1(\inq_ary[14][31] ), .A2(n3325), .A3(\inq_ary[4][31] ), 
        .A4(n3321), .Y(n2028) );
  AO22X1_RVT U2227 ( .A1(\inq_ary[7][31] ), .A2(n3322), .A3(\inq_ary[11][31] ), 
        .A4(n3316), .Y(n2027) );
  NOR4X1_RVT U2228 ( .A1(n2030), .A2(n2029), .A3(n2028), .A4(n2027), .Y(n2036)
         );
  AO22X1_RVT U2229 ( .A1(\inq_ary[2][31] ), .A2(n3271), .A3(\inq_ary[15][31] ), 
        .A4(n3312), .Y(n2034) );
  AO22X1_RVT U2230 ( .A1(\inq_ary[10][31] ), .A2(n3326), .A3(\inq_ary[13][31] ), .A4(n3323), .Y(n2033) );
  AO22X1_RVT U2231 ( .A1(\inq_ary[0][31] ), .A2(n3315), .A3(\inq_ary[5][31] ), 
        .A4(n3298), .Y(n2032) );
  AO22X1_RVT U2232 ( .A1(\inq_ary[9][31] ), .A2(n3314), .A3(\inq_ary[6][31] ), 
        .A4(n3311), .Y(n2031) );
  NOR4X1_RVT U2233 ( .A1(n2034), .A2(n2033), .A3(n2032), .A4(n2031), .Y(n2035)
         );
  NAND2X0_RVT U2234 ( .A1(n2036), .A2(n2035), .Y(N292) );
  AO22X1_RVT U2235 ( .A1(\inq_ary[9][32] ), .A2(n3314), .A3(\inq_ary[12][32] ), 
        .A4(n3303), .Y(n2040) );
  AO22X1_RVT U2236 ( .A1(\inq_ary[14][32] ), .A2(n3325), .A3(\inq_ary[7][32] ), 
        .A4(n3322), .Y(n2039) );
  AO22X1_RVT U2237 ( .A1(\inq_ary[1][32] ), .A2(n3324), .A3(\inq_ary[13][32] ), 
        .A4(n3323), .Y(n2038) );
  AO22X1_RVT U2238 ( .A1(\inq_ary[0][32] ), .A2(n3315), .A3(\inq_ary[5][32] ), 
        .A4(n3298), .Y(n2037) );
  NOR4X1_RVT U2239 ( .A1(n2040), .A2(n2039), .A3(n2038), .A4(n2037), .Y(n2046)
         );
  AO22X1_RVT U2240 ( .A1(\inq_ary[3][32] ), .A2(n3310), .A3(\inq_ary[4][32] ), 
        .A4(n3321), .Y(n2044) );
  AO22X1_RVT U2241 ( .A1(\inq_ary[10][32] ), .A2(n3326), .A3(\inq_ary[8][32] ), 
        .A4(n3313), .Y(n2043) );
  AO22X1_RVT U2242 ( .A1(\inq_ary[11][32] ), .A2(n3316), .A3(\inq_ary[6][32] ), 
        .A4(n3311), .Y(n2042) );
  AO22X1_RVT U2243 ( .A1(\inq_ary[15][32] ), .A2(n3312), .A3(\inq_ary[2][32] ), 
        .A4(n3271), .Y(n2041) );
  NOR4X1_RVT U2244 ( .A1(n2044), .A2(n2043), .A3(n2042), .A4(n2041), .Y(n2045)
         );
  NAND2X0_RVT U2245 ( .A1(n2046), .A2(n2045), .Y(N293) );
  AO22X1_RVT U2246 ( .A1(\inq_ary[1][33] ), .A2(n3324), .A3(\inq_ary[4][33] ), 
        .A4(n3321), .Y(n2050) );
  AO22X1_RVT U2247 ( .A1(\inq_ary[12][33] ), .A2(n3303), .A3(\inq_ary[11][33] ), .A4(n3316), .Y(n2049) );
  AO22X1_RVT U2248 ( .A1(\inq_ary[9][33] ), .A2(n3314), .A3(\inq_ary[6][33] ), 
        .A4(n3311), .Y(n2048) );
  AO22X1_RVT U2249 ( .A1(\inq_ary[8][33] ), .A2(n3313), .A3(\inq_ary[14][33] ), 
        .A4(n3325), .Y(n2047) );
  NOR4X1_RVT U2250 ( .A1(n2050), .A2(n2049), .A3(n2048), .A4(n2047), .Y(n2056)
         );
  AO22X1_RVT U2251 ( .A1(\inq_ary[2][33] ), .A2(n3271), .A3(\inq_ary[3][33] ), 
        .A4(n3310), .Y(n2054) );
  AO22X1_RVT U2252 ( .A1(\inq_ary[5][33] ), .A2(n3298), .A3(\inq_ary[7][33] ), 
        .A4(n3322), .Y(n2053) );
  AO22X1_RVT U2253 ( .A1(\inq_ary[0][33] ), .A2(n3315), .A3(\inq_ary[10][33] ), 
        .A4(n3326), .Y(n2052) );
  AO22X1_RVT U2254 ( .A1(\inq_ary[13][33] ), .A2(n3323), .A3(\inq_ary[15][33] ), .A4(n3312), .Y(n2051) );
  NOR4X1_RVT U2255 ( .A1(n2054), .A2(n2053), .A3(n2052), .A4(n2051), .Y(n2055)
         );
  NAND2X0_RVT U2256 ( .A1(n2056), .A2(n2055), .Y(N294) );
  AO22X1_RVT U2257 ( .A1(\inq_ary[3][34] ), .A2(n3310), .A3(\inq_ary[12][34] ), 
        .A4(n3303), .Y(n2060) );
  AO22X1_RVT U2258 ( .A1(\inq_ary[7][34] ), .A2(n3322), .A3(\inq_ary[15][34] ), 
        .A4(n3312), .Y(n2059) );
  AO22X1_RVT U2259 ( .A1(\inq_ary[11][34] ), .A2(n3316), .A3(\inq_ary[1][34] ), 
        .A4(n3324), .Y(n2058) );
  AO22X1_RVT U2260 ( .A1(\inq_ary[0][34] ), .A2(n3315), .A3(\inq_ary[5][34] ), 
        .A4(n3298), .Y(n2057) );
  NOR4X1_RVT U2261 ( .A1(n2060), .A2(n2059), .A3(n2058), .A4(n2057), .Y(n2066)
         );
  AO22X1_RVT U2262 ( .A1(\inq_ary[9][34] ), .A2(n3314), .A3(\inq_ary[13][34] ), 
        .A4(n3323), .Y(n2064) );
  AO22X1_RVT U2263 ( .A1(\inq_ary[8][34] ), .A2(n3313), .A3(\inq_ary[10][34] ), 
        .A4(n3326), .Y(n2063) );
  AO22X1_RVT U2264 ( .A1(\inq_ary[14][34] ), .A2(n3325), .A3(\inq_ary[6][34] ), 
        .A4(n3311), .Y(n2062) );
  AO22X1_RVT U2265 ( .A1(\inq_ary[2][34] ), .A2(n3271), .A3(\inq_ary[4][34] ), 
        .A4(n3321), .Y(n2061) );
  NOR4X1_RVT U2266 ( .A1(n2064), .A2(n2063), .A3(n2062), .A4(n2061), .Y(n2065)
         );
  NAND2X0_RVT U2267 ( .A1(n2066), .A2(n2065), .Y(N295) );
  AO22X1_RVT U2268 ( .A1(\inq_ary[10][35] ), .A2(n3326), .A3(\inq_ary[8][35] ), 
        .A4(n3313), .Y(n2070) );
  AO22X1_RVT U2269 ( .A1(\inq_ary[9][35] ), .A2(n3314), .A3(\inq_ary[14][35] ), 
        .A4(n3325), .Y(n2069) );
  AO22X1_RVT U2270 ( .A1(\inq_ary[13][35] ), .A2(n3323), .A3(\inq_ary[6][35] ), 
        .A4(n3311), .Y(n2068) );
  AO22X1_RVT U2271 ( .A1(\inq_ary[2][35] ), .A2(n3271), .A3(\inq_ary[5][35] ), 
        .A4(n3298), .Y(n2067) );
  NOR4X1_RVT U2272 ( .A1(n2070), .A2(n2069), .A3(n2068), .A4(n2067), .Y(n2076)
         );
  AO22X1_RVT U2273 ( .A1(\inq_ary[4][35] ), .A2(n3321), .A3(\inq_ary[0][35] ), 
        .A4(n3315), .Y(n2074) );
  AO22X1_RVT U2274 ( .A1(\inq_ary[12][35] ), .A2(n3303), .A3(\inq_ary[15][35] ), .A4(n3312), .Y(n2073) );
  AO22X1_RVT U2275 ( .A1(\inq_ary[3][35] ), .A2(n3310), .A3(\inq_ary[7][35] ), 
        .A4(n3322), .Y(n2072) );
  AO22X1_RVT U2276 ( .A1(\inq_ary[11][35] ), .A2(n3316), .A3(\inq_ary[1][35] ), 
        .A4(n3324), .Y(n2071) );
  NOR4X1_RVT U2277 ( .A1(n2074), .A2(n2073), .A3(n2072), .A4(n2071), .Y(n2075)
         );
  NAND2X0_RVT U2278 ( .A1(n2076), .A2(n2075), .Y(N296) );
  AO22X1_RVT U2279 ( .A1(\inq_ary[12][36] ), .A2(n3303), .A3(\inq_ary[6][36] ), 
        .A4(n3311), .Y(n2080) );
  AO22X1_RVT U2280 ( .A1(\inq_ary[2][36] ), .A2(n3271), .A3(\inq_ary[5][36] ), 
        .A4(n3298), .Y(n2079) );
  AO22X1_RVT U2281 ( .A1(\inq_ary[0][36] ), .A2(n3315), .A3(\inq_ary[15][36] ), 
        .A4(n3312), .Y(n2078) );
  AO22X1_RVT U2282 ( .A1(\inq_ary[1][36] ), .A2(n3324), .A3(\inq_ary[10][36] ), 
        .A4(n3326), .Y(n2077) );
  NOR4X1_RVT U2283 ( .A1(n2080), .A2(n2079), .A3(n2078), .A4(n2077), .Y(n2086)
         );
  AO22X1_RVT U2284 ( .A1(\inq_ary[11][36] ), .A2(n3316), .A3(\inq_ary[4][36] ), 
        .A4(n3321), .Y(n2084) );
  AO22X1_RVT U2285 ( .A1(\inq_ary[8][36] ), .A2(n3313), .A3(\inq_ary[9][36] ), 
        .A4(n3314), .Y(n2083) );
  AO22X1_RVT U2286 ( .A1(\inq_ary[7][36] ), .A2(n3322), .A3(\inq_ary[14][36] ), 
        .A4(n3325), .Y(n2082) );
  AO22X1_RVT U2287 ( .A1(\inq_ary[13][36] ), .A2(n3323), .A3(\inq_ary[3][36] ), 
        .A4(n3310), .Y(n2081) );
  NOR4X1_RVT U2288 ( .A1(n2084), .A2(n2083), .A3(n2082), .A4(n2081), .Y(n2085)
         );
  NAND2X0_RVT U2289 ( .A1(n2086), .A2(n2085), .Y(N297) );
  AO22X1_RVT U2290 ( .A1(\inq_ary[14][37] ), .A2(n3325), .A3(\inq_ary[8][37] ), 
        .A4(n3313), .Y(n2090) );
  AO22X1_RVT U2291 ( .A1(\inq_ary[4][37] ), .A2(n3321), .A3(\inq_ary[11][37] ), 
        .A4(n3316), .Y(n2089) );
  AO22X1_RVT U2292 ( .A1(\inq_ary[2][37] ), .A2(n3271), .A3(\inq_ary[15][37] ), 
        .A4(n3312), .Y(n2088) );
  AO22X1_RVT U2293 ( .A1(\inq_ary[12][37] ), .A2(n3303), .A3(\inq_ary[9][37] ), 
        .A4(n3314), .Y(n2087) );
  NOR4X1_RVT U2294 ( .A1(n2090), .A2(n2089), .A3(n2088), .A4(n2087), .Y(n2096)
         );
  AO22X1_RVT U2295 ( .A1(\inq_ary[13][37] ), .A2(n3323), .A3(\inq_ary[10][37] ), .A4(n3326), .Y(n2094) );
  AO22X1_RVT U2296 ( .A1(\inq_ary[6][37] ), .A2(n3311), .A3(\inq_ary[0][37] ), 
        .A4(n3315), .Y(n2093) );
  AO22X1_RVT U2297 ( .A1(\inq_ary[3][37] ), .A2(n3310), .A3(\inq_ary[5][37] ), 
        .A4(n3298), .Y(n2092) );
  AO22X1_RVT U2298 ( .A1(\inq_ary[1][37] ), .A2(n3324), .A3(\inq_ary[7][37] ), 
        .A4(n3322), .Y(n2091) );
  NOR4X1_RVT U2299 ( .A1(n2094), .A2(n2093), .A3(n2092), .A4(n2091), .Y(n2095)
         );
  NAND2X0_RVT U2300 ( .A1(n2096), .A2(n2095), .Y(N298) );
  AO22X1_RVT U2301 ( .A1(\inq_ary[13][38] ), .A2(n3323), .A3(\inq_ary[5][38] ), 
        .A4(n3298), .Y(n2100) );
  AO22X1_RVT U2302 ( .A1(\inq_ary[10][38] ), .A2(n3326), .A3(\inq_ary[8][38] ), 
        .A4(n3313), .Y(n2099) );
  AO22X1_RVT U2303 ( .A1(\inq_ary[11][38] ), .A2(n3316), .A3(\inq_ary[1][38] ), 
        .A4(n3324), .Y(n2098) );
  AO22X1_RVT U2304 ( .A1(\inq_ary[4][38] ), .A2(n3321), .A3(\inq_ary[2][38] ), 
        .A4(n3271), .Y(n2097) );
  NOR4X1_RVT U2305 ( .A1(n2100), .A2(n2099), .A3(n2098), .A4(n2097), .Y(n2106)
         );
  AO22X1_RVT U2306 ( .A1(\inq_ary[14][38] ), .A2(n3325), .A3(\inq_ary[12][38] ), .A4(n3303), .Y(n2104) );
  AO22X1_RVT U2307 ( .A1(\inq_ary[6][38] ), .A2(n3311), .A3(\inq_ary[0][38] ), 
        .A4(n3315), .Y(n2103) );
  AO22X1_RVT U2308 ( .A1(\inq_ary[9][38] ), .A2(n3314), .A3(\inq_ary[3][38] ), 
        .A4(n3310), .Y(n2102) );
  AO22X1_RVT U2309 ( .A1(\inq_ary[15][38] ), .A2(n3312), .A3(\inq_ary[7][38] ), 
        .A4(n3322), .Y(n2101) );
  NOR4X1_RVT U2310 ( .A1(n2104), .A2(n2103), .A3(n2102), .A4(n2101), .Y(n2105)
         );
  NAND2X0_RVT U2311 ( .A1(n2106), .A2(n2105), .Y(N299) );
  AO22X1_RVT U2312 ( .A1(\inq_ary[2][39] ), .A2(n3271), .A3(\inq_ary[10][39] ), 
        .A4(n3326), .Y(n2110) );
  AO22X1_RVT U2313 ( .A1(\inq_ary[1][39] ), .A2(n3324), .A3(\inq_ary[8][39] ), 
        .A4(n3313), .Y(n2109) );
  AO22X1_RVT U2314 ( .A1(\inq_ary[14][39] ), .A2(n3325), .A3(\inq_ary[12][39] ), .A4(n3303), .Y(n2108) );
  AO22X1_RVT U2315 ( .A1(\inq_ary[5][39] ), .A2(n3298), .A3(\inq_ary[7][39] ), 
        .A4(n3322), .Y(n2107) );
  NOR4X1_RVT U2316 ( .A1(n2110), .A2(n2109), .A3(n2108), .A4(n2107), .Y(n2116)
         );
  AO22X1_RVT U2317 ( .A1(\inq_ary[3][39] ), .A2(n3310), .A3(\inq_ary[13][39] ), 
        .A4(n3323), .Y(n2114) );
  AO22X1_RVT U2318 ( .A1(\inq_ary[4][39] ), .A2(n3321), .A3(\inq_ary[9][39] ), 
        .A4(n3314), .Y(n2113) );
  AO22X1_RVT U2319 ( .A1(\inq_ary[15][39] ), .A2(n3312), .A3(\inq_ary[6][39] ), 
        .A4(n3311), .Y(n2112) );
  AO22X1_RVT U2320 ( .A1(\inq_ary[11][39] ), .A2(n3316), .A3(\inq_ary[0][39] ), 
        .A4(n3315), .Y(n2111) );
  NOR4X1_RVT U2321 ( .A1(n2114), .A2(n2113), .A3(n2112), .A4(n2111), .Y(n2115)
         );
  NAND2X0_RVT U2322 ( .A1(n2116), .A2(n2115), .Y(N300) );
  AO22X1_RVT U2323 ( .A1(\inq_ary[13][40] ), .A2(n3323), .A3(\inq_ary[10][40] ), .A4(n3326), .Y(n2120) );
  AO22X1_RVT U2324 ( .A1(\inq_ary[6][40] ), .A2(n3311), .A3(\inq_ary[5][40] ), 
        .A4(n3298), .Y(n2119) );
  AO22X1_RVT U2325 ( .A1(\inq_ary[11][40] ), .A2(n3316), .A3(\inq_ary[1][40] ), 
        .A4(n3324), .Y(n2118) );
  AO22X1_RVT U2326 ( .A1(\inq_ary[4][40] ), .A2(n3321), .A3(\inq_ary[15][40] ), 
        .A4(n3312), .Y(n2117) );
  NOR4X1_RVT U2327 ( .A1(n2120), .A2(n2119), .A3(n2118), .A4(n2117), .Y(n2126)
         );
  AO22X1_RVT U2328 ( .A1(\inq_ary[7][40] ), .A2(n3322), .A3(\inq_ary[3][40] ), 
        .A4(n3310), .Y(n2124) );
  AO22X1_RVT U2329 ( .A1(\inq_ary[14][40] ), .A2(n3325), .A3(\inq_ary[0][40] ), 
        .A4(n3315), .Y(n2123) );
  AO22X1_RVT U2330 ( .A1(\inq_ary[12][40] ), .A2(n3303), .A3(\inq_ary[2][40] ), 
        .A4(n3271), .Y(n2122) );
  AO22X1_RVT U2331 ( .A1(\inq_ary[8][40] ), .A2(n3313), .A3(\inq_ary[9][40] ), 
        .A4(n3314), .Y(n2121) );
  NOR4X1_RVT U2332 ( .A1(n2124), .A2(n2123), .A3(n2122), .A4(n2121), .Y(n2125)
         );
  NAND2X0_RVT U2333 ( .A1(n2126), .A2(n2125), .Y(N301) );
  AO22X1_RVT U2334 ( .A1(\inq_ary[2][41] ), .A2(n3271), .A3(\inq_ary[8][41] ), 
        .A4(n3313), .Y(n2130) );
  AO22X1_RVT U2335 ( .A1(\inq_ary[13][41] ), .A2(n3323), .A3(\inq_ary[14][41] ), .A4(n3325), .Y(n2129) );
  AO22X1_RVT U2336 ( .A1(\inq_ary[7][41] ), .A2(n3322), .A3(\inq_ary[12][41] ), 
        .A4(n3303), .Y(n2128) );
  AO22X1_RVT U2337 ( .A1(\inq_ary[11][41] ), .A2(n3316), .A3(\inq_ary[1][41] ), 
        .A4(n3324), .Y(n2127) );
  NOR4X1_RVT U2338 ( .A1(n2130), .A2(n2129), .A3(n2128), .A4(n2127), .Y(n2136)
         );
  AO22X1_RVT U2339 ( .A1(\inq_ary[10][41] ), .A2(n3326), .A3(\inq_ary[9][41] ), 
        .A4(n3314), .Y(n2134) );
  AO22X1_RVT U2340 ( .A1(\inq_ary[6][41] ), .A2(n3311), .A3(\inq_ary[5][41] ), 
        .A4(n3298), .Y(n2133) );
  AO22X1_RVT U2341 ( .A1(\inq_ary[0][41] ), .A2(n3315), .A3(\inq_ary[15][41] ), 
        .A4(n3312), .Y(n2132) );
  AO22X1_RVT U2342 ( .A1(\inq_ary[3][41] ), .A2(n3310), .A3(\inq_ary[4][41] ), 
        .A4(n3321), .Y(n2131) );
  NOR4X1_RVT U2343 ( .A1(n2134), .A2(n2133), .A3(n2132), .A4(n2131), .Y(n2135)
         );
  NAND2X0_RVT U2344 ( .A1(n2136), .A2(n2135), .Y(N302) );
  AO22X1_RVT U2345 ( .A1(\inq_ary[11][42] ), .A2(n3316), .A3(\inq_ary[0][42] ), 
        .A4(n3315), .Y(n2140) );
  AO22X1_RVT U2346 ( .A1(\inq_ary[10][42] ), .A2(n3326), .A3(\inq_ary[13][42] ), .A4(n3323), .Y(n2139) );
  AO22X1_RVT U2347 ( .A1(\inq_ary[9][42] ), .A2(n3314), .A3(\inq_ary[3][42] ), 
        .A4(n3310), .Y(n2138) );
  AO22X1_RVT U2348 ( .A1(\inq_ary[4][42] ), .A2(n3321), .A3(\inq_ary[5][42] ), 
        .A4(n3298), .Y(n2137) );
  NOR4X1_RVT U2349 ( .A1(n2140), .A2(n2139), .A3(n2138), .A4(n2137), .Y(n2146)
         );
  AO22X1_RVT U2350 ( .A1(\inq_ary[15][42] ), .A2(n3312), .A3(\inq_ary[1][42] ), 
        .A4(n3324), .Y(n2144) );
  AO22X1_RVT U2351 ( .A1(\inq_ary[6][42] ), .A2(n3311), .A3(\inq_ary[7][42] ), 
        .A4(n3322), .Y(n2143) );
  AO22X1_RVT U2352 ( .A1(\inq_ary[2][42] ), .A2(n3271), .A3(\inq_ary[8][42] ), 
        .A4(n3313), .Y(n2142) );
  AO22X1_RVT U2353 ( .A1(\inq_ary[12][42] ), .A2(n3303), .A3(\inq_ary[14][42] ), .A4(n3325), .Y(n2141) );
  NOR4X1_RVT U2354 ( .A1(n2144), .A2(n2143), .A3(n2142), .A4(n2141), .Y(n2145)
         );
  NAND2X0_RVT U2355 ( .A1(n2146), .A2(n2145), .Y(N303) );
  AO22X1_RVT U2356 ( .A1(\inq_ary[8][43] ), .A2(n3313), .A3(\inq_ary[14][43] ), 
        .A4(n3325), .Y(n2150) );
  AO22X1_RVT U2357 ( .A1(\inq_ary[10][43] ), .A2(n3326), .A3(\inq_ary[13][43] ), .A4(n3323), .Y(n2149) );
  AO22X1_RVT U2358 ( .A1(\inq_ary[2][43] ), .A2(n3271), .A3(\inq_ary[6][43] ), 
        .A4(n3311), .Y(n2148) );
  AO22X1_RVT U2359 ( .A1(\inq_ary[1][43] ), .A2(n3324), .A3(\inq_ary[5][43] ), 
        .A4(n3298), .Y(n2147) );
  NOR4X1_RVT U2360 ( .A1(n2150), .A2(n2149), .A3(n2148), .A4(n2147), .Y(n2156)
         );
  AO22X1_RVT U2361 ( .A1(\inq_ary[15][43] ), .A2(n3312), .A3(\inq_ary[12][43] ), .A4(n3303), .Y(n2154) );
  AO22X1_RVT U2362 ( .A1(\inq_ary[9][43] ), .A2(n3314), .A3(\inq_ary[7][43] ), 
        .A4(n3322), .Y(n2153) );
  AO22X1_RVT U2363 ( .A1(\inq_ary[0][43] ), .A2(n3315), .A3(\inq_ary[4][43] ), 
        .A4(n3321), .Y(n2152) );
  AO22X1_RVT U2364 ( .A1(\inq_ary[3][43] ), .A2(n3310), .A3(\inq_ary[11][43] ), 
        .A4(n3316), .Y(n2151) );
  NOR4X1_RVT U2365 ( .A1(n2154), .A2(n2153), .A3(n2152), .A4(n2151), .Y(n2155)
         );
  NAND2X0_RVT U2366 ( .A1(n2156), .A2(n2155), .Y(N304) );
  AO22X1_RVT U2367 ( .A1(\inq_ary[12][44] ), .A2(n3303), .A3(\inq_ary[8][44] ), 
        .A4(n3313), .Y(n2160) );
  AO22X1_RVT U2368 ( .A1(\inq_ary[1][44] ), .A2(n3324), .A3(\inq_ary[14][44] ), 
        .A4(n3325), .Y(n2159) );
  AO22X1_RVT U2369 ( .A1(\inq_ary[10][44] ), .A2(n3326), .A3(\inq_ary[5][44] ), 
        .A4(n3298), .Y(n2158) );
  AO22X1_RVT U2370 ( .A1(\inq_ary[11][44] ), .A2(n3316), .A3(\inq_ary[3][44] ), 
        .A4(n3310), .Y(n2157) );
  NOR4X1_RVT U2371 ( .A1(n2160), .A2(n2159), .A3(n2158), .A4(n2157), .Y(n2166)
         );
  AO22X1_RVT U2372 ( .A1(\inq_ary[4][44] ), .A2(n3321), .A3(\inq_ary[13][44] ), 
        .A4(n3323), .Y(n2164) );
  AO22X1_RVT U2373 ( .A1(\inq_ary[6][44] ), .A2(n3311), .A3(\inq_ary[7][44] ), 
        .A4(n3322), .Y(n2163) );
  AO22X1_RVT U2374 ( .A1(\inq_ary[9][44] ), .A2(n3314), .A3(\inq_ary[0][44] ), 
        .A4(n3315), .Y(n2162) );
  AO22X1_RVT U2375 ( .A1(\inq_ary[15][44] ), .A2(n3312), .A3(\inq_ary[2][44] ), 
        .A4(n3271), .Y(n2161) );
  NOR4X1_RVT U2376 ( .A1(n2164), .A2(n2163), .A3(n2162), .A4(n2161), .Y(n2165)
         );
  NAND2X0_RVT U2377 ( .A1(n2166), .A2(n2165), .Y(N305) );
  AO22X1_RVT U2378 ( .A1(\inq_ary[5][45] ), .A2(n3298), .A3(\inq_ary[2][45] ), 
        .A4(n3271), .Y(n2170) );
  AO22X1_RVT U2379 ( .A1(\inq_ary[12][45] ), .A2(n3303), .A3(\inq_ary[3][45] ), 
        .A4(n3310), .Y(n2169) );
  AO22X1_RVT U2380 ( .A1(\inq_ary[8][45] ), .A2(n3313), .A3(\inq_ary[14][45] ), 
        .A4(n3325), .Y(n2168) );
  AO22X1_RVT U2381 ( .A1(\inq_ary[7][45] ), .A2(n3322), .A3(\inq_ary[1][45] ), 
        .A4(n3324), .Y(n2167) );
  NOR4X1_RVT U2382 ( .A1(n2170), .A2(n2169), .A3(n2168), .A4(n2167), .Y(n2176)
         );
  AO22X1_RVT U2383 ( .A1(\inq_ary[4][45] ), .A2(n3321), .A3(\inq_ary[11][45] ), 
        .A4(n3316), .Y(n2174) );
  AO22X1_RVT U2384 ( .A1(\inq_ary[0][45] ), .A2(n3315), .A3(\inq_ary[9][45] ), 
        .A4(n3314), .Y(n2173) );
  AO22X1_RVT U2385 ( .A1(\inq_ary[10][45] ), .A2(n3326), .A3(\inq_ary[13][45] ), .A4(n3323), .Y(n2172) );
  AO22X1_RVT U2386 ( .A1(\inq_ary[6][45] ), .A2(n3311), .A3(\inq_ary[15][45] ), 
        .A4(n3312), .Y(n2171) );
  NOR4X1_RVT U2387 ( .A1(n2174), .A2(n2173), .A3(n2172), .A4(n2171), .Y(n2175)
         );
  NAND2X0_RVT U2388 ( .A1(n2176), .A2(n2175), .Y(N306) );
  AO22X1_RVT U2389 ( .A1(\inq_ary[4][46] ), .A2(n3321), .A3(\inq_ary[15][46] ), 
        .A4(n3312), .Y(n2180) );
  AO22X1_RVT U2390 ( .A1(\inq_ary[14][46] ), .A2(n3325), .A3(\inq_ary[0][46] ), 
        .A4(n3315), .Y(n2179) );
  AO22X1_RVT U2391 ( .A1(\inq_ary[2][46] ), .A2(n3271), .A3(\inq_ary[5][46] ), 
        .A4(n3298), .Y(n2178) );
  AO22X1_RVT U2392 ( .A1(\inq_ary[10][46] ), .A2(n3326), .A3(\inq_ary[9][46] ), 
        .A4(n3314), .Y(n2177) );
  NOR4X1_RVT U2393 ( .A1(n2180), .A2(n2179), .A3(n2178), .A4(n2177), .Y(n2186)
         );
  AO22X1_RVT U2394 ( .A1(\inq_ary[6][46] ), .A2(n3311), .A3(\inq_ary[3][46] ), 
        .A4(n3310), .Y(n2184) );
  AO22X1_RVT U2395 ( .A1(\inq_ary[13][46] ), .A2(n3323), .A3(\inq_ary[7][46] ), 
        .A4(n3322), .Y(n2183) );
  AO22X1_RVT U2396 ( .A1(\inq_ary[8][46] ), .A2(n3313), .A3(\inq_ary[12][46] ), 
        .A4(n3303), .Y(n2182) );
  AO22X1_RVT U2397 ( .A1(\inq_ary[1][46] ), .A2(n3324), .A3(\inq_ary[11][46] ), 
        .A4(n3316), .Y(n2181) );
  NOR4X1_RVT U2398 ( .A1(n2184), .A2(n2183), .A3(n2182), .A4(n2181), .Y(n2185)
         );
  NAND2X0_RVT U2399 ( .A1(n2186), .A2(n2185), .Y(N307) );
  AO22X1_RVT U2400 ( .A1(\inq_ary[2][47] ), .A2(n3271), .A3(\inq_ary[10][47] ), 
        .A4(n3326), .Y(n2190) );
  AO22X1_RVT U2401 ( .A1(\inq_ary[15][47] ), .A2(n3312), .A3(\inq_ary[5][47] ), 
        .A4(n3298), .Y(n2189) );
  AO22X1_RVT U2402 ( .A1(\inq_ary[0][47] ), .A2(n3315), .A3(\inq_ary[6][47] ), 
        .A4(n3311), .Y(n2188) );
  AO22X1_RVT U2403 ( .A1(\inq_ary[4][47] ), .A2(n3321), .A3(\inq_ary[11][47] ), 
        .A4(n3316), .Y(n2187) );
  NOR4X1_RVT U2404 ( .A1(n2190), .A2(n2189), .A3(n2188), .A4(n2187), .Y(n2196)
         );
  AO22X1_RVT U2405 ( .A1(\inq_ary[8][47] ), .A2(n3313), .A3(\inq_ary[9][47] ), 
        .A4(n3314), .Y(n2194) );
  AO22X1_RVT U2406 ( .A1(\inq_ary[13][47] ), .A2(n3323), .A3(\inq_ary[3][47] ), 
        .A4(n3310), .Y(n2193) );
  AO22X1_RVT U2407 ( .A1(\inq_ary[1][47] ), .A2(n3324), .A3(\inq_ary[7][47] ), 
        .A4(n3322), .Y(n2192) );
  AO22X1_RVT U2408 ( .A1(\inq_ary[14][47] ), .A2(n3325), .A3(\inq_ary[12][47] ), .A4(n3303), .Y(n2191) );
  NOR4X1_RVT U2409 ( .A1(n2194), .A2(n2193), .A3(n2192), .A4(n2191), .Y(n2195)
         );
  NAND2X0_RVT U2410 ( .A1(n2196), .A2(n2195), .Y(N308) );
  AO22X1_RVT U2411 ( .A1(\inq_ary[0][48] ), .A2(n3315), .A3(\inq_ary[5][48] ), 
        .A4(n3298), .Y(n2200) );
  AO22X1_RVT U2412 ( .A1(\inq_ary[12][48] ), .A2(n3303), .A3(\inq_ary[13][48] ), .A4(n3323), .Y(n2199) );
  AO22X1_RVT U2413 ( .A1(\inq_ary[8][48] ), .A2(n3313), .A3(\inq_ary[14][48] ), 
        .A4(n3325), .Y(n2198) );
  AO22X1_RVT U2414 ( .A1(\inq_ary[11][48] ), .A2(n3316), .A3(\inq_ary[3][48] ), 
        .A4(n3310), .Y(n2197) );
  NOR4X1_RVT U2415 ( .A1(n2200), .A2(n2199), .A3(n2198), .A4(n2197), .Y(n2206)
         );
  AO22X1_RVT U2416 ( .A1(\inq_ary[7][48] ), .A2(n3322), .A3(\inq_ary[9][48] ), 
        .A4(n3314), .Y(n2204) );
  AO22X1_RVT U2417 ( .A1(\inq_ary[15][48] ), .A2(n3312), .A3(\inq_ary[4][48] ), 
        .A4(n3321), .Y(n2203) );
  AO22X1_RVT U2418 ( .A1(\inq_ary[1][48] ), .A2(n3324), .A3(\inq_ary[2][48] ), 
        .A4(n3271), .Y(n2202) );
  AO22X1_RVT U2419 ( .A1(\inq_ary[10][48] ), .A2(n3326), .A3(\inq_ary[6][48] ), 
        .A4(n3311), .Y(n2201) );
  NOR4X1_RVT U2420 ( .A1(n2204), .A2(n2203), .A3(n2202), .A4(n2201), .Y(n2205)
         );
  NAND2X0_RVT U2421 ( .A1(n2206), .A2(n2205), .Y(N309) );
  AO22X1_RVT U2422 ( .A1(\inq_ary[3][49] ), .A2(n3310), .A3(\inq_ary[11][49] ), 
        .A4(n3316), .Y(n2210) );
  AO22X1_RVT U2423 ( .A1(\inq_ary[10][49] ), .A2(n3326), .A3(\inq_ary[14][49] ), .A4(n3325), .Y(n2209) );
  AO22X1_RVT U2424 ( .A1(\inq_ary[2][49] ), .A2(n3271), .A3(\inq_ary[15][49] ), 
        .A4(n3312), .Y(n2208) );
  AO22X1_RVT U2425 ( .A1(\inq_ary[4][49] ), .A2(n3321), .A3(\inq_ary[7][49] ), 
        .A4(n3322), .Y(n2207) );
  NOR4X1_RVT U2426 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), .Y(n2216)
         );
  AO22X1_RVT U2427 ( .A1(\inq_ary[9][49] ), .A2(n3314), .A3(\inq_ary[1][49] ), 
        .A4(n3324), .Y(n2214) );
  AO22X1_RVT U2428 ( .A1(\inq_ary[13][49] ), .A2(n3323), .A3(\inq_ary[0][49] ), 
        .A4(n3315), .Y(n2213) );
  AO22X1_RVT U2429 ( .A1(\inq_ary[5][49] ), .A2(n3298), .A3(\inq_ary[12][49] ), 
        .A4(n3303), .Y(n2212) );
  AO22X1_RVT U2430 ( .A1(\inq_ary[6][49] ), .A2(n3311), .A3(\inq_ary[8][49] ), 
        .A4(n3313), .Y(n2211) );
  NOR4X1_RVT U2431 ( .A1(n2214), .A2(n2213), .A3(n2212), .A4(n2211), .Y(n2215)
         );
  NAND2X0_RVT U2432 ( .A1(n2216), .A2(n2215), .Y(N310) );
  AO22X1_RVT U2433 ( .A1(\inq_ary[4][50] ), .A2(n3321), .A3(\inq_ary[15][50] ), 
        .A4(n3312), .Y(n2220) );
  AO22X1_RVT U2434 ( .A1(\inq_ary[10][50] ), .A2(n3326), .A3(\inq_ary[6][50] ), 
        .A4(n3311), .Y(n2219) );
  AO22X1_RVT U2435 ( .A1(\inq_ary[14][50] ), .A2(n3325), .A3(\inq_ary[0][50] ), 
        .A4(n3315), .Y(n2218) );
  AO22X1_RVT U2436 ( .A1(\inq_ary[5][50] ), .A2(n3298), .A3(\inq_ary[7][50] ), 
        .A4(n3322), .Y(n2217) );
  NOR4X1_RVT U2437 ( .A1(n2220), .A2(n2219), .A3(n2218), .A4(n2217), .Y(n2226)
         );
  AO22X1_RVT U2438 ( .A1(\inq_ary[3][50] ), .A2(n3310), .A3(\inq_ary[11][50] ), 
        .A4(n3316), .Y(n2224) );
  AO22X1_RVT U2439 ( .A1(\inq_ary[2][50] ), .A2(n3271), .A3(\inq_ary[9][50] ), 
        .A4(n3314), .Y(n2223) );
  AO22X1_RVT U2440 ( .A1(\inq_ary[13][50] ), .A2(n3323), .A3(\inq_ary[8][50] ), 
        .A4(n3313), .Y(n2222) );
  AO22X1_RVT U2441 ( .A1(\inq_ary[1][50] ), .A2(n3324), .A3(\inq_ary[12][50] ), 
        .A4(n3303), .Y(n2221) );
  NOR4X1_RVT U2442 ( .A1(n2224), .A2(n2223), .A3(n2222), .A4(n2221), .Y(n2225)
         );
  NAND2X0_RVT U2443 ( .A1(n2226), .A2(n2225), .Y(N311) );
  AO22X1_RVT U2444 ( .A1(\inq_ary[5][51] ), .A2(n3298), .A3(\inq_ary[10][51] ), 
        .A4(n3326), .Y(n2230) );
  AO22X1_RVT U2445 ( .A1(\inq_ary[11][51] ), .A2(n3316), .A3(\inq_ary[3][51] ), 
        .A4(n3310), .Y(n2229) );
  AO22X1_RVT U2446 ( .A1(\inq_ary[13][51] ), .A2(n3323), .A3(\inq_ary[0][51] ), 
        .A4(n3315), .Y(n2228) );
  AO22X1_RVT U2447 ( .A1(\inq_ary[12][51] ), .A2(n3303), .A3(\inq_ary[9][51] ), 
        .A4(n3314), .Y(n2227) );
  NOR4X1_RVT U2448 ( .A1(n2230), .A2(n2229), .A3(n2228), .A4(n2227), .Y(n2236)
         );
  AO22X1_RVT U2449 ( .A1(\inq_ary[2][51] ), .A2(n3271), .A3(\inq_ary[1][51] ), 
        .A4(n3324), .Y(n2234) );
  AO22X1_RVT U2450 ( .A1(\inq_ary[15][51] ), .A2(n3312), .A3(\inq_ary[6][51] ), 
        .A4(n3311), .Y(n2233) );
  AO22X1_RVT U2451 ( .A1(\inq_ary[7][51] ), .A2(n3322), .A3(\inq_ary[4][51] ), 
        .A4(n3321), .Y(n2232) );
  AO22X1_RVT U2452 ( .A1(\inq_ary[8][51] ), .A2(n3313), .A3(\inq_ary[14][51] ), 
        .A4(n3325), .Y(n2231) );
  NOR4X1_RVT U2453 ( .A1(n2234), .A2(n2233), .A3(n2232), .A4(n2231), .Y(n2235)
         );
  NAND2X0_RVT U2454 ( .A1(n2236), .A2(n2235), .Y(N312) );
  AO22X1_RVT U2455 ( .A1(\inq_ary[15][52] ), .A2(n3312), .A3(\inq_ary[2][52] ), 
        .A4(n3271), .Y(n2240) );
  AO22X1_RVT U2456 ( .A1(\inq_ary[13][52] ), .A2(n3323), .A3(\inq_ary[0][52] ), 
        .A4(n3315), .Y(n2239) );
  AO22X1_RVT U2457 ( .A1(\inq_ary[5][52] ), .A2(n3298), .A3(\inq_ary[8][52] ), 
        .A4(n3313), .Y(n2238) );
  AO22X1_RVT U2458 ( .A1(\inq_ary[7][52] ), .A2(n3322), .A3(\inq_ary[9][52] ), 
        .A4(n3314), .Y(n2237) );
  NOR4X1_RVT U2459 ( .A1(n2240), .A2(n2239), .A3(n2238), .A4(n2237), .Y(n2246)
         );
  AO22X1_RVT U2460 ( .A1(\inq_ary[10][52] ), .A2(n3326), .A3(\inq_ary[12][52] ), .A4(n3303), .Y(n2244) );
  AO22X1_RVT U2461 ( .A1(\inq_ary[11][52] ), .A2(n3316), .A3(\inq_ary[3][52] ), 
        .A4(n3310), .Y(n2243) );
  AO22X1_RVT U2462 ( .A1(\inq_ary[14][52] ), .A2(n3325), .A3(\inq_ary[1][52] ), 
        .A4(n3324), .Y(n2242) );
  AO22X1_RVT U2463 ( .A1(\inq_ary[4][52] ), .A2(n3321), .A3(\inq_ary[6][52] ), 
        .A4(n3311), .Y(n2241) );
  NOR4X1_RVT U2464 ( .A1(n2244), .A2(n2243), .A3(n2242), .A4(n2241), .Y(n2245)
         );
  NAND2X0_RVT U2465 ( .A1(n2246), .A2(n2245), .Y(N313) );
  AO22X1_RVT U2466 ( .A1(\inq_ary[9][53] ), .A2(n3314), .A3(\inq_ary[4][53] ), 
        .A4(n3321), .Y(n2250) );
  AO22X1_RVT U2467 ( .A1(\inq_ary[13][53] ), .A2(n3323), .A3(\inq_ary[3][53] ), 
        .A4(n3310), .Y(n2249) );
  AO22X1_RVT U2468 ( .A1(\inq_ary[1][53] ), .A2(n3324), .A3(\inq_ary[15][53] ), 
        .A4(n3312), .Y(n2248) );
  AO22X1_RVT U2469 ( .A1(\inq_ary[6][53] ), .A2(n3311), .A3(\inq_ary[8][53] ), 
        .A4(n3313), .Y(n2247) );
  NOR4X1_RVT U2470 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .Y(n2256)
         );
  AO22X1_RVT U2471 ( .A1(\inq_ary[14][53] ), .A2(n3325), .A3(\inq_ary[5][53] ), 
        .A4(n3298), .Y(n2254) );
  AO22X1_RVT U2472 ( .A1(\inq_ary[0][53] ), .A2(n3315), .A3(\inq_ary[12][53] ), 
        .A4(n3303), .Y(n2253) );
  AO22X1_RVT U2473 ( .A1(\inq_ary[2][53] ), .A2(n3271), .A3(\inq_ary[7][53] ), 
        .A4(n3322), .Y(n2252) );
  AO22X1_RVT U2474 ( .A1(\inq_ary[10][53] ), .A2(n3326), .A3(\inq_ary[11][53] ), .A4(n3316), .Y(n2251) );
  NOR4X1_RVT U2475 ( .A1(n2254), .A2(n2253), .A3(n2252), .A4(n2251), .Y(n2255)
         );
  NAND2X0_RVT U2476 ( .A1(n2256), .A2(n2255), .Y(N314) );
  AO22X1_RVT U2477 ( .A1(\inq_ary[13][54] ), .A2(n3323), .A3(\inq_ary[8][54] ), 
        .A4(n3313), .Y(n2260) );
  AO22X1_RVT U2478 ( .A1(\inq_ary[14][54] ), .A2(n3325), .A3(\inq_ary[2][54] ), 
        .A4(n3271), .Y(n2259) );
  AO22X1_RVT U2479 ( .A1(\inq_ary[10][54] ), .A2(n3326), .A3(\inq_ary[9][54] ), 
        .A4(n3314), .Y(n2258) );
  AO22X1_RVT U2480 ( .A1(\inq_ary[7][54] ), .A2(n3322), .A3(\inq_ary[11][54] ), 
        .A4(n3316), .Y(n2257) );
  NOR4X1_RVT U2481 ( .A1(n2260), .A2(n2259), .A3(n2258), .A4(n2257), .Y(n2266)
         );
  AO22X1_RVT U2482 ( .A1(\inq_ary[0][54] ), .A2(n3315), .A3(\inq_ary[12][54] ), 
        .A4(n3303), .Y(n2264) );
  AO22X1_RVT U2483 ( .A1(\inq_ary[6][54] ), .A2(n3311), .A3(\inq_ary[3][54] ), 
        .A4(n3310), .Y(n2263) );
  AO22X1_RVT U2484 ( .A1(\inq_ary[1][54] ), .A2(n3324), .A3(\inq_ary[5][54] ), 
        .A4(n3298), .Y(n2262) );
  AO22X1_RVT U2485 ( .A1(\inq_ary[4][54] ), .A2(n3321), .A3(\inq_ary[15][54] ), 
        .A4(n3312), .Y(n2261) );
  NOR4X1_RVT U2486 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2261), .Y(n2265)
         );
  NAND2X0_RVT U2487 ( .A1(n2266), .A2(n2265), .Y(N315) );
  AO22X1_RVT U2488 ( .A1(\inq_ary[11][55] ), .A2(n3316), .A3(\inq_ary[9][55] ), 
        .A4(n3314), .Y(n2270) );
  AO22X1_RVT U2489 ( .A1(\inq_ary[0][55] ), .A2(n3315), .A3(\inq_ary[1][55] ), 
        .A4(n3324), .Y(n2269) );
  AO22X1_RVT U2490 ( .A1(\inq_ary[15][55] ), .A2(n3312), .A3(\inq_ary[12][55] ), .A4(n3303), .Y(n2268) );
  AO22X1_RVT U2491 ( .A1(\inq_ary[3][55] ), .A2(n3310), .A3(\inq_ary[4][55] ), 
        .A4(n3321), .Y(n2267) );
  NOR4X1_RVT U2492 ( .A1(n2270), .A2(n2269), .A3(n2268), .A4(n2267), .Y(n2276)
         );
  AO22X1_RVT U2493 ( .A1(\inq_ary[14][55] ), .A2(n3325), .A3(\inq_ary[13][55] ), .A4(n3323), .Y(n2274) );
  AO22X1_RVT U2494 ( .A1(\inq_ary[6][55] ), .A2(n3311), .A3(\inq_ary[7][55] ), 
        .A4(n3322), .Y(n2273) );
  AO22X1_RVT U2495 ( .A1(\inq_ary[10][55] ), .A2(n3326), .A3(\inq_ary[8][55] ), 
        .A4(n3313), .Y(n2272) );
  AO22X1_RVT U2496 ( .A1(\inq_ary[5][55] ), .A2(n3298), .A3(\inq_ary[2][55] ), 
        .A4(n3271), .Y(n2271) );
  NOR4X1_RVT U2497 ( .A1(n2274), .A2(n2273), .A3(n2272), .A4(n2271), .Y(n2275)
         );
  NAND2X0_RVT U2498 ( .A1(n2276), .A2(n2275), .Y(N316) );
  AO22X1_RVT U2499 ( .A1(\inq_ary[12][56] ), .A2(n3303), .A3(\inq_ary[0][56] ), 
        .A4(n3315), .Y(n2280) );
  AO22X1_RVT U2500 ( .A1(\inq_ary[6][56] ), .A2(n3311), .A3(\inq_ary[5][56] ), 
        .A4(n3298), .Y(n2279) );
  AO22X1_RVT U2501 ( .A1(\inq_ary[1][56] ), .A2(n3324), .A3(\inq_ary[11][56] ), 
        .A4(n3316), .Y(n2278) );
  AO22X1_RVT U2502 ( .A1(\inq_ary[4][56] ), .A2(n3321), .A3(\inq_ary[10][56] ), 
        .A4(n3326), .Y(n2277) );
  NOR4X1_RVT U2503 ( .A1(n2280), .A2(n2279), .A3(n2278), .A4(n2277), .Y(n2286)
         );
  AO22X1_RVT U2504 ( .A1(\inq_ary[9][56] ), .A2(n3314), .A3(\inq_ary[7][56] ), 
        .A4(n3322), .Y(n2284) );
  AO22X1_RVT U2505 ( .A1(\inq_ary[13][56] ), .A2(n3323), .A3(\inq_ary[14][56] ), .A4(n3325), .Y(n2283) );
  AO22X1_RVT U2506 ( .A1(\inq_ary[8][56] ), .A2(n3313), .A3(\inq_ary[2][56] ), 
        .A4(n3271), .Y(n2282) );
  AO22X1_RVT U2507 ( .A1(\inq_ary[15][56] ), .A2(n3312), .A3(\inq_ary[3][56] ), 
        .A4(n3310), .Y(n2281) );
  NOR4X1_RVT U2508 ( .A1(n2284), .A2(n2283), .A3(n2282), .A4(n2281), .Y(n2285)
         );
  NAND2X0_RVT U2509 ( .A1(n2286), .A2(n2285), .Y(N317) );
  AO22X1_RVT U2510 ( .A1(\inq_ary[12][57] ), .A2(n3303), .A3(\inq_ary[2][57] ), 
        .A4(n3271), .Y(n2290) );
  AO22X1_RVT U2511 ( .A1(\inq_ary[4][57] ), .A2(n3321), .A3(\inq_ary[5][57] ), 
        .A4(n3298), .Y(n2289) );
  AO22X1_RVT U2512 ( .A1(\inq_ary[15][57] ), .A2(n3312), .A3(\inq_ary[13][57] ), .A4(n3323), .Y(n2288) );
  AO22X1_RVT U2513 ( .A1(\inq_ary[3][57] ), .A2(n3310), .A3(\inq_ary[7][57] ), 
        .A4(n3322), .Y(n2287) );
  NOR4X1_RVT U2514 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), .Y(n2296)
         );
  AO22X1_RVT U2515 ( .A1(\inq_ary[10][57] ), .A2(n3326), .A3(\inq_ary[0][57] ), 
        .A4(n3315), .Y(n2294) );
  AO22X1_RVT U2516 ( .A1(\inq_ary[9][57] ), .A2(n3314), .A3(\inq_ary[11][57] ), 
        .A4(n3316), .Y(n2293) );
  AO22X1_RVT U2517 ( .A1(\inq_ary[8][57] ), .A2(n3313), .A3(\inq_ary[6][57] ), 
        .A4(n3311), .Y(n2292) );
  AO22X1_RVT U2518 ( .A1(\inq_ary[1][57] ), .A2(n3324), .A3(\inq_ary[14][57] ), 
        .A4(n3325), .Y(n2291) );
  NOR4X1_RVT U2519 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), .Y(n2295)
         );
  NAND2X0_RVT U2520 ( .A1(n2296), .A2(n2295), .Y(N318) );
  AO22X1_RVT U2521 ( .A1(\inq_ary[8][58] ), .A2(n3313), .A3(\inq_ary[4][58] ), 
        .A4(n3321), .Y(n2300) );
  AO22X1_RVT U2522 ( .A1(\inq_ary[15][58] ), .A2(n3312), .A3(\inq_ary[7][58] ), 
        .A4(n3322), .Y(n2299) );
  AO22X1_RVT U2523 ( .A1(\inq_ary[14][58] ), .A2(n3325), .A3(\inq_ary[12][58] ), .A4(n3303), .Y(n2298) );
  AO22X1_RVT U2524 ( .A1(\inq_ary[6][58] ), .A2(n3311), .A3(\inq_ary[2][58] ), 
        .A4(n3271), .Y(n2297) );
  NOR4X1_RVT U2525 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .Y(n2306)
         );
  AO22X1_RVT U2526 ( .A1(\inq_ary[13][58] ), .A2(n3323), .A3(\inq_ary[1][58] ), 
        .A4(n3324), .Y(n2304) );
  AO22X1_RVT U2527 ( .A1(\inq_ary[10][58] ), .A2(n3326), .A3(\inq_ary[11][58] ), .A4(n3316), .Y(n2303) );
  AO22X1_RVT U2528 ( .A1(\inq_ary[5][58] ), .A2(n3298), .A3(\inq_ary[3][58] ), 
        .A4(n3310), .Y(n2302) );
  AO22X1_RVT U2529 ( .A1(\inq_ary[9][58] ), .A2(n3314), .A3(\inq_ary[0][58] ), 
        .A4(n3315), .Y(n2301) );
  NOR4X1_RVT U2530 ( .A1(n2304), .A2(n2303), .A3(n2302), .A4(n2301), .Y(n2305)
         );
  NAND2X0_RVT U2531 ( .A1(n2306), .A2(n2305), .Y(N319) );
  AO22X1_RVT U2532 ( .A1(\inq_ary[1][59] ), .A2(n3324), .A3(\inq_ary[0][59] ), 
        .A4(n3315), .Y(n2310) );
  AO22X1_RVT U2533 ( .A1(\inq_ary[11][59] ), .A2(n3316), .A3(\inq_ary[9][59] ), 
        .A4(n3314), .Y(n2309) );
  AO22X1_RVT U2534 ( .A1(\inq_ary[8][59] ), .A2(n3313), .A3(\inq_ary[12][59] ), 
        .A4(n3303), .Y(n2308) );
  AO22X1_RVT U2535 ( .A1(\inq_ary[5][59] ), .A2(n3298), .A3(\inq_ary[10][59] ), 
        .A4(n3326), .Y(n2307) );
  NOR4X1_RVT U2536 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), .Y(n2316)
         );
  AO22X1_RVT U2537 ( .A1(\inq_ary[4][59] ), .A2(n3321), .A3(\inq_ary[3][59] ), 
        .A4(n3310), .Y(n2314) );
  AO22X1_RVT U2538 ( .A1(\inq_ary[2][59] ), .A2(n3271), .A3(\inq_ary[7][59] ), 
        .A4(n3322), .Y(n2313) );
  AO22X1_RVT U2539 ( .A1(\inq_ary[14][59] ), .A2(n3325), .A3(\inq_ary[13][59] ), .A4(n3323), .Y(n2312) );
  AO22X1_RVT U2540 ( .A1(\inq_ary[6][59] ), .A2(n3311), .A3(\inq_ary[15][59] ), 
        .A4(n3312), .Y(n2311) );
  NOR4X1_RVT U2541 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .Y(n2315)
         );
  NAND2X0_RVT U2542 ( .A1(n2316), .A2(n2315), .Y(N320) );
  AO22X1_RVT U2543 ( .A1(\inq_ary[12][60] ), .A2(n3303), .A3(\inq_ary[11][60] ), .A4(n3316), .Y(n2320) );
  AO22X1_RVT U2544 ( .A1(\inq_ary[9][60] ), .A2(n3314), .A3(\inq_ary[5][60] ), 
        .A4(n3298), .Y(n2319) );
  AO22X1_RVT U2545 ( .A1(\inq_ary[15][60] ), .A2(n3312), .A3(\inq_ary[14][60] ), .A4(n3325), .Y(n2318) );
  AO22X1_RVT U2546 ( .A1(\inq_ary[13][60] ), .A2(n3323), .A3(\inq_ary[4][60] ), 
        .A4(n3321), .Y(n2317) );
  NOR4X1_RVT U2547 ( .A1(n2320), .A2(n2319), .A3(n2318), .A4(n2317), .Y(n2326)
         );
  AO22X1_RVT U2548 ( .A1(\inq_ary[3][60] ), .A2(n3310), .A3(\inq_ary[0][60] ), 
        .A4(n3315), .Y(n2324) );
  AO22X1_RVT U2549 ( .A1(\inq_ary[1][60] ), .A2(n3324), .A3(\inq_ary[10][60] ), 
        .A4(n3326), .Y(n2323) );
  AO22X1_RVT U2550 ( .A1(\inq_ary[8][60] ), .A2(n3313), .A3(\inq_ary[7][60] ), 
        .A4(n3322), .Y(n2322) );
  AO22X1_RVT U2551 ( .A1(\inq_ary[6][60] ), .A2(n3311), .A3(\inq_ary[2][60] ), 
        .A4(n3271), .Y(n2321) );
  NOR4X1_RVT U2552 ( .A1(n2324), .A2(n2323), .A3(n2322), .A4(n2321), .Y(n2325)
         );
  NAND2X0_RVT U2553 ( .A1(n2326), .A2(n2325), .Y(N321) );
  AO22X1_RVT U2554 ( .A1(\inq_ary[11][61] ), .A2(n3316), .A3(\inq_ary[15][61] ), .A4(n3312), .Y(n2330) );
  AO22X1_RVT U2555 ( .A1(\inq_ary[9][61] ), .A2(n3314), .A3(\inq_ary[14][61] ), 
        .A4(n3325), .Y(n2329) );
  AO22X1_RVT U2556 ( .A1(\inq_ary[3][61] ), .A2(n3310), .A3(\inq_ary[13][61] ), 
        .A4(n3323), .Y(n2328) );
  AO22X1_RVT U2557 ( .A1(\inq_ary[4][61] ), .A2(n3321), .A3(\inq_ary[1][61] ), 
        .A4(n3324), .Y(n2327) );
  NOR4X1_RVT U2558 ( .A1(n2330), .A2(n2329), .A3(n2328), .A4(n2327), .Y(n2336)
         );
  AO22X1_RVT U2559 ( .A1(\inq_ary[6][61] ), .A2(n3311), .A3(\inq_ary[2][61] ), 
        .A4(n3271), .Y(n2334) );
  AO22X1_RVT U2560 ( .A1(\inq_ary[8][61] ), .A2(n3313), .A3(\inq_ary[7][61] ), 
        .A4(n3322), .Y(n2333) );
  AO22X1_RVT U2561 ( .A1(\inq_ary[12][61] ), .A2(n3303), .A3(\inq_ary[0][61] ), 
        .A4(n3315), .Y(n2332) );
  AO22X1_RVT U2562 ( .A1(\inq_ary[10][61] ), .A2(n3326), .A3(\inq_ary[5][61] ), 
        .A4(n3298), .Y(n2331) );
  NOR4X1_RVT U2563 ( .A1(n2334), .A2(n2333), .A3(n2332), .A4(n2331), .Y(n2335)
         );
  NAND2X0_RVT U2564 ( .A1(n2336), .A2(n2335), .Y(N322) );
  AO22X1_RVT U2565 ( .A1(\inq_ary[14][62] ), .A2(n3325), .A3(\inq_ary[0][62] ), 
        .A4(n3315), .Y(n2340) );
  AO22X1_RVT U2566 ( .A1(\inq_ary[7][62] ), .A2(n3322), .A3(\inq_ary[12][62] ), 
        .A4(n3303), .Y(n2339) );
  AO22X1_RVT U2567 ( .A1(\inq_ary[15][62] ), .A2(n3312), .A3(\inq_ary[6][62] ), 
        .A4(n3311), .Y(n2338) );
  AO22X1_RVT U2568 ( .A1(\inq_ary[2][62] ), .A2(n3271), .A3(\inq_ary[8][62] ), 
        .A4(n3313), .Y(n2337) );
  NOR4X1_RVT U2569 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .Y(n2346)
         );
  AO22X1_RVT U2570 ( .A1(\inq_ary[10][62] ), .A2(n3326), .A3(\inq_ary[13][62] ), .A4(n3323), .Y(n2344) );
  AO22X1_RVT U2571 ( .A1(\inq_ary[4][62] ), .A2(n3321), .A3(\inq_ary[1][62] ), 
        .A4(n3324), .Y(n2343) );
  AO22X1_RVT U2572 ( .A1(\inq_ary[3][62] ), .A2(n3310), .A3(\inq_ary[11][62] ), 
        .A4(n3316), .Y(n2342) );
  AO22X1_RVT U2573 ( .A1(\inq_ary[5][62] ), .A2(n3298), .A3(\inq_ary[9][62] ), 
        .A4(n3314), .Y(n2341) );
  NOR4X1_RVT U2574 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .Y(n2345)
         );
  NAND2X0_RVT U2575 ( .A1(n2346), .A2(n2345), .Y(N323) );
  AO22X1_RVT U2576 ( .A1(\inq_ary[2][63] ), .A2(n3271), .A3(\inq_ary[1][63] ), 
        .A4(n3324), .Y(n2350) );
  AO22X1_RVT U2577 ( .A1(\inq_ary[4][63] ), .A2(n3321), .A3(\inq_ary[15][63] ), 
        .A4(n3312), .Y(n2349) );
  AO22X1_RVT U2578 ( .A1(\inq_ary[13][63] ), .A2(n3323), .A3(\inq_ary[10][63] ), .A4(n3326), .Y(n2348) );
  AO22X1_RVT U2579 ( .A1(\inq_ary[12][63] ), .A2(n3303), .A3(\inq_ary[11][63] ), .A4(n3316), .Y(n2347) );
  NOR4X1_RVT U2580 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .Y(n2356)
         );
  AO22X1_RVT U2581 ( .A1(\inq_ary[3][63] ), .A2(n3310), .A3(\inq_ary[5][63] ), 
        .A4(n3298), .Y(n2354) );
  AO22X1_RVT U2582 ( .A1(\inq_ary[6][63] ), .A2(n3311), .A3(\inq_ary[0][63] ), 
        .A4(n3315), .Y(n2353) );
  AO22X1_RVT U2583 ( .A1(\inq_ary[7][63] ), .A2(n3322), .A3(\inq_ary[8][63] ), 
        .A4(n3313), .Y(n2352) );
  AO22X1_RVT U2584 ( .A1(\inq_ary[14][63] ), .A2(n3325), .A3(\inq_ary[9][63] ), 
        .A4(n3314), .Y(n2351) );
  NOR4X1_RVT U2585 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), .Y(n2355)
         );
  NAND2X0_RVT U2586 ( .A1(n2356), .A2(n2355), .Y(N324) );
  AO22X1_RVT U2587 ( .A1(\inq_ary[0][64] ), .A2(n3315), .A3(\inq_ary[11][64] ), 
        .A4(n3316), .Y(n2360) );
  AO22X1_RVT U2588 ( .A1(\inq_ary[1][64] ), .A2(n3324), .A3(\inq_ary[14][64] ), 
        .A4(n3325), .Y(n2359) );
  AO22X1_RVT U2589 ( .A1(\inq_ary[2][64] ), .A2(n3271), .A3(\inq_ary[9][64] ), 
        .A4(n3314), .Y(n2358) );
  AO22X1_RVT U2590 ( .A1(\inq_ary[4][64] ), .A2(n3321), .A3(\inq_ary[7][64] ), 
        .A4(n3322), .Y(n2357) );
  NOR4X1_RVT U2591 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .Y(n2366)
         );
  AO22X1_RVT U2592 ( .A1(\inq_ary[5][64] ), .A2(n3298), .A3(\inq_ary[10][64] ), 
        .A4(n3326), .Y(n2364) );
  AO22X1_RVT U2593 ( .A1(\inq_ary[13][64] ), .A2(n3323), .A3(\inq_ary[6][64] ), 
        .A4(n3311), .Y(n2363) );
  AO22X1_RVT U2594 ( .A1(\inq_ary[15][64] ), .A2(n3312), .A3(\inq_ary[3][64] ), 
        .A4(n3310), .Y(n2362) );
  AO22X1_RVT U2595 ( .A1(\inq_ary[8][64] ), .A2(n3313), .A3(\inq_ary[12][64] ), 
        .A4(n3303), .Y(n2361) );
  NOR4X1_RVT U2596 ( .A1(n2364), .A2(n2363), .A3(n2362), .A4(n2361), .Y(n2365)
         );
  NAND2X0_RVT U2597 ( .A1(n2366), .A2(n2365), .Y(N325) );
  AO22X1_RVT U2598 ( .A1(\inq_ary[13][65] ), .A2(n3323), .A3(\inq_ary[9][65] ), 
        .A4(n3314), .Y(n2370) );
  AO22X1_RVT U2599 ( .A1(\inq_ary[8][65] ), .A2(n3313), .A3(\inq_ary[4][65] ), 
        .A4(n3321), .Y(n2369) );
  AO22X1_RVT U2600 ( .A1(\inq_ary[3][65] ), .A2(n3310), .A3(\inq_ary[11][65] ), 
        .A4(n3316), .Y(n2368) );
  AO22X1_RVT U2601 ( .A1(\inq_ary[1][65] ), .A2(n3324), .A3(\inq_ary[6][65] ), 
        .A4(n3311), .Y(n2367) );
  NOR4X1_RVT U2602 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .Y(n2376)
         );
  AO22X1_RVT U2603 ( .A1(\inq_ary[10][65] ), .A2(n3326), .A3(\inq_ary[15][65] ), .A4(n3312), .Y(n2374) );
  AO22X1_RVT U2604 ( .A1(\inq_ary[14][65] ), .A2(n3325), .A3(\inq_ary[5][65] ), 
        .A4(n3298), .Y(n2373) );
  AO22X1_RVT U2605 ( .A1(\inq_ary[7][65] ), .A2(n3322), .A3(\inq_ary[0][65] ), 
        .A4(n3315), .Y(n2372) );
  AO22X1_RVT U2606 ( .A1(\inq_ary[2][65] ), .A2(n3271), .A3(\inq_ary[12][65] ), 
        .A4(n3303), .Y(n2371) );
  NOR4X1_RVT U2607 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), .Y(n2375)
         );
  NAND2X0_RVT U2608 ( .A1(n2376), .A2(n2375), .Y(N326) );
  AO22X1_RVT U2609 ( .A1(\inq_ary[6][66] ), .A2(n3311), .A3(\inq_ary[2][66] ), 
        .A4(n3271), .Y(n2380) );
  AO22X1_RVT U2610 ( .A1(\inq_ary[7][66] ), .A2(n3322), .A3(\inq_ary[15][66] ), 
        .A4(n3312), .Y(n2379) );
  AO22X1_RVT U2611 ( .A1(\inq_ary[4][66] ), .A2(n3321), .A3(\inq_ary[3][66] ), 
        .A4(n3310), .Y(n2378) );
  AO22X1_RVT U2612 ( .A1(\inq_ary[8][66] ), .A2(n3313), .A3(\inq_ary[14][66] ), 
        .A4(n3325), .Y(n2377) );
  NOR4X1_RVT U2613 ( .A1(n2380), .A2(n2379), .A3(n2378), .A4(n2377), .Y(n2386)
         );
  AO22X1_RVT U2614 ( .A1(\inq_ary[11][66] ), .A2(n3316), .A3(\inq_ary[5][66] ), 
        .A4(n3298), .Y(n2384) );
  AO22X1_RVT U2615 ( .A1(\inq_ary[10][66] ), .A2(n3326), .A3(\inq_ary[0][66] ), 
        .A4(n3315), .Y(n2383) );
  AO22X1_RVT U2616 ( .A1(\inq_ary[1][66] ), .A2(n3324), .A3(\inq_ary[12][66] ), 
        .A4(n3303), .Y(n2382) );
  AO22X1_RVT U2617 ( .A1(\inq_ary[13][66] ), .A2(n3323), .A3(\inq_ary[9][66] ), 
        .A4(n3314), .Y(n2381) );
  NOR4X1_RVT U2618 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .Y(n2385)
         );
  NAND2X0_RVT U2619 ( .A1(n2386), .A2(n2385), .Y(N327) );
  AO22X1_RVT U2620 ( .A1(\inq_ary[15][67] ), .A2(n3312), .A3(\inq_ary[2][67] ), 
        .A4(n3271), .Y(n2390) );
  AO22X1_RVT U2621 ( .A1(\inq_ary[7][67] ), .A2(n3322), .A3(\inq_ary[4][67] ), 
        .A4(n3321), .Y(n2389) );
  AO22X1_RVT U2622 ( .A1(\inq_ary[14][67] ), .A2(n3325), .A3(\inq_ary[13][67] ), .A4(n3323), .Y(n2388) );
  AO22X1_RVT U2623 ( .A1(\inq_ary[11][67] ), .A2(n3316), .A3(\inq_ary[10][67] ), .A4(n3326), .Y(n2387) );
  NOR4X1_RVT U2624 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .Y(n2396)
         );
  AO22X1_RVT U2625 ( .A1(\inq_ary[6][67] ), .A2(n3311), .A3(\inq_ary[0][67] ), 
        .A4(n3315), .Y(n2394) );
  AO22X1_RVT U2626 ( .A1(\inq_ary[8][67] ), .A2(n3313), .A3(\inq_ary[9][67] ), 
        .A4(n3314), .Y(n2393) );
  AO22X1_RVT U2627 ( .A1(\inq_ary[12][67] ), .A2(n3303), .A3(\inq_ary[1][67] ), 
        .A4(n3324), .Y(n2392) );
  AO22X1_RVT U2628 ( .A1(\inq_ary[3][67] ), .A2(n3310), .A3(\inq_ary[5][67] ), 
        .A4(n3298), .Y(n2391) );
  NOR4X1_RVT U2629 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .Y(n2395)
         );
  NAND2X0_RVT U2630 ( .A1(n2396), .A2(n2395), .Y(N328) );
  AO22X1_RVT U2631 ( .A1(\inq_ary[6][68] ), .A2(n3311), .A3(\inq_ary[8][68] ), 
        .A4(n3313), .Y(n2400) );
  AO22X1_RVT U2632 ( .A1(\inq_ary[3][68] ), .A2(n3310), .A3(\inq_ary[5][68] ), 
        .A4(n3298), .Y(n2399) );
  AO22X1_RVT U2633 ( .A1(\inq_ary[12][68] ), .A2(n3303), .A3(\inq_ary[11][68] ), .A4(n3316), .Y(n2398) );
  AO22X1_RVT U2634 ( .A1(\inq_ary[9][68] ), .A2(n3314), .A3(\inq_ary[15][68] ), 
        .A4(n3312), .Y(n2397) );
  NOR4X1_RVT U2635 ( .A1(n2400), .A2(n2399), .A3(n2398), .A4(n2397), .Y(n2406)
         );
  AO22X1_RVT U2636 ( .A1(\inq_ary[7][68] ), .A2(n3322), .A3(\inq_ary[13][68] ), 
        .A4(n3323), .Y(n2404) );
  AO22X1_RVT U2637 ( .A1(\inq_ary[14][68] ), .A2(n3325), .A3(\inq_ary[2][68] ), 
        .A4(n3271), .Y(n2403) );
  AO22X1_RVT U2638 ( .A1(\inq_ary[10][68] ), .A2(n3326), .A3(\inq_ary[4][68] ), 
        .A4(n3321), .Y(n2402) );
  AO22X1_RVT U2639 ( .A1(\inq_ary[1][68] ), .A2(n3324), .A3(\inq_ary[0][68] ), 
        .A4(n3315), .Y(n2401) );
  NOR4X1_RVT U2640 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .Y(n2405)
         );
  NAND2X0_RVT U2641 ( .A1(n2406), .A2(n2405), .Y(N329) );
  AO22X1_RVT U2642 ( .A1(\inq_ary[5][69] ), .A2(n3298), .A3(\inq_ary[2][69] ), 
        .A4(n3271), .Y(n2410) );
  AO22X1_RVT U2643 ( .A1(\inq_ary[7][69] ), .A2(n3322), .A3(\inq_ary[3][69] ), 
        .A4(n3310), .Y(n2409) );
  AO22X1_RVT U2644 ( .A1(\inq_ary[9][69] ), .A2(n3314), .A3(\inq_ary[14][69] ), 
        .A4(n3325), .Y(n2408) );
  AO22X1_RVT U2645 ( .A1(\inq_ary[0][69] ), .A2(n3315), .A3(\inq_ary[8][69] ), 
        .A4(n3313), .Y(n2407) );
  NOR4X1_RVT U2646 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .Y(n2416)
         );
  AO22X1_RVT U2647 ( .A1(\inq_ary[4][69] ), .A2(n3321), .A3(\inq_ary[6][69] ), 
        .A4(n3311), .Y(n2414) );
  AO22X1_RVT U2648 ( .A1(\inq_ary[12][69] ), .A2(n3303), .A3(\inq_ary[10][69] ), .A4(n3326), .Y(n2413) );
  AO22X1_RVT U2649 ( .A1(\inq_ary[1][69] ), .A2(n3324), .A3(\inq_ary[13][69] ), 
        .A4(n3323), .Y(n2412) );
  AO22X1_RVT U2650 ( .A1(\inq_ary[15][69] ), .A2(n3312), .A3(\inq_ary[11][69] ), .A4(n3316), .Y(n2411) );
  NOR4X1_RVT U2651 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .Y(n2415)
         );
  NAND2X0_RVT U2652 ( .A1(n2416), .A2(n2415), .Y(N330) );
  AO22X1_RVT U2653 ( .A1(\inq_ary[12][70] ), .A2(n3303), .A3(\inq_ary[3][70] ), 
        .A4(n3310), .Y(n2420) );
  AO22X1_RVT U2654 ( .A1(\inq_ary[5][70] ), .A2(n3298), .A3(\inq_ary[0][70] ), 
        .A4(n3315), .Y(n2419) );
  AO22X1_RVT U2655 ( .A1(\inq_ary[1][70] ), .A2(n3324), .A3(\inq_ary[11][70] ), 
        .A4(n3316), .Y(n2418) );
  AO22X1_RVT U2656 ( .A1(\inq_ary[10][70] ), .A2(n3326), .A3(\inq_ary[7][70] ), 
        .A4(n3322), .Y(n2417) );
  NOR4X1_RVT U2657 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .Y(n2426)
         );
  AO22X1_RVT U2658 ( .A1(\inq_ary[4][70] ), .A2(n3321), .A3(\inq_ary[15][70] ), 
        .A4(n3312), .Y(n2424) );
  AO22X1_RVT U2659 ( .A1(\inq_ary[6][70] ), .A2(n3311), .A3(\inq_ary[14][70] ), 
        .A4(n3325), .Y(n2423) );
  AO22X1_RVT U2660 ( .A1(\inq_ary[2][70] ), .A2(n3271), .A3(\inq_ary[8][70] ), 
        .A4(n3313), .Y(n2422) );
  AO22X1_RVT U2661 ( .A1(\inq_ary[13][70] ), .A2(n3323), .A3(\inq_ary[9][70] ), 
        .A4(n3314), .Y(n2421) );
  NOR4X1_RVT U2662 ( .A1(n2424), .A2(n2423), .A3(n2422), .A4(n2421), .Y(n2425)
         );
  NAND2X0_RVT U2663 ( .A1(n2426), .A2(n2425), .Y(N331) );
  AO22X1_RVT U2664 ( .A1(\inq_ary[9][71] ), .A2(n3314), .A3(\inq_ary[10][71] ), 
        .A4(n3326), .Y(n2430) );
  AO22X1_RVT U2665 ( .A1(\inq_ary[8][71] ), .A2(n3313), .A3(\inq_ary[13][71] ), 
        .A4(n3323), .Y(n2429) );
  AO22X1_RVT U2666 ( .A1(\inq_ary[3][71] ), .A2(n3310), .A3(\inq_ary[12][71] ), 
        .A4(n3303), .Y(n2428) );
  AO22X1_RVT U2667 ( .A1(\inq_ary[15][71] ), .A2(n3312), .A3(\inq_ary[5][71] ), 
        .A4(n3298), .Y(n2427) );
  NOR4X1_RVT U2668 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .Y(n2436)
         );
  AO22X1_RVT U2669 ( .A1(\inq_ary[0][71] ), .A2(n3315), .A3(\inq_ary[14][71] ), 
        .A4(n3325), .Y(n2434) );
  AO22X1_RVT U2670 ( .A1(\inq_ary[11][71] ), .A2(n3316), .A3(\inq_ary[2][71] ), 
        .A4(n3271), .Y(n2433) );
  AO22X1_RVT U2671 ( .A1(\inq_ary[4][71] ), .A2(n3321), .A3(\inq_ary[6][71] ), 
        .A4(n3311), .Y(n2432) );
  AO22X1_RVT U2672 ( .A1(\inq_ary[7][71] ), .A2(n3322), .A3(\inq_ary[1][71] ), 
        .A4(n3324), .Y(n2431) );
  NOR4X1_RVT U2673 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .Y(n2435)
         );
  NAND2X0_RVT U2674 ( .A1(n2436), .A2(n2435), .Y(N332) );
  AO22X1_RVT U2675 ( .A1(\inq_ary[11][72] ), .A2(n3316), .A3(\inq_ary[13][72] ), .A4(n3323), .Y(n2440) );
  AO22X1_RVT U2676 ( .A1(\inq_ary[12][72] ), .A2(n3303), .A3(\inq_ary[3][72] ), 
        .A4(n3310), .Y(n2439) );
  AO22X1_RVT U2677 ( .A1(\inq_ary[5][72] ), .A2(n3298), .A3(\inq_ary[9][72] ), 
        .A4(n3314), .Y(n2438) );
  AO22X1_RVT U2678 ( .A1(\inq_ary[4][72] ), .A2(n3321), .A3(\inq_ary[10][72] ), 
        .A4(n3326), .Y(n2437) );
  NOR4X1_RVT U2679 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .Y(n2446)
         );
  AO22X1_RVT U2680 ( .A1(\inq_ary[14][72] ), .A2(n3325), .A3(\inq_ary[7][72] ), 
        .A4(n3322), .Y(n2444) );
  AO22X1_RVT U2681 ( .A1(\inq_ary[0][72] ), .A2(n3315), .A3(\inq_ary[2][72] ), 
        .A4(n3271), .Y(n2443) );
  AO22X1_RVT U2682 ( .A1(\inq_ary[1][72] ), .A2(n3324), .A3(\inq_ary[15][72] ), 
        .A4(n3312), .Y(n2442) );
  AO22X1_RVT U2683 ( .A1(\inq_ary[6][72] ), .A2(n3311), .A3(\inq_ary[8][72] ), 
        .A4(n3313), .Y(n2441) );
  NOR4X1_RVT U2684 ( .A1(n2444), .A2(n2443), .A3(n2442), .A4(n2441), .Y(n2445)
         );
  NAND2X0_RVT U2685 ( .A1(n2446), .A2(n2445), .Y(N333) );
  AO22X1_RVT U2686 ( .A1(\inq_ary[11][73] ), .A2(n3316), .A3(\inq_ary[1][73] ), 
        .A4(n3324), .Y(n2450) );
  AO22X1_RVT U2687 ( .A1(\inq_ary[8][73] ), .A2(n3313), .A3(\inq_ary[7][73] ), 
        .A4(n3322), .Y(n2449) );
  AO22X1_RVT U2688 ( .A1(\inq_ary[3][73] ), .A2(n3310), .A3(\inq_ary[10][73] ), 
        .A4(n3326), .Y(n2448) );
  AO22X1_RVT U2689 ( .A1(\inq_ary[12][73] ), .A2(n3303), .A3(\inq_ary[14][73] ), .A4(n3325), .Y(n2447) );
  NOR4X1_RVT U2690 ( .A1(n2450), .A2(n2449), .A3(n2448), .A4(n2447), .Y(n2456)
         );
  AO22X1_RVT U2691 ( .A1(\inq_ary[6][73] ), .A2(n3311), .A3(\inq_ary[13][73] ), 
        .A4(n3323), .Y(n2454) );
  AO22X1_RVT U2692 ( .A1(\inq_ary[9][73] ), .A2(n3314), .A3(\inq_ary[4][73] ), 
        .A4(n3321), .Y(n2453) );
  AO22X1_RVT U2693 ( .A1(\inq_ary[15][73] ), .A2(n3312), .A3(\inq_ary[0][73] ), 
        .A4(n3315), .Y(n2452) );
  AO22X1_RVT U2694 ( .A1(\inq_ary[2][73] ), .A2(n3271), .A3(\inq_ary[5][73] ), 
        .A4(n3298), .Y(n2451) );
  NOR4X1_RVT U2695 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .Y(n2455)
         );
  NAND2X0_RVT U2696 ( .A1(n2456), .A2(n2455), .Y(N334) );
  AO22X1_RVT U2697 ( .A1(\inq_ary[15][74] ), .A2(n3312), .A3(\inq_ary[12][74] ), .A4(n3303), .Y(n2460) );
  AO22X1_RVT U2698 ( .A1(\inq_ary[8][74] ), .A2(n3313), .A3(\inq_ary[9][74] ), 
        .A4(n3314), .Y(n2459) );
  AO22X1_RVT U2699 ( .A1(\inq_ary[4][74] ), .A2(n3321), .A3(\inq_ary[3][74] ), 
        .A4(n3310), .Y(n2458) );
  AO22X1_RVT U2700 ( .A1(\inq_ary[10][74] ), .A2(n3326), .A3(\inq_ary[7][74] ), 
        .A4(n3322), .Y(n2457) );
  NOR4X1_RVT U2701 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .Y(n2466)
         );
  AO22X1_RVT U2702 ( .A1(\inq_ary[14][74] ), .A2(n3325), .A3(\inq_ary[11][74] ), .A4(n3316), .Y(n2464) );
  AO22X1_RVT U2703 ( .A1(\inq_ary[1][74] ), .A2(n3324), .A3(\inq_ary[13][74] ), 
        .A4(n3323), .Y(n2463) );
  AO22X1_RVT U2704 ( .A1(\inq_ary[6][74] ), .A2(n3311), .A3(\inq_ary[0][74] ), 
        .A4(n3315), .Y(n2462) );
  AO22X1_RVT U2705 ( .A1(\inq_ary[5][74] ), .A2(n3298), .A3(\inq_ary[2][74] ), 
        .A4(n3271), .Y(n2461) );
  NOR4X1_RVT U2706 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .Y(n2465)
         );
  NAND2X0_RVT U2707 ( .A1(n2466), .A2(n2465), .Y(N335) );
  AO22X1_RVT U2708 ( .A1(\inq_ary[7][75] ), .A2(n3322), .A3(\inq_ary[12][75] ), 
        .A4(n3303), .Y(n2470) );
  AO22X1_RVT U2709 ( .A1(\inq_ary[0][75] ), .A2(n3315), .A3(\inq_ary[3][75] ), 
        .A4(n3310), .Y(n2469) );
  AO22X1_RVT U2710 ( .A1(\inq_ary[14][75] ), .A2(n3325), .A3(\inq_ary[9][75] ), 
        .A4(n3314), .Y(n2468) );
  AO22X1_RVT U2711 ( .A1(\inq_ary[8][75] ), .A2(n3313), .A3(\inq_ary[5][75] ), 
        .A4(n3298), .Y(n2467) );
  NOR4X1_RVT U2712 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .Y(n2476)
         );
  AO22X1_RVT U2713 ( .A1(\inq_ary[15][75] ), .A2(n3312), .A3(\inq_ary[1][75] ), 
        .A4(n3324), .Y(n2474) );
  AO22X1_RVT U2714 ( .A1(\inq_ary[11][75] ), .A2(n3316), .A3(\inq_ary[2][75] ), 
        .A4(n3271), .Y(n2473) );
  AO22X1_RVT U2715 ( .A1(\inq_ary[6][75] ), .A2(n3311), .A3(\inq_ary[10][75] ), 
        .A4(n3326), .Y(n2472) );
  AO22X1_RVT U2716 ( .A1(\inq_ary[4][75] ), .A2(n3321), .A3(\inq_ary[13][75] ), 
        .A4(n3323), .Y(n2471) );
  NOR4X1_RVT U2717 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .Y(n2475)
         );
  NAND2X0_RVT U2718 ( .A1(n2476), .A2(n2475), .Y(N336) );
  AO22X1_RVT U2719 ( .A1(\inq_ary[5][76] ), .A2(n3298), .A3(\inq_ary[9][76] ), 
        .A4(n3314), .Y(n2480) );
  AO22X1_RVT U2720 ( .A1(\inq_ary[6][76] ), .A2(n3311), .A3(\inq_ary[7][76] ), 
        .A4(n3322), .Y(n2479) );
  AO22X1_RVT U2721 ( .A1(\inq_ary[10][76] ), .A2(n3326), .A3(\inq_ary[11][76] ), .A4(n3316), .Y(n2478) );
  AO22X1_RVT U2722 ( .A1(\inq_ary[15][76] ), .A2(n3312), .A3(\inq_ary[4][76] ), 
        .A4(n3321), .Y(n2477) );
  NOR4X1_RVT U2723 ( .A1(n2480), .A2(n2479), .A3(n2478), .A4(n2477), .Y(n2486)
         );
  AO22X1_RVT U2724 ( .A1(\inq_ary[0][76] ), .A2(n3315), .A3(\inq_ary[14][76] ), 
        .A4(n3325), .Y(n2484) );
  AO22X1_RVT U2725 ( .A1(\inq_ary[3][76] ), .A2(n3310), .A3(\inq_ary[8][76] ), 
        .A4(n3313), .Y(n2483) );
  AO22X1_RVT U2726 ( .A1(\inq_ary[1][76] ), .A2(n3324), .A3(\inq_ary[2][76] ), 
        .A4(n3271), .Y(n2482) );
  AO22X1_RVT U2727 ( .A1(\inq_ary[13][76] ), .A2(n3323), .A3(\inq_ary[12][76] ), .A4(n3303), .Y(n2481) );
  NOR4X1_RVT U2728 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .Y(n2485)
         );
  NAND2X0_RVT U2729 ( .A1(n2486), .A2(n2485), .Y(N337) );
  AO22X1_RVT U2730 ( .A1(\inq_ary[1][77] ), .A2(n3324), .A3(\inq_ary[10][77] ), 
        .A4(n3326), .Y(n2490) );
  AO22X1_RVT U2731 ( .A1(\inq_ary[8][77] ), .A2(n3313), .A3(\inq_ary[5][77] ), 
        .A4(n3298), .Y(n2489) );
  AO22X1_RVT U2732 ( .A1(\inq_ary[11][77] ), .A2(n3316), .A3(\inq_ary[6][77] ), 
        .A4(n3311), .Y(n2488) );
  AO22X1_RVT U2733 ( .A1(\inq_ary[4][77] ), .A2(n3321), .A3(\inq_ary[14][77] ), 
        .A4(n3325), .Y(n2487) );
  NOR4X1_RVT U2734 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .Y(n2496)
         );
  AO22X1_RVT U2735 ( .A1(\inq_ary[3][77] ), .A2(n3310), .A3(\inq_ary[7][77] ), 
        .A4(n3322), .Y(n2494) );
  AO22X1_RVT U2736 ( .A1(\inq_ary[12][77] ), .A2(n3303), .A3(\inq_ary[13][77] ), .A4(n3323), .Y(n2493) );
  AO22X1_RVT U2737 ( .A1(\inq_ary[15][77] ), .A2(n3312), .A3(\inq_ary[0][77] ), 
        .A4(n3315), .Y(n2492) );
  AO22X1_RVT U2738 ( .A1(\inq_ary[9][77] ), .A2(n3314), .A3(\inq_ary[2][77] ), 
        .A4(n3271), .Y(n2491) );
  NOR4X1_RVT U2739 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), .Y(n2495)
         );
  NAND2X0_RVT U2740 ( .A1(n2496), .A2(n2495), .Y(N338) );
  AO22X1_RVT U2741 ( .A1(\inq_ary[15][78] ), .A2(n3312), .A3(\inq_ary[7][78] ), 
        .A4(n3322), .Y(n2500) );
  AO22X1_RVT U2742 ( .A1(\inq_ary[1][78] ), .A2(n3324), .A3(\inq_ary[14][78] ), 
        .A4(n3325), .Y(n2499) );
  AO22X1_RVT U2743 ( .A1(\inq_ary[3][78] ), .A2(n3310), .A3(\inq_ary[2][78] ), 
        .A4(n3271), .Y(n2498) );
  AO22X1_RVT U2744 ( .A1(\inq_ary[10][78] ), .A2(n3326), .A3(\inq_ary[13][78] ), .A4(n3323), .Y(n2497) );
  NOR4X1_RVT U2745 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .Y(n2506)
         );
  AO22X1_RVT U2746 ( .A1(\inq_ary[9][78] ), .A2(n3314), .A3(\inq_ary[6][78] ), 
        .A4(n3311), .Y(n2504) );
  AO22X1_RVT U2747 ( .A1(\inq_ary[12][78] ), .A2(n3303), .A3(\inq_ary[11][78] ), .A4(n3316), .Y(n2503) );
  AO22X1_RVT U2748 ( .A1(\inq_ary[5][78] ), .A2(n3298), .A3(\inq_ary[4][78] ), 
        .A4(n3321), .Y(n2502) );
  AO22X1_RVT U2749 ( .A1(\inq_ary[8][78] ), .A2(n3313), .A3(\inq_ary[0][78] ), 
        .A4(n3315), .Y(n2501) );
  NOR4X1_RVT U2750 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .Y(n2505)
         );
  NAND2X0_RVT U2751 ( .A1(n2506), .A2(n2505), .Y(N339) );
  AO22X1_RVT U2752 ( .A1(\inq_ary[11][79] ), .A2(n3316), .A3(\inq_ary[1][79] ), 
        .A4(n3324), .Y(n2510) );
  AO22X1_RVT U2753 ( .A1(\inq_ary[0][79] ), .A2(n3315), .A3(\inq_ary[12][79] ), 
        .A4(n3303), .Y(n2509) );
  AO22X1_RVT U2754 ( .A1(\inq_ary[6][79] ), .A2(n3311), .A3(\inq_ary[9][79] ), 
        .A4(n3314), .Y(n2508) );
  AO22X1_RVT U2755 ( .A1(\inq_ary[13][79] ), .A2(n3323), .A3(\inq_ary[14][79] ), .A4(n3325), .Y(n2507) );
  NOR4X1_RVT U2756 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .Y(n2516)
         );
  AO22X1_RVT U2757 ( .A1(\inq_ary[8][79] ), .A2(n3313), .A3(\inq_ary[5][79] ), 
        .A4(n3298), .Y(n2514) );
  AO22X1_RVT U2758 ( .A1(\inq_ary[4][79] ), .A2(n3321), .A3(\inq_ary[2][79] ), 
        .A4(n3271), .Y(n2513) );
  AO22X1_RVT U2759 ( .A1(\inq_ary[3][79] ), .A2(n3310), .A3(\inq_ary[10][79] ), 
        .A4(n3326), .Y(n2512) );
  AO22X1_RVT U2760 ( .A1(\inq_ary[15][79] ), .A2(n3312), .A3(\inq_ary[7][79] ), 
        .A4(n3322), .Y(n2511) );
  NOR4X1_RVT U2761 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .Y(n2515)
         );
  NAND2X0_RVT U2762 ( .A1(n2516), .A2(n2515), .Y(N340) );
  AO22X1_RVT U2763 ( .A1(\inq_ary[12][80] ), .A2(n3303), .A3(\inq_ary[11][80] ), .A4(n3316), .Y(n2520) );
  AO22X1_RVT U2764 ( .A1(\inq_ary[5][80] ), .A2(n3298), .A3(\inq_ary[2][80] ), 
        .A4(n3271), .Y(n2519) );
  AO22X1_RVT U2765 ( .A1(\inq_ary[3][80] ), .A2(n3310), .A3(\inq_ary[0][80] ), 
        .A4(n3315), .Y(n2518) );
  AO22X1_RVT U2766 ( .A1(\inq_ary[15][80] ), .A2(n3312), .A3(\inq_ary[8][80] ), 
        .A4(n3313), .Y(n2517) );
  NOR4X1_RVT U2767 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .Y(n2526)
         );
  AO22X1_RVT U2768 ( .A1(\inq_ary[14][80] ), .A2(n3325), .A3(\inq_ary[13][80] ), .A4(n3323), .Y(n2524) );
  AO22X1_RVT U2769 ( .A1(\inq_ary[7][80] ), .A2(n3322), .A3(\inq_ary[10][80] ), 
        .A4(n3326), .Y(n2523) );
  AO22X1_RVT U2770 ( .A1(\inq_ary[1][80] ), .A2(n3324), .A3(\inq_ary[4][80] ), 
        .A4(n3321), .Y(n2522) );
  AO22X1_RVT U2771 ( .A1(\inq_ary[6][80] ), .A2(n3311), .A3(\inq_ary[9][80] ), 
        .A4(n3314), .Y(n2521) );
  NOR4X1_RVT U2772 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .Y(n2525)
         );
  NAND2X0_RVT U2773 ( .A1(n2526), .A2(n2525), .Y(N341) );
  AO22X1_RVT U2774 ( .A1(\inq_ary[12][81] ), .A2(n3303), .A3(\inq_ary[0][81] ), 
        .A4(n3315), .Y(n2530) );
  AO22X1_RVT U2775 ( .A1(\inq_ary[6][81] ), .A2(n3311), .A3(\inq_ary[1][81] ), 
        .A4(n3324), .Y(n2529) );
  AO22X1_RVT U2776 ( .A1(\inq_ary[9][81] ), .A2(n3314), .A3(\inq_ary[8][81] ), 
        .A4(n3313), .Y(n2528) );
  AO22X1_RVT U2777 ( .A1(\inq_ary[10][81] ), .A2(n3326), .A3(\inq_ary[7][81] ), 
        .A4(n3322), .Y(n2527) );
  NOR4X1_RVT U2778 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .Y(n2536)
         );
  AO22X1_RVT U2779 ( .A1(\inq_ary[14][81] ), .A2(n3325), .A3(\inq_ary[3][81] ), 
        .A4(n3310), .Y(n2534) );
  AO22X1_RVT U2780 ( .A1(\inq_ary[13][81] ), .A2(n3323), .A3(\inq_ary[5][81] ), 
        .A4(n3298), .Y(n2533) );
  AO22X1_RVT U2781 ( .A1(\inq_ary[4][81] ), .A2(n3321), .A3(\inq_ary[2][81] ), 
        .A4(n3271), .Y(n2532) );
  AO22X1_RVT U2782 ( .A1(\inq_ary[15][81] ), .A2(n3312), .A3(\inq_ary[11][81] ), .A4(n3316), .Y(n2531) );
  NOR4X1_RVT U2783 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), .Y(n2535)
         );
  NAND2X0_RVT U2784 ( .A1(n2536), .A2(n2535), .Y(N342) );
  AO22X1_RVT U2785 ( .A1(\inq_ary[4][82] ), .A2(n3321), .A3(\inq_ary[1][82] ), 
        .A4(n3324), .Y(n2540) );
  AO22X1_RVT U2786 ( .A1(\inq_ary[13][82] ), .A2(n3323), .A3(\inq_ary[5][82] ), 
        .A4(n3298), .Y(n2539) );
  AO22X1_RVT U2787 ( .A1(\inq_ary[9][82] ), .A2(n3314), .A3(\inq_ary[12][82] ), 
        .A4(n3303), .Y(n2538) );
  AO22X1_RVT U2788 ( .A1(\inq_ary[10][82] ), .A2(n3326), .A3(\inq_ary[11][82] ), .A4(n3316), .Y(n2537) );
  NOR4X1_RVT U2789 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .Y(n2546)
         );
  AO22X1_RVT U2790 ( .A1(\inq_ary[14][82] ), .A2(n3325), .A3(\inq_ary[6][82] ), 
        .A4(n3311), .Y(n2544) );
  AO22X1_RVT U2791 ( .A1(\inq_ary[15][82] ), .A2(n3312), .A3(\inq_ary[7][82] ), 
        .A4(n3322), .Y(n2543) );
  AO22X1_RVT U2792 ( .A1(\inq_ary[8][82] ), .A2(n3313), .A3(\inq_ary[3][82] ), 
        .A4(n3310), .Y(n2542) );
  AO22X1_RVT U2793 ( .A1(\inq_ary[0][82] ), .A2(n3315), .A3(\inq_ary[2][82] ), 
        .A4(n3271), .Y(n2541) );
  NOR4X1_RVT U2794 ( .A1(n2544), .A2(n2543), .A3(n2542), .A4(n2541), .Y(n2545)
         );
  NAND2X0_RVT U2795 ( .A1(n2546), .A2(n2545), .Y(N343) );
  AO22X1_RVT U2796 ( .A1(\inq_ary[12][83] ), .A2(n3303), .A3(\inq_ary[0][83] ), 
        .A4(n3315), .Y(n2550) );
  AO22X1_RVT U2797 ( .A1(\inq_ary[5][83] ), .A2(n3298), .A3(\inq_ary[8][83] ), 
        .A4(n3313), .Y(n2549) );
  AO22X1_RVT U2798 ( .A1(\inq_ary[15][83] ), .A2(n3312), .A3(\inq_ary[1][83] ), 
        .A4(n3324), .Y(n2548) );
  AO22X1_RVT U2799 ( .A1(\inq_ary[14][83] ), .A2(n3325), .A3(\inq_ary[9][83] ), 
        .A4(n3314), .Y(n2547) );
  NOR4X1_RVT U2800 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .Y(n2556)
         );
  AO22X1_RVT U2801 ( .A1(\inq_ary[2][83] ), .A2(n3271), .A3(\inq_ary[4][83] ), 
        .A4(n3321), .Y(n2554) );
  AO22X1_RVT U2802 ( .A1(\inq_ary[3][83] ), .A2(n3310), .A3(\inq_ary[6][83] ), 
        .A4(n3311), .Y(n2553) );
  AO22X1_RVT U2803 ( .A1(\inq_ary[11][83] ), .A2(n3316), .A3(\inq_ary[13][83] ), .A4(n3323), .Y(n2552) );
  AO22X1_RVT U2804 ( .A1(\inq_ary[7][83] ), .A2(n3322), .A3(\inq_ary[10][83] ), 
        .A4(n3326), .Y(n2551) );
  NOR4X1_RVT U2805 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .Y(n2555)
         );
  NAND2X0_RVT U2806 ( .A1(n2556), .A2(n2555), .Y(N344) );
  AO22X1_RVT U2807 ( .A1(\inq_ary[8][84] ), .A2(n3313), .A3(\inq_ary[15][84] ), 
        .A4(n3312), .Y(n2560) );
  AO22X1_RVT U2808 ( .A1(\inq_ary[14][84] ), .A2(n3325), .A3(\inq_ary[7][84] ), 
        .A4(n3322), .Y(n2559) );
  AO22X1_RVT U2809 ( .A1(\inq_ary[12][84] ), .A2(n3303), .A3(\inq_ary[10][84] ), .A4(n3326), .Y(n2558) );
  AO22X1_RVT U2810 ( .A1(\inq_ary[3][84] ), .A2(n3310), .A3(\inq_ary[5][84] ), 
        .A4(n3298), .Y(n2557) );
  NOR4X1_RVT U2811 ( .A1(n2560), .A2(n2559), .A3(n2558), .A4(n2557), .Y(n2566)
         );
  AO22X1_RVT U2812 ( .A1(\inq_ary[2][84] ), .A2(n3271), .A3(\inq_ary[4][84] ), 
        .A4(n3321), .Y(n2564) );
  AO22X1_RVT U2813 ( .A1(\inq_ary[6][84] ), .A2(n3311), .A3(\inq_ary[1][84] ), 
        .A4(n3324), .Y(n2563) );
  AO22X1_RVT U2814 ( .A1(\inq_ary[11][84] ), .A2(n3316), .A3(\inq_ary[13][84] ), .A4(n3323), .Y(n2562) );
  AO22X1_RVT U2815 ( .A1(\inq_ary[0][84] ), .A2(n3315), .A3(\inq_ary[9][84] ), 
        .A4(n3314), .Y(n2561) );
  NOR4X1_RVT U2816 ( .A1(n2564), .A2(n2563), .A3(n2562), .A4(n2561), .Y(n2565)
         );
  NAND2X0_RVT U2817 ( .A1(n2566), .A2(n2565), .Y(N345) );
  AO22X1_RVT U2818 ( .A1(\inq_ary[1][85] ), .A2(n3324), .A3(\inq_ary[15][85] ), 
        .A4(n3312), .Y(n2570) );
  AO22X1_RVT U2819 ( .A1(\inq_ary[7][85] ), .A2(n3322), .A3(\inq_ary[11][85] ), 
        .A4(n3316), .Y(n2569) );
  AO22X1_RVT U2820 ( .A1(\inq_ary[6][85] ), .A2(n3311), .A3(\inq_ary[13][85] ), 
        .A4(n3323), .Y(n2568) );
  AO22X1_RVT U2821 ( .A1(\inq_ary[3][85] ), .A2(n3310), .A3(\inq_ary[8][85] ), 
        .A4(n3313), .Y(n2567) );
  NOR4X1_RVT U2822 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), .Y(n2576)
         );
  AO22X1_RVT U2823 ( .A1(\inq_ary[5][85] ), .A2(n3298), .A3(\inq_ary[9][85] ), 
        .A4(n3314), .Y(n2574) );
  AO22X1_RVT U2824 ( .A1(\inq_ary[12][85] ), .A2(n3303), .A3(\inq_ary[0][85] ), 
        .A4(n3315), .Y(n2573) );
  AO22X1_RVT U2825 ( .A1(\inq_ary[2][85] ), .A2(n3271), .A3(\inq_ary[4][85] ), 
        .A4(n3321), .Y(n2572) );
  AO22X1_RVT U2826 ( .A1(\inq_ary[14][85] ), .A2(n3325), .A3(\inq_ary[10][85] ), .A4(n3326), .Y(n2571) );
  NOR4X1_RVT U2827 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .Y(n2575)
         );
  NAND2X0_RVT U2828 ( .A1(n2576), .A2(n2575), .Y(N346) );
  AO22X1_RVT U2829 ( .A1(\inq_ary[5][86] ), .A2(n3298), .A3(\inq_ary[13][86] ), 
        .A4(n3323), .Y(n2580) );
  AO22X1_RVT U2830 ( .A1(\inq_ary[4][86] ), .A2(n3321), .A3(\inq_ary[0][86] ), 
        .A4(n3315), .Y(n2579) );
  AO22X1_RVT U2831 ( .A1(\inq_ary[14][86] ), .A2(n3325), .A3(\inq_ary[11][86] ), .A4(n3316), .Y(n2578) );
  AO22X1_RVT U2832 ( .A1(\inq_ary[7][86] ), .A2(n3322), .A3(\inq_ary[1][86] ), 
        .A4(n3324), .Y(n2577) );
  NOR4X1_RVT U2833 ( .A1(n2580), .A2(n2579), .A3(n2578), .A4(n2577), .Y(n2586)
         );
  AO22X1_RVT U2834 ( .A1(\inq_ary[12][86] ), .A2(n3303), .A3(\inq_ary[2][86] ), 
        .A4(n3271), .Y(n2584) );
  AO22X1_RVT U2835 ( .A1(\inq_ary[9][86] ), .A2(n3314), .A3(\inq_ary[10][86] ), 
        .A4(n3326), .Y(n2583) );
  AO22X1_RVT U2836 ( .A1(\inq_ary[8][86] ), .A2(n3313), .A3(\inq_ary[6][86] ), 
        .A4(n3311), .Y(n2582) );
  AO22X1_RVT U2837 ( .A1(\inq_ary[3][86] ), .A2(n3310), .A3(\inq_ary[15][86] ), 
        .A4(n3312), .Y(n2581) );
  NOR4X1_RVT U2838 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .Y(n2585)
         );
  NAND2X0_RVT U2839 ( .A1(n2586), .A2(n2585), .Y(N347) );
  AO22X1_RVT U2840 ( .A1(\inq_ary[14][87] ), .A2(n3325), .A3(\inq_ary[11][87] ), .A4(n3316), .Y(n2590) );
  AO22X1_RVT U2841 ( .A1(\inq_ary[15][87] ), .A2(n3312), .A3(\inq_ary[1][87] ), 
        .A4(n3324), .Y(n2589) );
  AO22X1_RVT U2842 ( .A1(\inq_ary[0][87] ), .A2(n3315), .A3(\inq_ary[3][87] ), 
        .A4(n3310), .Y(n2588) );
  AO22X1_RVT U2843 ( .A1(\inq_ary[9][87] ), .A2(n3314), .A3(\inq_ary[5][87] ), 
        .A4(n3298), .Y(n2587) );
  NOR4X1_RVT U2844 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .Y(n2596)
         );
  AO22X1_RVT U2845 ( .A1(\inq_ary[7][87] ), .A2(n3322), .A3(\inq_ary[2][87] ), 
        .A4(n3271), .Y(n2594) );
  AO22X1_RVT U2846 ( .A1(\inq_ary[13][87] ), .A2(n3323), .A3(\inq_ary[10][87] ), .A4(n3326), .Y(n2593) );
  AO22X1_RVT U2847 ( .A1(\inq_ary[8][87] ), .A2(n3313), .A3(\inq_ary[12][87] ), 
        .A4(n3303), .Y(n2592) );
  AO22X1_RVT U2848 ( .A1(\inq_ary[4][87] ), .A2(n3321), .A3(\inq_ary[6][87] ), 
        .A4(n3311), .Y(n2591) );
  NOR4X1_RVT U2849 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .Y(n2595)
         );
  NAND2X0_RVT U2850 ( .A1(n2596), .A2(n2595), .Y(N348) );
  AO22X1_RVT U2851 ( .A1(\inq_ary[1][88] ), .A2(n3324), .A3(\inq_ary[11][88] ), 
        .A4(n3316), .Y(n2600) );
  AO22X1_RVT U2852 ( .A1(\inq_ary[9][88] ), .A2(n3314), .A3(\inq_ary[10][88] ), 
        .A4(n3326), .Y(n2599) );
  AO22X1_RVT U2853 ( .A1(\inq_ary[2][88] ), .A2(n3271), .A3(\inq_ary[14][88] ), 
        .A4(n3325), .Y(n2598) );
  AO22X1_RVT U2854 ( .A1(\inq_ary[4][88] ), .A2(n3321), .A3(\inq_ary[3][88] ), 
        .A4(n3310), .Y(n2597) );
  NOR4X1_RVT U2855 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .Y(n2606)
         );
  AO22X1_RVT U2856 ( .A1(\inq_ary[12][88] ), .A2(n3303), .A3(\inq_ary[13][88] ), .A4(n3323), .Y(n2604) );
  AO22X1_RVT U2857 ( .A1(\inq_ary[6][88] ), .A2(n3311), .A3(\inq_ary[5][88] ), 
        .A4(n3298), .Y(n2603) );
  AO22X1_RVT U2858 ( .A1(\inq_ary[7][88] ), .A2(n3322), .A3(\inq_ary[8][88] ), 
        .A4(n3313), .Y(n2602) );
  AO22X1_RVT U2859 ( .A1(\inq_ary[0][88] ), .A2(n3315), .A3(\inq_ary[15][88] ), 
        .A4(n3312), .Y(n2601) );
  NOR4X1_RVT U2860 ( .A1(n2604), .A2(n2603), .A3(n2602), .A4(n2601), .Y(n2605)
         );
  NAND2X0_RVT U2861 ( .A1(n2606), .A2(n2605), .Y(N349) );
  AO22X1_RVT U2862 ( .A1(\inq_ary[4][89] ), .A2(n3321), .A3(\inq_ary[1][89] ), 
        .A4(n3324), .Y(n2610) );
  AO22X1_RVT U2863 ( .A1(\inq_ary[5][89] ), .A2(n3298), .A3(\inq_ary[9][89] ), 
        .A4(n3314), .Y(n2609) );
  AO22X1_RVT U2864 ( .A1(\inq_ary[0][89] ), .A2(n3315), .A3(\inq_ary[2][89] ), 
        .A4(n3271), .Y(n2608) );
  AO22X1_RVT U2865 ( .A1(\inq_ary[3][89] ), .A2(n3310), .A3(\inq_ary[7][89] ), 
        .A4(n3322), .Y(n2607) );
  NOR4X1_RVT U2866 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .Y(n2616)
         );
  AO22X1_RVT U2867 ( .A1(\inq_ary[13][89] ), .A2(n3323), .A3(\inq_ary[11][89] ), .A4(n3316), .Y(n2614) );
  AO22X1_RVT U2868 ( .A1(\inq_ary[14][89] ), .A2(n3325), .A3(\inq_ary[8][89] ), 
        .A4(n3313), .Y(n2613) );
  AO22X1_RVT U2869 ( .A1(\inq_ary[10][89] ), .A2(n3326), .A3(\inq_ary[15][89] ), .A4(n3312), .Y(n2612) );
  AO22X1_RVT U2870 ( .A1(\inq_ary[12][89] ), .A2(n3303), .A3(\inq_ary[6][89] ), 
        .A4(n3311), .Y(n2611) );
  NOR4X1_RVT U2871 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .Y(n2615)
         );
  NAND2X0_RVT U2872 ( .A1(n2616), .A2(n2615), .Y(N350) );
  AO22X1_RVT U2873 ( .A1(\inq_ary[5][90] ), .A2(n3298), .A3(\inq_ary[4][90] ), 
        .A4(n3321), .Y(n2620) );
  AO22X1_RVT U2874 ( .A1(\inq_ary[10][90] ), .A2(n3326), .A3(\inq_ary[1][90] ), 
        .A4(n3324), .Y(n2619) );
  AO22X1_RVT U2875 ( .A1(\inq_ary[0][90] ), .A2(n3315), .A3(\inq_ary[11][90] ), 
        .A4(n3316), .Y(n2618) );
  AO22X1_RVT U2876 ( .A1(\inq_ary[14][90] ), .A2(n3325), .A3(\inq_ary[12][90] ), .A4(n3303), .Y(n2617) );
  NOR4X1_RVT U2877 ( .A1(n2620), .A2(n2619), .A3(n2618), .A4(n2617), .Y(n2626)
         );
  AO22X1_RVT U2878 ( .A1(\inq_ary[6][90] ), .A2(n3311), .A3(\inq_ary[8][90] ), 
        .A4(n3313), .Y(n2624) );
  AO22X1_RVT U2879 ( .A1(\inq_ary[13][90] ), .A2(n3323), .A3(\inq_ary[3][90] ), 
        .A4(n3310), .Y(n2623) );
  AO22X1_RVT U2880 ( .A1(\inq_ary[7][90] ), .A2(n3322), .A3(\inq_ary[15][90] ), 
        .A4(n3312), .Y(n2622) );
  AO22X1_RVT U2881 ( .A1(\inq_ary[2][90] ), .A2(n3271), .A3(\inq_ary[9][90] ), 
        .A4(n3314), .Y(n2621) );
  NOR4X1_RVT U2882 ( .A1(n2624), .A2(n2623), .A3(n2622), .A4(n2621), .Y(n2625)
         );
  NAND2X0_RVT U2883 ( .A1(n2626), .A2(n2625), .Y(N351) );
  AO22X1_RVT U2884 ( .A1(\inq_ary[0][91] ), .A2(n3315), .A3(\inq_ary[4][91] ), 
        .A4(n3321), .Y(n2630) );
  AO22X1_RVT U2885 ( .A1(\inq_ary[3][91] ), .A2(n3310), .A3(\inq_ary[12][91] ), 
        .A4(n3303), .Y(n2629) );
  AO22X1_RVT U2886 ( .A1(\inq_ary[6][91] ), .A2(n3311), .A3(\inq_ary[13][91] ), 
        .A4(n3323), .Y(n2628) );
  AO22X1_RVT U2887 ( .A1(\inq_ary[7][91] ), .A2(n3322), .A3(\inq_ary[14][91] ), 
        .A4(n3325), .Y(n2627) );
  NOR4X1_RVT U2888 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .Y(n2636)
         );
  AO22X1_RVT U2889 ( .A1(\inq_ary[1][91] ), .A2(n3324), .A3(\inq_ary[9][91] ), 
        .A4(n3314), .Y(n2634) );
  AO22X1_RVT U2890 ( .A1(\inq_ary[8][91] ), .A2(n3313), .A3(\inq_ary[11][91] ), 
        .A4(n3316), .Y(n2633) );
  AO22X1_RVT U2891 ( .A1(\inq_ary[15][91] ), .A2(n3312), .A3(\inq_ary[5][91] ), 
        .A4(n3298), .Y(n2632) );
  AO22X1_RVT U2892 ( .A1(\inq_ary[10][91] ), .A2(n3326), .A3(\inq_ary[2][91] ), 
        .A4(n3271), .Y(n2631) );
  NOR4X1_RVT U2893 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .Y(n2635)
         );
  NAND2X0_RVT U2894 ( .A1(n2636), .A2(n2635), .Y(N352) );
  AO22X1_RVT U2895 ( .A1(\inq_ary[4][92] ), .A2(n3321), .A3(\inq_ary[1][92] ), 
        .A4(n3324), .Y(n2640) );
  AO22X1_RVT U2896 ( .A1(\inq_ary[7][92] ), .A2(n3322), .A3(\inq_ary[5][92] ), 
        .A4(n3298), .Y(n2639) );
  AO22X1_RVT U2897 ( .A1(\inq_ary[8][92] ), .A2(n3313), .A3(\inq_ary[11][92] ), 
        .A4(n3316), .Y(n2638) );
  AO22X1_RVT U2898 ( .A1(\inq_ary[13][92] ), .A2(n3323), .A3(\inq_ary[9][92] ), 
        .A4(n3314), .Y(n2637) );
  NOR4X1_RVT U2899 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .Y(n2646)
         );
  AO22X1_RVT U2900 ( .A1(\inq_ary[12][92] ), .A2(n3303), .A3(\inq_ary[0][92] ), 
        .A4(n3315), .Y(n2644) );
  AO22X1_RVT U2901 ( .A1(\inq_ary[14][92] ), .A2(n3325), .A3(\inq_ary[6][92] ), 
        .A4(n3311), .Y(n2643) );
  AO22X1_RVT U2902 ( .A1(\inq_ary[2][92] ), .A2(n3271), .A3(\inq_ary[15][92] ), 
        .A4(n3312), .Y(n2642) );
  AO22X1_RVT U2903 ( .A1(\inq_ary[10][92] ), .A2(n3326), .A3(\inq_ary[3][92] ), 
        .A4(n3310), .Y(n2641) );
  NOR4X1_RVT U2904 ( .A1(n2644), .A2(n2643), .A3(n2642), .A4(n2641), .Y(n2645)
         );
  NAND2X0_RVT U2905 ( .A1(n2646), .A2(n2645), .Y(N353) );
  AO22X1_RVT U2906 ( .A1(\inq_ary[12][93] ), .A2(n3303), .A3(\inq_ary[4][93] ), 
        .A4(n3321), .Y(n2650) );
  AO22X1_RVT U2907 ( .A1(\inq_ary[5][93] ), .A2(n3298), .A3(\inq_ary[10][93] ), 
        .A4(n3326), .Y(n2649) );
  AO22X1_RVT U2908 ( .A1(\inq_ary[1][93] ), .A2(n3324), .A3(\inq_ary[15][93] ), 
        .A4(n3312), .Y(n2648) );
  AO22X1_RVT U2909 ( .A1(\inq_ary[3][93] ), .A2(n3310), .A3(\inq_ary[11][93] ), 
        .A4(n3316), .Y(n2647) );
  NOR4X1_RVT U2910 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .Y(n2656)
         );
  AO22X1_RVT U2911 ( .A1(\inq_ary[9][93] ), .A2(n3314), .A3(\inq_ary[6][93] ), 
        .A4(n3311), .Y(n2654) );
  AO22X1_RVT U2912 ( .A1(\inq_ary[14][93] ), .A2(n3325), .A3(\inq_ary[0][93] ), 
        .A4(n3315), .Y(n2653) );
  AO22X1_RVT U2913 ( .A1(\inq_ary[13][93] ), .A2(n3323), .A3(\inq_ary[7][93] ), 
        .A4(n3322), .Y(n2652) );
  AO22X1_RVT U2914 ( .A1(\inq_ary[2][93] ), .A2(n3271), .A3(\inq_ary[8][93] ), 
        .A4(n3313), .Y(n2651) );
  NOR4X1_RVT U2915 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .Y(n2655)
         );
  NAND2X0_RVT U2916 ( .A1(n2656), .A2(n2655), .Y(N354) );
  AO22X1_RVT U2917 ( .A1(\inq_ary[13][94] ), .A2(n3323), .A3(\inq_ary[11][94] ), .A4(n3316), .Y(n2660) );
  AO22X1_RVT U2918 ( .A1(\inq_ary[15][94] ), .A2(n3312), .A3(\inq_ary[4][94] ), 
        .A4(n3321), .Y(n2659) );
  AO22X1_RVT U2919 ( .A1(\inq_ary[7][94] ), .A2(n3322), .A3(\inq_ary[3][94] ), 
        .A4(n3310), .Y(n2658) );
  AO22X1_RVT U2920 ( .A1(\inq_ary[6][94] ), .A2(n3311), .A3(\inq_ary[8][94] ), 
        .A4(n3313), .Y(n2657) );
  NOR4X1_RVT U2921 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .Y(n2666)
         );
  AO22X1_RVT U2922 ( .A1(\inq_ary[1][94] ), .A2(n3324), .A3(\inq_ary[0][94] ), 
        .A4(n3315), .Y(n2664) );
  AO22X1_RVT U2923 ( .A1(\inq_ary[2][94] ), .A2(n3271), .A3(\inq_ary[10][94] ), 
        .A4(n3326), .Y(n2663) );
  AO22X1_RVT U2924 ( .A1(\inq_ary[12][94] ), .A2(n3303), .A3(\inq_ary[5][94] ), 
        .A4(n3298), .Y(n2662) );
  AO22X1_RVT U2925 ( .A1(\inq_ary[14][94] ), .A2(n3325), .A3(\inq_ary[9][94] ), 
        .A4(n3314), .Y(n2661) );
  NOR4X1_RVT U2926 ( .A1(n2664), .A2(n2663), .A3(n2662), .A4(n2661), .Y(n2665)
         );
  NAND2X0_RVT U2927 ( .A1(n2666), .A2(n2665), .Y(N355) );
  AO22X1_RVT U2928 ( .A1(\inq_ary[9][95] ), .A2(n3314), .A3(\inq_ary[0][95] ), 
        .A4(n3315), .Y(n2670) );
  AO22X1_RVT U2929 ( .A1(\inq_ary[2][95] ), .A2(n3271), .A3(\inq_ary[14][95] ), 
        .A4(n3325), .Y(n2669) );
  AO22X1_RVT U2930 ( .A1(\inq_ary[8][95] ), .A2(n3313), .A3(\inq_ary[13][95] ), 
        .A4(n3323), .Y(n2668) );
  AO22X1_RVT U2931 ( .A1(\inq_ary[11][95] ), .A2(n3316), .A3(\inq_ary[15][95] ), .A4(n3312), .Y(n2667) );
  NOR4X1_RVT U2932 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .Y(n2676)
         );
  AO22X1_RVT U2933 ( .A1(\inq_ary[1][95] ), .A2(n3324), .A3(\inq_ary[6][95] ), 
        .A4(n3311), .Y(n2674) );
  AO22X1_RVT U2934 ( .A1(\inq_ary[12][95] ), .A2(n3303), .A3(\inq_ary[4][95] ), 
        .A4(n3321), .Y(n2673) );
  AO22X1_RVT U2935 ( .A1(\inq_ary[7][95] ), .A2(n3322), .A3(\inq_ary[10][95] ), 
        .A4(n3326), .Y(n2672) );
  AO22X1_RVT U2936 ( .A1(\inq_ary[5][95] ), .A2(n3298), .A3(\inq_ary[3][95] ), 
        .A4(n3310), .Y(n2671) );
  NOR4X1_RVT U2937 ( .A1(n2674), .A2(n2673), .A3(n2672), .A4(n2671), .Y(n2675)
         );
  NAND2X0_RVT U2938 ( .A1(n2676), .A2(n2675), .Y(N356) );
  AO22X1_RVT U2939 ( .A1(\inq_ary[2][96] ), .A2(n3271), .A3(\inq_ary[10][96] ), 
        .A4(n3326), .Y(n2680) );
  AO22X1_RVT U2940 ( .A1(\inq_ary[11][96] ), .A2(n3316), .A3(\inq_ary[9][96] ), 
        .A4(n3314), .Y(n2679) );
  AO22X1_RVT U2941 ( .A1(\inq_ary[3][96] ), .A2(n3310), .A3(\inq_ary[13][96] ), 
        .A4(n3323), .Y(n2678) );
  AO22X1_RVT U2942 ( .A1(\inq_ary[4][96] ), .A2(n3321), .A3(\inq_ary[5][96] ), 
        .A4(n3298), .Y(n2677) );
  NOR4X1_RVT U2943 ( .A1(n2680), .A2(n2679), .A3(n2678), .A4(n2677), .Y(n2686)
         );
  AO22X1_RVT U2944 ( .A1(\inq_ary[8][96] ), .A2(n3313), .A3(\inq_ary[6][96] ), 
        .A4(n3311), .Y(n2684) );
  AO22X1_RVT U2945 ( .A1(\inq_ary[1][96] ), .A2(n3324), .A3(\inq_ary[0][96] ), 
        .A4(n3315), .Y(n2683) );
  AO22X1_RVT U2946 ( .A1(\inq_ary[14][96] ), .A2(n3325), .A3(\inq_ary[12][96] ), .A4(n3303), .Y(n2682) );
  AO22X1_RVT U2947 ( .A1(\inq_ary[7][96] ), .A2(n3322), .A3(\inq_ary[15][96] ), 
        .A4(n3312), .Y(n2681) );
  NOR4X1_RVT U2948 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .Y(n2685)
         );
  NAND2X0_RVT U2949 ( .A1(n2686), .A2(n2685), .Y(N357) );
  AO22X1_RVT U2950 ( .A1(\inq_ary[0][97] ), .A2(n3315), .A3(\inq_ary[5][97] ), 
        .A4(n3298), .Y(n2690) );
  AO22X1_RVT U2951 ( .A1(\inq_ary[2][97] ), .A2(n3271), .A3(\inq_ary[14][97] ), 
        .A4(n3325), .Y(n2689) );
  AO22X1_RVT U2952 ( .A1(\inq_ary[9][97] ), .A2(n3314), .A3(\inq_ary[8][97] ), 
        .A4(n3313), .Y(n2688) );
  AO22X1_RVT U2953 ( .A1(\inq_ary[7][97] ), .A2(n3322), .A3(\inq_ary[11][97] ), 
        .A4(n3316), .Y(n2687) );
  NOR4X1_RVT U2954 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .Y(n2696)
         );
  AO22X1_RVT U2955 ( .A1(\inq_ary[10][97] ), .A2(n3326), .A3(\inq_ary[12][97] ), .A4(n3303), .Y(n2694) );
  AO22X1_RVT U2956 ( .A1(\inq_ary[13][97] ), .A2(n3323), .A3(\inq_ary[1][97] ), 
        .A4(n3324), .Y(n2693) );
  AO22X1_RVT U2957 ( .A1(\inq_ary[6][97] ), .A2(n3311), .A3(\inq_ary[15][97] ), 
        .A4(n3312), .Y(n2692) );
  AO22X1_RVT U2958 ( .A1(\inq_ary[3][97] ), .A2(n3310), .A3(\inq_ary[4][97] ), 
        .A4(n3321), .Y(n2691) );
  NOR4X1_RVT U2959 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .Y(n2695)
         );
  NAND2X0_RVT U2960 ( .A1(n2696), .A2(n2695), .Y(N358) );
  AO22X1_RVT U2961 ( .A1(\inq_ary[15][98] ), .A2(n3312), .A3(\inq_ary[12][98] ), .A4(n3303), .Y(n2700) );
  AO22X1_RVT U2962 ( .A1(\inq_ary[7][98] ), .A2(n3322), .A3(\inq_ary[9][98] ), 
        .A4(n3314), .Y(n2699) );
  AO22X1_RVT U2963 ( .A1(\inq_ary[10][98] ), .A2(n3326), .A3(\inq_ary[14][98] ), .A4(n3325), .Y(n2698) );
  AO22X1_RVT U2964 ( .A1(\inq_ary[0][98] ), .A2(n3315), .A3(\inq_ary[6][98] ), 
        .A4(n3311), .Y(n2697) );
  NOR4X1_RVT U2965 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .Y(n2706)
         );
  AO22X1_RVT U2966 ( .A1(\inq_ary[1][98] ), .A2(n3324), .A3(\inq_ary[5][98] ), 
        .A4(n3298), .Y(n2704) );
  AO22X1_RVT U2967 ( .A1(\inq_ary[11][98] ), .A2(n3316), .A3(\inq_ary[4][98] ), 
        .A4(n3321), .Y(n2703) );
  AO22X1_RVT U2968 ( .A1(\inq_ary[3][98] ), .A2(n3310), .A3(\inq_ary[8][98] ), 
        .A4(n3313), .Y(n2702) );
  AO22X1_RVT U2969 ( .A1(\inq_ary[13][98] ), .A2(n3323), .A3(\inq_ary[2][98] ), 
        .A4(n3271), .Y(n2701) );
  NOR4X1_RVT U2970 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .Y(n2705)
         );
  NAND2X0_RVT U2971 ( .A1(n2706), .A2(n2705), .Y(N359) );
  AO22X1_RVT U2972 ( .A1(\inq_ary[5][99] ), .A2(n3298), .A3(\inq_ary[10][99] ), 
        .A4(n3326), .Y(n2710) );
  AO22X1_RVT U2973 ( .A1(\inq_ary[8][99] ), .A2(n3313), .A3(\inq_ary[4][99] ), 
        .A4(n3321), .Y(n2709) );
  AO22X1_RVT U2974 ( .A1(\inq_ary[15][99] ), .A2(n3312), .A3(\inq_ary[9][99] ), 
        .A4(n3314), .Y(n2708) );
  AO22X1_RVT U2975 ( .A1(\inq_ary[0][99] ), .A2(n3315), .A3(\inq_ary[3][99] ), 
        .A4(n3310), .Y(n2707) );
  NOR4X1_RVT U2976 ( .A1(n2710), .A2(n2709), .A3(n2708), .A4(n2707), .Y(n2716)
         );
  AO22X1_RVT U2977 ( .A1(\inq_ary[6][99] ), .A2(n3311), .A3(\inq_ary[2][99] ), 
        .A4(n3271), .Y(n2714) );
  AO22X1_RVT U2978 ( .A1(\inq_ary[11][99] ), .A2(n3316), .A3(\inq_ary[12][99] ), .A4(n3303), .Y(n2713) );
  AO22X1_RVT U2979 ( .A1(\inq_ary[1][99] ), .A2(n3324), .A3(\inq_ary[14][99] ), 
        .A4(n3325), .Y(n2712) );
  AO22X1_RVT U2980 ( .A1(\inq_ary[7][99] ), .A2(n3322), .A3(\inq_ary[13][99] ), 
        .A4(n3323), .Y(n2711) );
  NOR4X1_RVT U2981 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .Y(n2715)
         );
  NAND2X0_RVT U2982 ( .A1(n2716), .A2(n2715), .Y(N361) );
  AO22X1_RVT U2983 ( .A1(\inq_ary[8][100] ), .A2(n3313), .A3(
        \inq_ary[14][100] ), .A4(n3325), .Y(n2720) );
  AO22X1_RVT U2984 ( .A1(\inq_ary[3][100] ), .A2(n3310), .A3(
        \inq_ary[10][100] ), .A4(n3326), .Y(n2719) );
  AO22X1_RVT U2985 ( .A1(\inq_ary[9][100] ), .A2(n3314), .A3(\inq_ary[7][100] ), .A4(n3322), .Y(n2718) );
  AO22X1_RVT U2986 ( .A1(\inq_ary[12][100] ), .A2(n3303), .A3(
        \inq_ary[0][100] ), .A4(n3315), .Y(n2717) );
  NOR4X1_RVT U2987 ( .A1(n2720), .A2(n2719), .A3(n2718), .A4(n2717), .Y(n2726)
         );
  AO22X1_RVT U2988 ( .A1(\inq_ary[2][100] ), .A2(n3271), .A3(
        \inq_ary[15][100] ), .A4(n3312), .Y(n2724) );
  AO22X1_RVT U2989 ( .A1(\inq_ary[11][100] ), .A2(n3316), .A3(
        \inq_ary[4][100] ), .A4(n3321), .Y(n2723) );
  AO22X1_RVT U2990 ( .A1(\inq_ary[1][100] ), .A2(n3324), .A3(\inq_ary[5][100] ), .A4(n3298), .Y(n2722) );
  AO22X1_RVT U2991 ( .A1(\inq_ary[6][100] ), .A2(n3311), .A3(
        \inq_ary[13][100] ), .A4(n3323), .Y(n2721) );
  NOR4X1_RVT U2992 ( .A1(n2724), .A2(n2723), .A3(n2722), .A4(n2721), .Y(n2725)
         );
  NAND2X0_RVT U2993 ( .A1(n2726), .A2(n2725), .Y(N362) );
  AO22X1_RVT U2994 ( .A1(\inq_ary[14][101] ), .A2(n3325), .A3(
        \inq_ary[8][101] ), .A4(n3313), .Y(n2730) );
  AO22X1_RVT U2995 ( .A1(\inq_ary[10][101] ), .A2(n3326), .A3(
        \inq_ary[9][101] ), .A4(n3314), .Y(n2729) );
  AO22X1_RVT U2996 ( .A1(\inq_ary[13][101] ), .A2(n3323), .A3(
        \inq_ary[1][101] ), .A4(n3324), .Y(n2728) );
  AO22X1_RVT U2997 ( .A1(\inq_ary[11][101] ), .A2(n3316), .A3(
        \inq_ary[2][101] ), .A4(n3271), .Y(n2727) );
  NOR4X1_RVT U2998 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .Y(n2736)
         );
  AO22X1_RVT U2999 ( .A1(\inq_ary[3][101] ), .A2(n3310), .A3(
        \inq_ary[15][101] ), .A4(n3312), .Y(n2734) );
  AO22X1_RVT U3000 ( .A1(\inq_ary[6][101] ), .A2(n3311), .A3(\inq_ary[7][101] ), .A4(n3322), .Y(n2733) );
  AO22X1_RVT U3001 ( .A1(\inq_ary[12][101] ), .A2(n3303), .A3(
        \inq_ary[5][101] ), .A4(n3298), .Y(n2732) );
  AO22X1_RVT U3002 ( .A1(\inq_ary[4][101] ), .A2(n3321), .A3(\inq_ary[0][101] ), .A4(n3315), .Y(n2731) );
  NOR4X1_RVT U3003 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .Y(n2735)
         );
  NAND2X0_RVT U3004 ( .A1(n2736), .A2(n2735), .Y(N363) );
  AO22X1_RVT U3005 ( .A1(\inq_ary[1][102] ), .A2(n3324), .A3(\inq_ary[0][102] ), .A4(n3315), .Y(n2740) );
  AO22X1_RVT U3006 ( .A1(\inq_ary[8][102] ), .A2(n3313), .A3(\inq_ary[6][102] ), .A4(n3311), .Y(n2739) );
  AO22X1_RVT U3007 ( .A1(\inq_ary[14][102] ), .A2(n3325), .A3(
        \inq_ary[2][102] ), .A4(n3271), .Y(n2738) );
  AO22X1_RVT U3008 ( .A1(\inq_ary[3][102] ), .A2(n3310), .A3(
        \inq_ary[10][102] ), .A4(n3326), .Y(n2737) );
  NOR4X1_RVT U3009 ( .A1(n2740), .A2(n2739), .A3(n2738), .A4(n2737), .Y(n2746)
         );
  AO22X1_RVT U3010 ( .A1(\inq_ary[9][102] ), .A2(n3314), .A3(
        \inq_ary[13][102] ), .A4(n3323), .Y(n2744) );
  AO22X1_RVT U3011 ( .A1(\inq_ary[4][102] ), .A2(n3321), .A3(\inq_ary[7][102] ), .A4(n3322), .Y(n2743) );
  AO22X1_RVT U3012 ( .A1(\inq_ary[11][102] ), .A2(n3316), .A3(
        \inq_ary[12][102] ), .A4(n3303), .Y(n2742) );
  AO22X1_RVT U3013 ( .A1(\inq_ary[15][102] ), .A2(n3312), .A3(
        \inq_ary[5][102] ), .A4(n3298), .Y(n2741) );
  NOR4X1_RVT U3014 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .Y(n2745)
         );
  NAND2X0_RVT U3015 ( .A1(n2746), .A2(n2745), .Y(N364) );
  AO22X1_RVT U3016 ( .A1(\inq_ary[11][103] ), .A2(n3316), .A3(
        \inq_ary[13][103] ), .A4(n3323), .Y(n2750) );
  AO22X1_RVT U3017 ( .A1(\inq_ary[15][103] ), .A2(n3312), .A3(
        \inq_ary[6][103] ), .A4(n3311), .Y(n2749) );
  AO22X1_RVT U3018 ( .A1(\inq_ary[12][103] ), .A2(n3303), .A3(
        \inq_ary[2][103] ), .A4(n3271), .Y(n2748) );
  AO22X1_RVT U3019 ( .A1(\inq_ary[9][103] ), .A2(n3314), .A3(\inq_ary[3][103] ), .A4(n3310), .Y(n2747) );
  NOR4X1_RVT U3020 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .Y(n2756)
         );
  AO22X1_RVT U3021 ( .A1(\inq_ary[1][103] ), .A2(n3324), .A3(\inq_ary[8][103] ), .A4(n3313), .Y(n2754) );
  AO22X1_RVT U3022 ( .A1(\inq_ary[0][103] ), .A2(n3315), .A3(
        \inq_ary[14][103] ), .A4(n3325), .Y(n2753) );
  AO22X1_RVT U3023 ( .A1(\inq_ary[4][103] ), .A2(n3321), .A3(
        \inq_ary[10][103] ), .A4(n3326), .Y(n2752) );
  AO22X1_RVT U3024 ( .A1(\inq_ary[7][103] ), .A2(n3322), .A3(\inq_ary[5][103] ), .A4(n3298), .Y(n2751) );
  NOR4X1_RVT U3025 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), .Y(n2755)
         );
  NAND2X0_RVT U3026 ( .A1(n2756), .A2(n2755), .Y(N365) );
  AO22X1_RVT U3027 ( .A1(\inq_ary[3][104] ), .A2(n3310), .A3(
        \inq_ary[14][104] ), .A4(n3325), .Y(n2760) );
  AO22X1_RVT U3028 ( .A1(\inq_ary[2][104] ), .A2(n3271), .A3(
        \inq_ary[15][104] ), .A4(n3312), .Y(n2759) );
  AO22X1_RVT U3029 ( .A1(\inq_ary[12][104] ), .A2(n3303), .A3(
        \inq_ary[7][104] ), .A4(n3322), .Y(n2758) );
  AO22X1_RVT U3030 ( .A1(\inq_ary[9][104] ), .A2(n3314), .A3(\inq_ary[1][104] ), .A4(n3324), .Y(n2757) );
  NOR4X1_RVT U3031 ( .A1(n2760), .A2(n2759), .A3(n2758), .A4(n2757), .Y(n2766)
         );
  AO22X1_RVT U3032 ( .A1(\inq_ary[8][104] ), .A2(n3313), .A3(\inq_ary[0][104] ), .A4(n3315), .Y(n2764) );
  AO22X1_RVT U3033 ( .A1(\inq_ary[11][104] ), .A2(n3316), .A3(
        \inq_ary[5][104] ), .A4(n3298), .Y(n2763) );
  AO22X1_RVT U3034 ( .A1(\inq_ary[10][104] ), .A2(n3326), .A3(
        \inq_ary[6][104] ), .A4(n3311), .Y(n2762) );
  AO22X1_RVT U3035 ( .A1(\inq_ary[13][104] ), .A2(n3323), .A3(
        \inq_ary[4][104] ), .A4(n3321), .Y(n2761) );
  NOR4X1_RVT U3036 ( .A1(n2764), .A2(n2763), .A3(n2762), .A4(n2761), .Y(n2765)
         );
  NAND2X0_RVT U3037 ( .A1(n2766), .A2(n2765), .Y(N366) );
  AO22X1_RVT U3038 ( .A1(\inq_ary[3][105] ), .A2(n3310), .A3(\inq_ary[9][105] ), .A4(n3314), .Y(n2770) );
  AO22X1_RVT U3039 ( .A1(\inq_ary[7][105] ), .A2(n3322), .A3(\inq_ary[0][105] ), .A4(n3315), .Y(n2769) );
  AO22X1_RVT U3040 ( .A1(\inq_ary[6][105] ), .A2(n3311), .A3(
        \inq_ary[11][105] ), .A4(n3316), .Y(n2768) );
  AO22X1_RVT U3041 ( .A1(\inq_ary[12][105] ), .A2(n3303), .A3(
        \inq_ary[8][105] ), .A4(n3313), .Y(n2767) );
  NOR4X1_RVT U3042 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), .Y(n2776)
         );
  AO22X1_RVT U3043 ( .A1(\inq_ary[14][105] ), .A2(n3325), .A3(
        \inq_ary[10][105] ), .A4(n3326), .Y(n2774) );
  AO22X1_RVT U3044 ( .A1(\inq_ary[15][105] ), .A2(n3312), .A3(
        \inq_ary[5][105] ), .A4(n3298), .Y(n2773) );
  AO22X1_RVT U3045 ( .A1(\inq_ary[13][105] ), .A2(n3323), .A3(
        \inq_ary[1][105] ), .A4(n3324), .Y(n2772) );
  AO22X1_RVT U3046 ( .A1(\inq_ary[4][105] ), .A2(n3321), .A3(\inq_ary[2][105] ), .A4(n3271), .Y(n2771) );
  NOR4X1_RVT U3047 ( .A1(n2774), .A2(n2773), .A3(n2772), .A4(n2771), .Y(n2775)
         );
  NAND2X0_RVT U3048 ( .A1(n2776), .A2(n2775), .Y(N367) );
  AO22X1_RVT U3049 ( .A1(\inq_ary[0][106] ), .A2(n3315), .A3(\inq_ary[6][106] ), .A4(n3311), .Y(n2780) );
  AO22X1_RVT U3050 ( .A1(\inq_ary[2][106] ), .A2(n3271), .A3(
        \inq_ary[11][106] ), .A4(n3316), .Y(n2779) );
  AO22X1_RVT U3051 ( .A1(\inq_ary[1][106] ), .A2(n3324), .A3(\inq_ary[5][106] ), .A4(n3298), .Y(n2778) );
  AO22X1_RVT U3052 ( .A1(\inq_ary[9][106] ), .A2(n3314), .A3(\inq_ary[3][106] ), .A4(n3310), .Y(n2777) );
  NOR4X1_RVT U3053 ( .A1(n2780), .A2(n2779), .A3(n2778), .A4(n2777), .Y(n2786)
         );
  AO22X1_RVT U3054 ( .A1(\inq_ary[14][106] ), .A2(n3325), .A3(
        \inq_ary[12][106] ), .A4(n3303), .Y(n2784) );
  AO22X1_RVT U3055 ( .A1(\inq_ary[13][106] ), .A2(n3323), .A3(
        \inq_ary[7][106] ), .A4(n3322), .Y(n2783) );
  AO22X1_RVT U3056 ( .A1(\inq_ary[15][106] ), .A2(n3312), .A3(
        \inq_ary[8][106] ), .A4(n3313), .Y(n2782) );
  AO22X1_RVT U3057 ( .A1(\inq_ary[4][106] ), .A2(n3321), .A3(
        \inq_ary[10][106] ), .A4(n3326), .Y(n2781) );
  NOR4X1_RVT U3058 ( .A1(n2784), .A2(n2783), .A3(n2782), .A4(n2781), .Y(n2785)
         );
  NAND2X0_RVT U3059 ( .A1(n2786), .A2(n2785), .Y(N368) );
  AO22X1_RVT U3060 ( .A1(\inq_ary[9][107] ), .A2(n3314), .A3(\inq_ary[4][107] ), .A4(n3321), .Y(n2790) );
  AO22X1_RVT U3061 ( .A1(\inq_ary[2][107] ), .A2(n3271), .A3(\inq_ary[0][107] ), .A4(n3315), .Y(n2789) );
  AO22X1_RVT U3062 ( .A1(\inq_ary[10][107] ), .A2(n3326), .A3(
        \inq_ary[8][107] ), .A4(n3313), .Y(n2788) );
  AO22X1_RVT U3063 ( .A1(\inq_ary[14][107] ), .A2(n3325), .A3(
        \inq_ary[12][107] ), .A4(n3303), .Y(n2787) );
  NOR4X1_RVT U3064 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .Y(n2796)
         );
  AO22X1_RVT U3065 ( .A1(\inq_ary[7][107] ), .A2(n3322), .A3(
        \inq_ary[13][107] ), .A4(n3323), .Y(n2794) );
  AO22X1_RVT U3066 ( .A1(\inq_ary[1][107] ), .A2(n3324), .A3(
        \inq_ary[15][107] ), .A4(n3312), .Y(n2793) );
  AO22X1_RVT U3067 ( .A1(\inq_ary[5][107] ), .A2(n3298), .A3(\inq_ary[3][107] ), .A4(n3310), .Y(n2792) );
  AO22X1_RVT U3068 ( .A1(\inq_ary[6][107] ), .A2(n3311), .A3(
        \inq_ary[11][107] ), .A4(n3316), .Y(n2791) );
  NOR4X1_RVT U3069 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), .Y(n2795)
         );
  NAND2X0_RVT U3070 ( .A1(n2796), .A2(n2795), .Y(N369) );
  AO22X1_RVT U3071 ( .A1(\inq_ary[11][108] ), .A2(n3316), .A3(
        \inq_ary[6][108] ), .A4(n3311), .Y(n2800) );
  AO22X1_RVT U3072 ( .A1(\inq_ary[13][108] ), .A2(n3323), .A3(
        \inq_ary[5][108] ), .A4(n3298), .Y(n2799) );
  AO22X1_RVT U3073 ( .A1(\inq_ary[2][108] ), .A2(n3271), .A3(
        \inq_ary[14][108] ), .A4(n3325), .Y(n2798) );
  AO22X1_RVT U3074 ( .A1(\inq_ary[15][108] ), .A2(n3312), .A3(
        \inq_ary[10][108] ), .A4(n3326), .Y(n2797) );
  NOR4X1_RVT U3075 ( .A1(n2800), .A2(n2799), .A3(n2798), .A4(n2797), .Y(n2806)
         );
  AO22X1_RVT U3076 ( .A1(\inq_ary[8][108] ), .A2(n3313), .A3(\inq_ary[9][108] ), .A4(n3314), .Y(n2804) );
  AO22X1_RVT U3077 ( .A1(\inq_ary[4][108] ), .A2(n3321), .A3(\inq_ary[1][108] ), .A4(n3324), .Y(n2803) );
  AO22X1_RVT U3078 ( .A1(\inq_ary[0][108] ), .A2(n3315), .A3(\inq_ary[3][108] ), .A4(n3310), .Y(n2802) );
  AO22X1_RVT U3079 ( .A1(\inq_ary[7][108] ), .A2(n3322), .A3(
        \inq_ary[12][108] ), .A4(n3303), .Y(n2801) );
  NOR4X1_RVT U3080 ( .A1(n2804), .A2(n2803), .A3(n2802), .A4(n2801), .Y(n2805)
         );
  NAND2X0_RVT U3081 ( .A1(n2806), .A2(n2805), .Y(N370) );
  AO22X1_RVT U3082 ( .A1(\inq_ary[1][109] ), .A2(n3324), .A3(\inq_ary[9][109] ), .A4(n3314), .Y(n2810) );
  AO22X1_RVT U3083 ( .A1(\inq_ary[0][109] ), .A2(n3315), .A3(
        \inq_ary[10][109] ), .A4(n3326), .Y(n2809) );
  AO22X1_RVT U3084 ( .A1(\inq_ary[13][109] ), .A2(n3323), .A3(
        \inq_ary[8][109] ), .A4(n3313), .Y(n2808) );
  AO22X1_RVT U3085 ( .A1(\inq_ary[14][109] ), .A2(n3325), .A3(
        \inq_ary[3][109] ), .A4(n3310), .Y(n2807) );
  NOR4X1_RVT U3086 ( .A1(n2810), .A2(n2809), .A3(n2808), .A4(n2807), .Y(n2816)
         );
  AO22X1_RVT U3087 ( .A1(\inq_ary[4][109] ), .A2(n3321), .A3(\inq_ary[5][109] ), .A4(n3298), .Y(n2814) );
  AO22X1_RVT U3088 ( .A1(\inq_ary[12][109] ), .A2(n3303), .A3(
        \inq_ary[7][109] ), .A4(n3322), .Y(n2813) );
  AO22X1_RVT U3089 ( .A1(\inq_ary[6][109] ), .A2(n3311), .A3(\inq_ary[2][109] ), .A4(n3271), .Y(n2812) );
  AO22X1_RVT U3090 ( .A1(\inq_ary[11][109] ), .A2(n3316), .A3(
        \inq_ary[15][109] ), .A4(n3312), .Y(n2811) );
  NOR4X1_RVT U3091 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .Y(n2815)
         );
  NAND2X0_RVT U3092 ( .A1(n2816), .A2(n2815), .Y(N371) );
  AO22X1_RVT U3093 ( .A1(\inq_ary[1][110] ), .A2(n3324), .A3(
        \inq_ary[12][110] ), .A4(n3303), .Y(n2820) );
  AO22X1_RVT U3094 ( .A1(\inq_ary[5][110] ), .A2(n3298), .A3(
        \inq_ary[13][110] ), .A4(n3323), .Y(n2819) );
  AO22X1_RVT U3095 ( .A1(\inq_ary[15][110] ), .A2(n3312), .A3(
        \inq_ary[14][110] ), .A4(n3325), .Y(n2818) );
  AO22X1_RVT U3096 ( .A1(\inq_ary[11][110] ), .A2(n3316), .A3(
        \inq_ary[2][110] ), .A4(n3271), .Y(n2817) );
  NOR4X1_RVT U3097 ( .A1(n2820), .A2(n2819), .A3(n2818), .A4(n2817), .Y(n2826)
         );
  AO22X1_RVT U3098 ( .A1(\inq_ary[9][110] ), .A2(n3314), .A3(\inq_ary[4][110] ), .A4(n3321), .Y(n2824) );
  AO22X1_RVT U3099 ( .A1(\inq_ary[6][110] ), .A2(n3311), .A3(\inq_ary[8][110] ), .A4(n3313), .Y(n2823) );
  AO22X1_RVT U3100 ( .A1(\inq_ary[3][110] ), .A2(n3310), .A3(\inq_ary[7][110] ), .A4(n3322), .Y(n2822) );
  AO22X1_RVT U3101 ( .A1(\inq_ary[10][110] ), .A2(n3326), .A3(
        \inq_ary[0][110] ), .A4(n3315), .Y(n2821) );
  NOR4X1_RVT U3102 ( .A1(n2824), .A2(n2823), .A3(n2822), .A4(n2821), .Y(n2825)
         );
  NAND2X0_RVT U3103 ( .A1(n2826), .A2(n2825), .Y(N372) );
  AO22X1_RVT U3104 ( .A1(\inq_ary[3][111] ), .A2(n3310), .A3(\inq_ary[1][111] ), .A4(n3324), .Y(n2830) );
  AO22X1_RVT U3105 ( .A1(\inq_ary[4][111] ), .A2(n3321), .A3(\inq_ary[9][111] ), .A4(n3314), .Y(n2829) );
  AO22X1_RVT U3106 ( .A1(\inq_ary[5][111] ), .A2(n3298), .A3(
        \inq_ary[15][111] ), .A4(n3312), .Y(n2828) );
  AO22X1_RVT U3107 ( .A1(\inq_ary[7][111] ), .A2(n3322), .A3(
        \inq_ary[14][111] ), .A4(n3325), .Y(n2827) );
  NOR4X1_RVT U3108 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .Y(n2836)
         );
  AO22X1_RVT U3109 ( .A1(\inq_ary[0][111] ), .A2(n3315), .A3(\inq_ary[8][111] ), .A4(n3313), .Y(n2834) );
  AO22X1_RVT U3110 ( .A1(\inq_ary[10][111] ), .A2(n3326), .A3(
        \inq_ary[13][111] ), .A4(n3323), .Y(n2833) );
  AO22X1_RVT U3111 ( .A1(\inq_ary[12][111] ), .A2(n3303), .A3(
        \inq_ary[2][111] ), .A4(n3271), .Y(n2832) );
  AO22X1_RVT U3112 ( .A1(\inq_ary[6][111] ), .A2(n3311), .A3(
        \inq_ary[11][111] ), .A4(n3316), .Y(n2831) );
  NOR4X1_RVT U3113 ( .A1(n2834), .A2(n2833), .A3(n2832), .A4(n2831), .Y(n2835)
         );
  NAND2X0_RVT U3114 ( .A1(n2836), .A2(n2835), .Y(N373) );
  AO22X1_RVT U3115 ( .A1(\inq_ary[13][112] ), .A2(n3323), .A3(
        \inq_ary[3][112] ), .A4(n3310), .Y(n2840) );
  AO22X1_RVT U3116 ( .A1(\inq_ary[11][112] ), .A2(n3316), .A3(
        \inq_ary[8][112] ), .A4(n3313), .Y(n2839) );
  AO22X1_RVT U3117 ( .A1(\inq_ary[10][112] ), .A2(n3326), .A3(
        \inq_ary[6][112] ), .A4(n3311), .Y(n2838) );
  AO22X1_RVT U3118 ( .A1(\inq_ary[0][112] ), .A2(n3315), .A3(\inq_ary[4][112] ), .A4(n3321), .Y(n2837) );
  NOR4X1_RVT U3119 ( .A1(n2840), .A2(n2839), .A3(n2838), .A4(n2837), .Y(n2846)
         );
  AO22X1_RVT U3120 ( .A1(\inq_ary[14][112] ), .A2(n3325), .A3(
        \inq_ary[9][112] ), .A4(n3314), .Y(n2844) );
  AO22X1_RVT U3121 ( .A1(\inq_ary[15][112] ), .A2(n3312), .A3(
        \inq_ary[1][112] ), .A4(n3324), .Y(n2843) );
  AO22X1_RVT U3122 ( .A1(\inq_ary[7][112] ), .A2(n3322), .A3(
        \inq_ary[12][112] ), .A4(n3303), .Y(n2842) );
  AO22X1_RVT U3123 ( .A1(\inq_ary[2][112] ), .A2(n3271), .A3(\inq_ary[5][112] ), .A4(n3298), .Y(n2841) );
  NOR4X1_RVT U3124 ( .A1(n2844), .A2(n2843), .A3(n2842), .A4(n2841), .Y(n2845)
         );
  NAND2X0_RVT U3125 ( .A1(n2846), .A2(n2845), .Y(N374) );
  AO22X1_RVT U3126 ( .A1(\inq_ary[15][113] ), .A2(n3312), .A3(
        \inq_ary[9][113] ), .A4(n3314), .Y(n2850) );
  AO22X1_RVT U3127 ( .A1(\inq_ary[7][113] ), .A2(n3322), .A3(\inq_ary[3][113] ), .A4(n3310), .Y(n2849) );
  AO22X1_RVT U3128 ( .A1(\inq_ary[8][113] ), .A2(n3313), .A3(\inq_ary[4][113] ), .A4(n3321), .Y(n2848) );
  AO22X1_RVT U3129 ( .A1(\inq_ary[10][113] ), .A2(n3326), .A3(
        \inq_ary[12][113] ), .A4(n3303), .Y(n2847) );
  NOR4X1_RVT U3130 ( .A1(n2850), .A2(n2849), .A3(n2848), .A4(n2847), .Y(n2856)
         );
  AO22X1_RVT U3131 ( .A1(\inq_ary[2][113] ), .A2(n3271), .A3(\inq_ary[0][113] ), .A4(n3315), .Y(n2854) );
  AO22X1_RVT U3132 ( .A1(\inq_ary[13][113] ), .A2(n3323), .A3(
        \inq_ary[5][113] ), .A4(n3298), .Y(n2853) );
  AO22X1_RVT U3133 ( .A1(\inq_ary[14][113] ), .A2(n3325), .A3(
        \inq_ary[11][113] ), .A4(n3316), .Y(n2852) );
  AO22X1_RVT U3134 ( .A1(\inq_ary[1][113] ), .A2(n3324), .A3(\inq_ary[6][113] ), .A4(n3311), .Y(n2851) );
  NOR4X1_RVT U3135 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), .Y(n2855)
         );
  NAND2X0_RVT U3136 ( .A1(n2856), .A2(n2855), .Y(N375) );
  AO22X1_RVT U3137 ( .A1(\inq_ary[2][114] ), .A2(n3271), .A3(\inq_ary[5][114] ), .A4(n3298), .Y(n2860) );
  AO22X1_RVT U3138 ( .A1(\inq_ary[9][114] ), .A2(n3314), .A3(\inq_ary[1][114] ), .A4(n3324), .Y(n2859) );
  AO22X1_RVT U3139 ( .A1(\inq_ary[4][114] ), .A2(n3321), .A3(
        \inq_ary[13][114] ), .A4(n3323), .Y(n2858) );
  AO22X1_RVT U3140 ( .A1(\inq_ary[14][114] ), .A2(n3325), .A3(
        \inq_ary[7][114] ), .A4(n3322), .Y(n2857) );
  NOR4X1_RVT U3141 ( .A1(n2860), .A2(n2859), .A3(n2858), .A4(n2857), .Y(n2866)
         );
  AO22X1_RVT U3142 ( .A1(\inq_ary[15][114] ), .A2(n3312), .A3(
        \inq_ary[0][114] ), .A4(n3315), .Y(n2864) );
  AO22X1_RVT U3143 ( .A1(\inq_ary[8][114] ), .A2(n3313), .A3(
        \inq_ary[12][114] ), .A4(n3303), .Y(n2863) );
  AO22X1_RVT U3144 ( .A1(\inq_ary[3][114] ), .A2(n3310), .A3(
        \inq_ary[11][114] ), .A4(n3316), .Y(n2862) );
  AO22X1_RVT U3145 ( .A1(\inq_ary[6][114] ), .A2(n3311), .A3(
        \inq_ary[10][114] ), .A4(n3326), .Y(n2861) );
  NOR4X1_RVT U3146 ( .A1(n2864), .A2(n2863), .A3(n2862), .A4(n2861), .Y(n2865)
         );
  NAND2X0_RVT U3147 ( .A1(n2866), .A2(n2865), .Y(N376) );
  AO22X1_RVT U3148 ( .A1(\inq_ary[8][115] ), .A2(n3313), .A3(\inq_ary[5][115] ), .A4(n3298), .Y(n2870) );
  AO22X1_RVT U3149 ( .A1(\inq_ary[9][115] ), .A2(n3314), .A3(\inq_ary[2][115] ), .A4(n3271), .Y(n2869) );
  AO22X1_RVT U3150 ( .A1(\inq_ary[14][115] ), .A2(n3325), .A3(
        \inq_ary[4][115] ), .A4(n3321), .Y(n2868) );
  AO22X1_RVT U3151 ( .A1(\inq_ary[7][115] ), .A2(n3322), .A3(
        \inq_ary[10][115] ), .A4(n3326), .Y(n2867) );
  NOR4X1_RVT U3152 ( .A1(n2870), .A2(n2869), .A3(n2868), .A4(n2867), .Y(n2876)
         );
  AO22X1_RVT U3153 ( .A1(\inq_ary[1][115] ), .A2(n3324), .A3(\inq_ary[3][115] ), .A4(n3310), .Y(n2874) );
  AO22X1_RVT U3154 ( .A1(\inq_ary[11][115] ), .A2(n3316), .A3(
        \inq_ary[12][115] ), .A4(n3303), .Y(n2873) );
  AO22X1_RVT U3155 ( .A1(\inq_ary[15][115] ), .A2(n3312), .A3(
        \inq_ary[0][115] ), .A4(n3315), .Y(n2872) );
  AO22X1_RVT U3156 ( .A1(\inq_ary[6][115] ), .A2(n3311), .A3(
        \inq_ary[13][115] ), .A4(n3323), .Y(n2871) );
  NOR4X1_RVT U3157 ( .A1(n2874), .A2(n2873), .A3(n2872), .A4(n2871), .Y(n2875)
         );
  NAND2X0_RVT U3158 ( .A1(n2876), .A2(n2875), .Y(N377) );
  AO22X1_RVT U3159 ( .A1(\inq_ary[8][116] ), .A2(n3313), .A3(
        \inq_ary[14][116] ), .A4(n3325), .Y(n2880) );
  AO22X1_RVT U3160 ( .A1(\inq_ary[12][116] ), .A2(n3303), .A3(
        \inq_ary[9][116] ), .A4(n3314), .Y(n2879) );
  AO22X1_RVT U3161 ( .A1(\inq_ary[11][116] ), .A2(n3316), .A3(
        \inq_ary[1][116] ), .A4(n3324), .Y(n2878) );
  AO22X1_RVT U3162 ( .A1(\inq_ary[10][116] ), .A2(n3326), .A3(
        \inq_ary[13][116] ), .A4(n3323), .Y(n2877) );
  NOR4X1_RVT U3163 ( .A1(n2880), .A2(n2879), .A3(n2878), .A4(n2877), .Y(n2886)
         );
  AO22X1_RVT U3164 ( .A1(\inq_ary[3][116] ), .A2(n3310), .A3(\inq_ary[4][116] ), .A4(n3321), .Y(n2884) );
  AO22X1_RVT U3165 ( .A1(\inq_ary[15][116] ), .A2(n3312), .A3(
        \inq_ary[5][116] ), .A4(n3298), .Y(n2883) );
  AO22X1_RVT U3166 ( .A1(\inq_ary[6][116] ), .A2(n3311), .A3(\inq_ary[0][116] ), .A4(n3315), .Y(n2882) );
  AO22X1_RVT U3167 ( .A1(\inq_ary[2][116] ), .A2(n3271), .A3(\inq_ary[7][116] ), .A4(n3322), .Y(n2881) );
  NOR4X1_RVT U3168 ( .A1(n2884), .A2(n2883), .A3(n2882), .A4(n2881), .Y(n2885)
         );
  NAND2X0_RVT U3169 ( .A1(n2886), .A2(n2885), .Y(N378) );
  AO22X1_RVT U3170 ( .A1(\inq_ary[14][117] ), .A2(n3325), .A3(
        \inq_ary[15][117] ), .A4(n3312), .Y(n2890) );
  AO22X1_RVT U3171 ( .A1(\inq_ary[11][117] ), .A2(n3316), .A3(
        \inq_ary[1][117] ), .A4(n3324), .Y(n2889) );
  AO22X1_RVT U3172 ( .A1(\inq_ary[8][117] ), .A2(n3313), .A3(\inq_ary[2][117] ), .A4(n3271), .Y(n2888) );
  AO22X1_RVT U3173 ( .A1(\inq_ary[4][117] ), .A2(n3321), .A3(\inq_ary[6][117] ), .A4(n3311), .Y(n2887) );
  NOR4X1_RVT U3174 ( .A1(n2890), .A2(n2889), .A3(n2888), .A4(n2887), .Y(n2896)
         );
  AO22X1_RVT U3175 ( .A1(\inq_ary[0][117] ), .A2(n3315), .A3(\inq_ary[9][117] ), .A4(n3314), .Y(n2894) );
  AO22X1_RVT U3176 ( .A1(\inq_ary[10][117] ), .A2(n3326), .A3(
        \inq_ary[12][117] ), .A4(n3303), .Y(n2893) );
  AO22X1_RVT U3177 ( .A1(\inq_ary[7][117] ), .A2(n3322), .A3(\inq_ary[5][117] ), .A4(n3298), .Y(n2892) );
  AO22X1_RVT U3178 ( .A1(\inq_ary[3][117] ), .A2(n3310), .A3(
        \inq_ary[13][117] ), .A4(n3323), .Y(n2891) );
  NOR4X1_RVT U3179 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .Y(n2895)
         );
  NAND2X0_RVT U3180 ( .A1(n2896), .A2(n2895), .Y(N379) );
  AO22X1_RVT U3181 ( .A1(\inq_ary[1][118] ), .A2(n3324), .A3(
        \inq_ary[14][118] ), .A4(n3325), .Y(n2900) );
  AO22X1_RVT U3182 ( .A1(\inq_ary[15][118] ), .A2(n3312), .A3(
        \inq_ary[4][118] ), .A4(n3321), .Y(n2899) );
  AO22X1_RVT U3183 ( .A1(\inq_ary[8][118] ), .A2(n3313), .A3(\inq_ary[5][118] ), .A4(n3298), .Y(n2898) );
  AO22X1_RVT U3184 ( .A1(\inq_ary[6][118] ), .A2(n3311), .A3(\inq_ary[9][118] ), .A4(n3314), .Y(n2897) );
  NOR4X1_RVT U3185 ( .A1(n2900), .A2(n2899), .A3(n2898), .A4(n2897), .Y(n2906)
         );
  AO22X1_RVT U3186 ( .A1(\inq_ary[10][118] ), .A2(n3326), .A3(
        \inq_ary[7][118] ), .A4(n3322), .Y(n2904) );
  AO22X1_RVT U3187 ( .A1(\inq_ary[11][118] ), .A2(n3316), .A3(
        \inq_ary[13][118] ), .A4(n3323), .Y(n2903) );
  AO22X1_RVT U3188 ( .A1(\inq_ary[0][118] ), .A2(n3315), .A3(\inq_ary[3][118] ), .A4(n3310), .Y(n2902) );
  AO22X1_RVT U3189 ( .A1(\inq_ary[2][118] ), .A2(n3271), .A3(
        \inq_ary[12][118] ), .A4(n3303), .Y(n2901) );
  NOR4X1_RVT U3190 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .Y(n2905)
         );
  NAND2X0_RVT U3191 ( .A1(n2906), .A2(n2905), .Y(N380) );
  AO22X1_RVT U3192 ( .A1(\inq_ary[9][119] ), .A2(n3314), .A3(
        \inq_ary[10][119] ), .A4(n3326), .Y(n2910) );
  AO22X1_RVT U3193 ( .A1(\inq_ary[7][119] ), .A2(n3322), .A3(
        \inq_ary[13][119] ), .A4(n3323), .Y(n2909) );
  AO22X1_RVT U3194 ( .A1(\inq_ary[8][119] ), .A2(n3313), .A3(
        \inq_ary[12][119] ), .A4(n3303), .Y(n2908) );
  AO22X1_RVT U3195 ( .A1(\inq_ary[0][119] ), .A2(n3315), .A3(
        \inq_ary[14][119] ), .A4(n3325), .Y(n2907) );
  NOR4X1_RVT U3196 ( .A1(n2910), .A2(n2909), .A3(n2908), .A4(n2907), .Y(n2916)
         );
  AO22X1_RVT U3197 ( .A1(\inq_ary[3][119] ), .A2(n3310), .A3(\inq_ary[1][119] ), .A4(n3324), .Y(n2914) );
  AO22X1_RVT U3198 ( .A1(\inq_ary[6][119] ), .A2(n3311), .A3(\inq_ary[4][119] ), .A4(n3321), .Y(n2913) );
  AO22X1_RVT U3199 ( .A1(\inq_ary[15][119] ), .A2(n3312), .A3(
        \inq_ary[2][119] ), .A4(n3271), .Y(n2912) );
  AO22X1_RVT U3200 ( .A1(\inq_ary[5][119] ), .A2(n3298), .A3(
        \inq_ary[11][119] ), .A4(n3316), .Y(n2911) );
  NOR4X1_RVT U3201 ( .A1(n2914), .A2(n2913), .A3(n2912), .A4(n2911), .Y(n2915)
         );
  NAND2X0_RVT U3202 ( .A1(n2916), .A2(n2915), .Y(N381) );
  AO22X1_RVT U3203 ( .A1(\inq_ary[1][120] ), .A2(n3324), .A3(\inq_ary[8][120] ), .A4(n3313), .Y(n2920) );
  AO22X1_RVT U3204 ( .A1(\inq_ary[9][120] ), .A2(n3314), .A3(\inq_ary[7][120] ), .A4(n3322), .Y(n2919) );
  AO22X1_RVT U3205 ( .A1(\inq_ary[5][120] ), .A2(n3298), .A3(
        \inq_ary[15][120] ), .A4(n3312), .Y(n2918) );
  AO22X1_RVT U3206 ( .A1(\inq_ary[4][120] ), .A2(n3321), .A3(\inq_ary[6][120] ), .A4(n3311), .Y(n2917) );
  NOR4X1_RVT U3207 ( .A1(n2920), .A2(n2919), .A3(n2918), .A4(n2917), .Y(n2926)
         );
  AO22X1_RVT U3208 ( .A1(\inq_ary[10][120] ), .A2(n3326), .A3(
        \inq_ary[2][120] ), .A4(n3271), .Y(n2924) );
  AO22X1_RVT U3209 ( .A1(\inq_ary[3][120] ), .A2(n3310), .A3(
        \inq_ary[11][120] ), .A4(n3316), .Y(n2923) );
  AO22X1_RVT U3210 ( .A1(\inq_ary[0][120] ), .A2(n3315), .A3(
        \inq_ary[13][120] ), .A4(n3323), .Y(n2922) );
  AO22X1_RVT U3211 ( .A1(\inq_ary[14][120] ), .A2(n3325), .A3(
        \inq_ary[12][120] ), .A4(n3303), .Y(n2921) );
  NOR4X1_RVT U3212 ( .A1(n2924), .A2(n2923), .A3(n2922), .A4(n2921), .Y(n2925)
         );
  NAND2X0_RVT U3213 ( .A1(n2926), .A2(n2925), .Y(N382) );
  AO22X1_RVT U3214 ( .A1(\inq_ary[14][121] ), .A2(n3325), .A3(
        \inq_ary[7][121] ), .A4(n3322), .Y(n2930) );
  AO22X1_RVT U3215 ( .A1(\inq_ary[3][121] ), .A2(n3310), .A3(
        \inq_ary[11][121] ), .A4(n3316), .Y(n2929) );
  AO22X1_RVT U3216 ( .A1(\inq_ary[12][121] ), .A2(n3303), .A3(
        \inq_ary[0][121] ), .A4(n3315), .Y(n2928) );
  AO22X1_RVT U3217 ( .A1(\inq_ary[8][121] ), .A2(n3313), .A3(
        \inq_ary[10][121] ), .A4(n3326), .Y(n2927) );
  NOR4X1_RVT U3218 ( .A1(n2930), .A2(n2929), .A3(n2928), .A4(n2927), .Y(n2936)
         );
  AO22X1_RVT U3219 ( .A1(\inq_ary[5][121] ), .A2(n3298), .A3(\inq_ary[4][121] ), .A4(n3321), .Y(n2934) );
  AO22X1_RVT U3220 ( .A1(\inq_ary[6][121] ), .A2(n3311), .A3(
        \inq_ary[13][121] ), .A4(n3323), .Y(n2933) );
  AO22X1_RVT U3221 ( .A1(\inq_ary[1][121] ), .A2(n3324), .A3(\inq_ary[9][121] ), .A4(n3314), .Y(n2932) );
  AO22X1_RVT U3222 ( .A1(\inq_ary[15][121] ), .A2(n3312), .A3(
        \inq_ary[2][121] ), .A4(n3271), .Y(n2931) );
  NOR4X1_RVT U3223 ( .A1(n2934), .A2(n2933), .A3(n2932), .A4(n2931), .Y(n2935)
         );
  NAND2X0_RVT U3224 ( .A1(n2936), .A2(n2935), .Y(N383) );
  AO22X1_RVT U3225 ( .A1(\inq_ary[10][122] ), .A2(n3326), .A3(
        \inq_ary[5][122] ), .A4(n3298), .Y(n2940) );
  AO22X1_RVT U3226 ( .A1(\inq_ary[1][122] ), .A2(n3324), .A3(\inq_ary[7][122] ), .A4(n3322), .Y(n2939) );
  AO22X1_RVT U3227 ( .A1(\inq_ary[2][122] ), .A2(n3271), .A3(
        \inq_ary[12][122] ), .A4(n3303), .Y(n2938) );
  AO22X1_RVT U3228 ( .A1(\inq_ary[15][122] ), .A2(n3312), .A3(
        \inq_ary[6][122] ), .A4(n3311), .Y(n2937) );
  NOR4X1_RVT U3229 ( .A1(n2940), .A2(n2939), .A3(n2938), .A4(n2937), .Y(n2946)
         );
  AO22X1_RVT U3230 ( .A1(\inq_ary[13][122] ), .A2(n3323), .A3(
        \inq_ary[4][122] ), .A4(n3321), .Y(n2944) );
  AO22X1_RVT U3231 ( .A1(\inq_ary[14][122] ), .A2(n3325), .A3(
        \inq_ary[0][122] ), .A4(n3315), .Y(n2943) );
  AO22X1_RVT U3232 ( .A1(\inq_ary[11][122] ), .A2(n3316), .A3(
        \inq_ary[9][122] ), .A4(n3314), .Y(n2942) );
  AO22X1_RVT U3233 ( .A1(\inq_ary[8][122] ), .A2(n3313), .A3(\inq_ary[3][122] ), .A4(n3310), .Y(n2941) );
  NOR4X1_RVT U3234 ( .A1(n2944), .A2(n2943), .A3(n2942), .A4(n2941), .Y(n2945)
         );
  NAND2X0_RVT U3235 ( .A1(n2946), .A2(n2945), .Y(N384) );
  AO22X1_RVT U3236 ( .A1(\inq_ary[8][123] ), .A2(n3313), .A3(
        \inq_ary[13][123] ), .A4(n3323), .Y(n2950) );
  AO22X1_RVT U3237 ( .A1(\inq_ary[14][123] ), .A2(n3325), .A3(
        \inq_ary[7][123] ), .A4(n3322), .Y(n2949) );
  AO22X1_RVT U3238 ( .A1(\inq_ary[15][123] ), .A2(n3312), .A3(
        \inq_ary[3][123] ), .A4(n3310), .Y(n2948) );
  AO22X1_RVT U3239 ( .A1(\inq_ary[2][123] ), .A2(n3271), .A3(
        \inq_ary[12][123] ), .A4(n3303), .Y(n2947) );
  NOR4X1_RVT U3240 ( .A1(n2950), .A2(n2949), .A3(n2948), .A4(n2947), .Y(n2956)
         );
  AO22X1_RVT U3241 ( .A1(\inq_ary[5][123] ), .A2(n3298), .A3(\inq_ary[6][123] ), .A4(n3311), .Y(n2954) );
  AO22X1_RVT U3242 ( .A1(\inq_ary[11][123] ), .A2(n3316), .A3(
        \inq_ary[9][123] ), .A4(n3314), .Y(n2953) );
  AO22X1_RVT U3243 ( .A1(\inq_ary[4][123] ), .A2(n3321), .A3(
        \inq_ary[10][123] ), .A4(n3326), .Y(n2952) );
  AO22X1_RVT U3244 ( .A1(\inq_ary[1][123] ), .A2(n3324), .A3(\inq_ary[0][123] ), .A4(n3315), .Y(n2951) );
  NOR4X1_RVT U3245 ( .A1(n2954), .A2(n2953), .A3(n2952), .A4(n2951), .Y(n2955)
         );
  NAND2X0_RVT U3246 ( .A1(n2956), .A2(n2955), .Y(N385) );
  AO22X1_RVT U3247 ( .A1(\inq_ary[6][124] ), .A2(n3311), .A3(
        \inq_ary[11][124] ), .A4(n3316), .Y(n2960) );
  AO22X1_RVT U3248 ( .A1(\inq_ary[10][124] ), .A2(n3326), .A3(
        \inq_ary[14][124] ), .A4(n3325), .Y(n2959) );
  AO22X1_RVT U3249 ( .A1(\inq_ary[4][124] ), .A2(n3321), .A3(
        \inq_ary[13][124] ), .A4(n3323), .Y(n2958) );
  AO22X1_RVT U3250 ( .A1(\inq_ary[9][124] ), .A2(n3314), .A3(\inq_ary[5][124] ), .A4(n3298), .Y(n2957) );
  NOR4X1_RVT U3251 ( .A1(n2960), .A2(n2959), .A3(n2958), .A4(n2957), .Y(n2966)
         );
  AO22X1_RVT U3252 ( .A1(\inq_ary[12][124] ), .A2(n3303), .A3(
        \inq_ary[3][124] ), .A4(n3310), .Y(n2964) );
  AO22X1_RVT U3253 ( .A1(\inq_ary[2][124] ), .A2(n3271), .A3(\inq_ary[8][124] ), .A4(n3313), .Y(n2963) );
  AO22X1_RVT U3254 ( .A1(\inq_ary[7][124] ), .A2(n3322), .A3(\inq_ary[0][124] ), .A4(n3315), .Y(n2962) );
  AO22X1_RVT U3255 ( .A1(\inq_ary[1][124] ), .A2(n3324), .A3(
        \inq_ary[15][124] ), .A4(n3312), .Y(n2961) );
  NOR4X1_RVT U3256 ( .A1(n2964), .A2(n2963), .A3(n2962), .A4(n2961), .Y(n2965)
         );
  NAND2X0_RVT U3257 ( .A1(n2966), .A2(n2965), .Y(N386) );
  AO22X1_RVT U3258 ( .A1(\inq_ary[5][125] ), .A2(n3298), .A3(
        \inq_ary[10][125] ), .A4(n3326), .Y(n2970) );
  AO22X1_RVT U3259 ( .A1(\inq_ary[15][125] ), .A2(n3312), .A3(
        \inq_ary[0][125] ), .A4(n3315), .Y(n2969) );
  AO22X1_RVT U3260 ( .A1(\inq_ary[14][125] ), .A2(n3325), .A3(
        \inq_ary[11][125] ), .A4(n3316), .Y(n2968) );
  AO22X1_RVT U3261 ( .A1(\inq_ary[8][125] ), .A2(n3313), .A3(\inq_ary[4][125] ), .A4(n3321), .Y(n2967) );
  NOR4X1_RVT U3262 ( .A1(n2970), .A2(n2969), .A3(n2968), .A4(n2967), .Y(n2976)
         );
  AO22X1_RVT U3263 ( .A1(\inq_ary[2][125] ), .A2(n3271), .A3(\inq_ary[3][125] ), .A4(n3310), .Y(n2974) );
  AO22X1_RVT U3264 ( .A1(\inq_ary[7][125] ), .A2(n3322), .A3(
        \inq_ary[13][125] ), .A4(n3323), .Y(n2973) );
  AO22X1_RVT U3265 ( .A1(\inq_ary[12][125] ), .A2(n3303), .A3(
        \inq_ary[6][125] ), .A4(n3311), .Y(n2972) );
  AO22X1_RVT U3266 ( .A1(\inq_ary[1][125] ), .A2(n3324), .A3(\inq_ary[9][125] ), .A4(n3314), .Y(n2971) );
  NOR4X1_RVT U3267 ( .A1(n2974), .A2(n2973), .A3(n2972), .A4(n2971), .Y(n2975)
         );
  NAND2X0_RVT U3268 ( .A1(n2976), .A2(n2975), .Y(N387) );
  AO22X1_RVT U3269 ( .A1(\inq_ary[6][126] ), .A2(n3311), .A3(\inq_ary[0][126] ), .A4(n3315), .Y(n2980) );
  AO22X1_RVT U3270 ( .A1(\inq_ary[3][126] ), .A2(n3310), .A3(\inq_ary[7][126] ), .A4(n3322), .Y(n2979) );
  AO22X1_RVT U3271 ( .A1(\inq_ary[9][126] ), .A2(n3314), .A3(
        \inq_ary[12][126] ), .A4(n3303), .Y(n2978) );
  AO22X1_RVT U3272 ( .A1(\inq_ary[15][126] ), .A2(n3312), .A3(
        \inq_ary[8][126] ), .A4(n3313), .Y(n2977) );
  NOR4X1_RVT U3273 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .Y(n2986)
         );
  AO22X1_RVT U3274 ( .A1(\inq_ary[13][126] ), .A2(n3323), .A3(
        \inq_ary[5][126] ), .A4(n3298), .Y(n2984) );
  AO22X1_RVT U3275 ( .A1(\inq_ary[4][126] ), .A2(n3321), .A3(
        \inq_ary[11][126] ), .A4(n3316), .Y(n2983) );
  AO22X1_RVT U3276 ( .A1(\inq_ary[2][126] ), .A2(n3271), .A3(\inq_ary[1][126] ), .A4(n3324), .Y(n2982) );
  AO22X1_RVT U3277 ( .A1(\inq_ary[14][126] ), .A2(n3325), .A3(
        \inq_ary[10][126] ), .A4(n3326), .Y(n2981) );
  NOR4X1_RVT U3278 ( .A1(n2984), .A2(n2983), .A3(n2982), .A4(n2981), .Y(n2985)
         );
  NAND2X0_RVT U3279 ( .A1(n2986), .A2(n2985), .Y(N388) );
  AO22X1_RVT U3280 ( .A1(\inq_ary[7][127] ), .A2(n3322), .A3(\inq_ary[1][127] ), .A4(n3324), .Y(n2990) );
  AO22X1_RVT U3281 ( .A1(\inq_ary[11][127] ), .A2(n3316), .A3(
        \inq_ary[3][127] ), .A4(n3310), .Y(n2989) );
  AO22X1_RVT U3282 ( .A1(\inq_ary[14][127] ), .A2(n3325), .A3(
        \inq_ary[13][127] ), .A4(n3323), .Y(n2988) );
  AO22X1_RVT U3283 ( .A1(\inq_ary[4][127] ), .A2(n3321), .A3(
        \inq_ary[12][127] ), .A4(n3303), .Y(n2987) );
  NOR4X1_RVT U3284 ( .A1(n2990), .A2(n2989), .A3(n2988), .A4(n2987), .Y(n2996)
         );
  AO22X1_RVT U3285 ( .A1(\inq_ary[2][127] ), .A2(n3271), .A3(
        \inq_ary[10][127] ), .A4(n3326), .Y(n2994) );
  AO22X1_RVT U3286 ( .A1(\inq_ary[9][127] ), .A2(n3314), .A3(\inq_ary[8][127] ), .A4(n3313), .Y(n2993) );
  AO22X1_RVT U3287 ( .A1(\inq_ary[5][127] ), .A2(n3298), .A3(\inq_ary[0][127] ), .A4(n3315), .Y(n2992) );
  AO22X1_RVT U3288 ( .A1(\inq_ary[15][127] ), .A2(n3312), .A3(
        \inq_ary[6][127] ), .A4(n3311), .Y(n2991) );
  NOR4X1_RVT U3289 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .Y(n2995)
         );
  NAND2X0_RVT U3290 ( .A1(n2996), .A2(n2995), .Y(N389) );
  AO22X1_RVT U3291 ( .A1(\inq_ary[10][128] ), .A2(n3326), .A3(
        \inq_ary[15][128] ), .A4(n3312), .Y(n3000) );
  AO22X1_RVT U3292 ( .A1(\inq_ary[5][128] ), .A2(n3298), .A3(
        \inq_ary[13][128] ), .A4(n3323), .Y(n2999) );
  AO22X1_RVT U3293 ( .A1(\inq_ary[0][128] ), .A2(n3315), .A3(\inq_ary[9][128] ), .A4(n3314), .Y(n2998) );
  AO22X1_RVT U3294 ( .A1(\inq_ary[11][128] ), .A2(n3316), .A3(
        \inq_ary[4][128] ), .A4(n3321), .Y(n2997) );
  NOR4X1_RVT U3295 ( .A1(n3000), .A2(n2999), .A3(n2998), .A4(n2997), .Y(n3006)
         );
  AO22X1_RVT U3296 ( .A1(\inq_ary[7][128] ), .A2(n3322), .A3(\inq_ary[3][128] ), .A4(n3310), .Y(n3004) );
  AO22X1_RVT U3297 ( .A1(\inq_ary[8][128] ), .A2(n3313), .A3(\inq_ary[2][128] ), .A4(n3271), .Y(n3003) );
  AO22X1_RVT U3298 ( .A1(\inq_ary[12][128] ), .A2(n3303), .A3(
        \inq_ary[14][128] ), .A4(n3325), .Y(n3002) );
  AO22X1_RVT U3299 ( .A1(\inq_ary[6][128] ), .A2(n3311), .A3(\inq_ary[1][128] ), .A4(n3324), .Y(n3001) );
  NOR4X1_RVT U3300 ( .A1(n3004), .A2(n3003), .A3(n3002), .A4(n3001), .Y(n3005)
         );
  NAND2X0_RVT U3301 ( .A1(n3006), .A2(n3005), .Y(N390) );
  AO22X1_RVT U3302 ( .A1(\inq_ary[7][129] ), .A2(n3322), .A3(
        \inq_ary[12][129] ), .A4(n3303), .Y(n3010) );
  AO22X1_RVT U3303 ( .A1(\inq_ary[15][129] ), .A2(n3312), .A3(
        \inq_ary[2][129] ), .A4(n3271), .Y(n3009) );
  AO22X1_RVT U3304 ( .A1(\inq_ary[1][129] ), .A2(n3324), .A3(
        \inq_ary[14][129] ), .A4(n3325), .Y(n3008) );
  AO22X1_RVT U3305 ( .A1(\inq_ary[3][129] ), .A2(n3310), .A3(
        \inq_ary[11][129] ), .A4(n3316), .Y(n3007) );
  NOR4X1_RVT U3306 ( .A1(n3010), .A2(n3009), .A3(n3008), .A4(n3007), .Y(n3016)
         );
  AO22X1_RVT U3307 ( .A1(\inq_ary[9][129] ), .A2(n3314), .A3(
        \inq_ary[10][129] ), .A4(n3326), .Y(n3014) );
  AO22X1_RVT U3308 ( .A1(\inq_ary[8][129] ), .A2(n3313), .A3(\inq_ary[5][129] ), .A4(n3298), .Y(n3013) );
  AO22X1_RVT U3309 ( .A1(\inq_ary[13][129] ), .A2(n3323), .A3(
        \inq_ary[0][129] ), .A4(n3315), .Y(n3012) );
  AO22X1_RVT U3310 ( .A1(\inq_ary[4][129] ), .A2(n3321), .A3(\inq_ary[6][129] ), .A4(n3311), .Y(n3011) );
  NOR4X1_RVT U3311 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .Y(n3015)
         );
  NAND2X0_RVT U3312 ( .A1(n3016), .A2(n3015), .Y(N391) );
  AO22X1_RVT U3313 ( .A1(\inq_ary[10][130] ), .A2(n3326), .A3(
        \inq_ary[6][130] ), .A4(n3311), .Y(n3020) );
  AO22X1_RVT U3314 ( .A1(\inq_ary[0][130] ), .A2(n3315), .A3(
        \inq_ary[12][130] ), .A4(n3303), .Y(n3019) );
  AO22X1_RVT U3315 ( .A1(\inq_ary[2][130] ), .A2(n3271), .A3(
        \inq_ary[11][130] ), .A4(n3316), .Y(n3018) );
  AO22X1_RVT U3316 ( .A1(\inq_ary[9][130] ), .A2(n3314), .A3(\inq_ary[5][130] ), .A4(n3298), .Y(n3017) );
  NOR4X1_RVT U3317 ( .A1(n3020), .A2(n3019), .A3(n3018), .A4(n3017), .Y(n3026)
         );
  AO22X1_RVT U3318 ( .A1(\inq_ary[4][130] ), .A2(n3321), .A3(\inq_ary[7][130] ), .A4(n3322), .Y(n3024) );
  AO22X1_RVT U3319 ( .A1(\inq_ary[15][130] ), .A2(n3312), .A3(
        \inq_ary[1][130] ), .A4(n3324), .Y(n3023) );
  AO22X1_RVT U3320 ( .A1(\inq_ary[3][130] ), .A2(n3310), .A3(\inq_ary[8][130] ), .A4(n3313), .Y(n3022) );
  AO22X1_RVT U3321 ( .A1(\inq_ary[13][130] ), .A2(n3323), .A3(
        \inq_ary[14][130] ), .A4(n3325), .Y(n3021) );
  NOR4X1_RVT U3322 ( .A1(n3024), .A2(n3023), .A3(n3022), .A4(n3021), .Y(n3025)
         );
  NAND2X0_RVT U3323 ( .A1(n3026), .A2(n3025), .Y(N392) );
  AO22X1_RVT U3324 ( .A1(\inq_ary[9][131] ), .A2(n3314), .A3(
        \inq_ary[10][131] ), .A4(n3326), .Y(n3030) );
  AO22X1_RVT U3325 ( .A1(\inq_ary[2][131] ), .A2(n3271), .A3(\inq_ary[8][131] ), .A4(n3313), .Y(n3029) );
  AO22X1_RVT U3326 ( .A1(\inq_ary[7][131] ), .A2(n3322), .A3(\inq_ary[4][131] ), .A4(n3321), .Y(n3028) );
  AO22X1_RVT U3327 ( .A1(\inq_ary[6][131] ), .A2(n3311), .A3(
        \inq_ary[11][131] ), .A4(n3316), .Y(n3027) );
  NOR4X1_RVT U3328 ( .A1(n3030), .A2(n3029), .A3(n3028), .A4(n3027), .Y(n3036)
         );
  AO22X1_RVT U3329 ( .A1(\inq_ary[1][131] ), .A2(n3324), .A3(\inq_ary[3][131] ), .A4(n3310), .Y(n3034) );
  AO22X1_RVT U3330 ( .A1(\inq_ary[13][131] ), .A2(n3323), .A3(
        \inq_ary[15][131] ), .A4(n3312), .Y(n3033) );
  AO22X1_RVT U3331 ( .A1(\inq_ary[14][131] ), .A2(n3325), .A3(
        \inq_ary[12][131] ), .A4(n3303), .Y(n3032) );
  AO22X1_RVT U3332 ( .A1(\inq_ary[0][131] ), .A2(n3315), .A3(\inq_ary[5][131] ), .A4(n3298), .Y(n3031) );
  NOR4X1_RVT U3333 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n3031), .Y(n3035)
         );
  NAND2X0_RVT U3334 ( .A1(n3036), .A2(n3035), .Y(N393) );
  AO22X1_RVT U3335 ( .A1(\inq_ary[5][132] ), .A2(n3298), .A3(
        \inq_ary[13][132] ), .A4(n3323), .Y(n3040) );
  AO22X1_RVT U3336 ( .A1(\inq_ary[2][132] ), .A2(n3271), .A3(
        \inq_ary[11][132] ), .A4(n3316), .Y(n3039) );
  AO22X1_RVT U3337 ( .A1(\inq_ary[12][132] ), .A2(n3303), .A3(
        \inq_ary[3][132] ), .A4(n3310), .Y(n3038) );
  AO22X1_RVT U3338 ( .A1(\inq_ary[0][132] ), .A2(n3315), .A3(
        \inq_ary[15][132] ), .A4(n3312), .Y(n3037) );
  NOR4X1_RVT U3339 ( .A1(n3040), .A2(n3039), .A3(n3038), .A4(n3037), .Y(n3046)
         );
  AO22X1_RVT U3340 ( .A1(\inq_ary[4][132] ), .A2(n3321), .A3(\inq_ary[8][132] ), .A4(n3313), .Y(n3044) );
  AO22X1_RVT U3341 ( .A1(\inq_ary[1][132] ), .A2(n3324), .A3(\inq_ary[6][132] ), .A4(n3311), .Y(n3043) );
  AO22X1_RVT U3342 ( .A1(\inq_ary[10][132] ), .A2(n3326), .A3(
        \inq_ary[14][132] ), .A4(n3325), .Y(n3042) );
  AO22X1_RVT U3343 ( .A1(\inq_ary[9][132] ), .A2(n3314), .A3(\inq_ary[7][132] ), .A4(n3322), .Y(n3041) );
  NOR4X1_RVT U3344 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .Y(n3045)
         );
  NAND2X0_RVT U3345 ( .A1(n3046), .A2(n3045), .Y(N394) );
  AO22X1_RVT U3346 ( .A1(\inq_ary[6][133] ), .A2(n3311), .A3(\inq_ary[1][133] ), .A4(n3324), .Y(n3050) );
  AO22X1_RVT U3347 ( .A1(\inq_ary[14][133] ), .A2(n3325), .A3(
        \inq_ary[13][133] ), .A4(n3323), .Y(n3049) );
  AO22X1_RVT U3348 ( .A1(\inq_ary[5][133] ), .A2(n3298), .A3(\inq_ary[2][133] ), .A4(n3271), .Y(n3048) );
  AO22X1_RVT U3349 ( .A1(\inq_ary[15][133] ), .A2(n3312), .A3(
        \inq_ary[3][133] ), .A4(n3310), .Y(n3047) );
  NOR4X1_RVT U3350 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .Y(n3056)
         );
  AO22X1_RVT U3351 ( .A1(\inq_ary[0][133] ), .A2(n3315), .A3(\inq_ary[8][133] ), .A4(n3313), .Y(n3054) );
  AO22X1_RVT U3352 ( .A1(\inq_ary[10][133] ), .A2(n3326), .A3(
        \inq_ary[4][133] ), .A4(n3321), .Y(n3053) );
  AO22X1_RVT U3353 ( .A1(\inq_ary[11][133] ), .A2(n3316), .A3(
        \inq_ary[7][133] ), .A4(n3322), .Y(n3052) );
  AO22X1_RVT U3354 ( .A1(\inq_ary[12][133] ), .A2(n3303), .A3(
        \inq_ary[9][133] ), .A4(n3314), .Y(n3051) );
  NOR4X1_RVT U3355 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .Y(n3055)
         );
  NAND2X0_RVT U3356 ( .A1(n3056), .A2(n3055), .Y(N395) );
  AO22X1_RVT U3357 ( .A1(\inq_ary[6][134] ), .A2(n3311), .A3(\inq_ary[3][134] ), .A4(n3310), .Y(n3060) );
  AO22X1_RVT U3358 ( .A1(\inq_ary[4][134] ), .A2(n3321), .A3(\inq_ary[5][134] ), .A4(n3298), .Y(n3059) );
  AO22X1_RVT U3359 ( .A1(\inq_ary[1][134] ), .A2(n3324), .A3(
        \inq_ary[12][134] ), .A4(n3303), .Y(n3058) );
  AO22X1_RVT U3360 ( .A1(\inq_ary[2][134] ), .A2(n3271), .A3(
        \inq_ary[10][134] ), .A4(n3326), .Y(n3057) );
  NOR4X1_RVT U3361 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), .Y(n3066)
         );
  AO22X1_RVT U3362 ( .A1(\inq_ary[14][134] ), .A2(n3325), .A3(
        \inq_ary[13][134] ), .A4(n3323), .Y(n3064) );
  AO22X1_RVT U3363 ( .A1(\inq_ary[15][134] ), .A2(n3312), .A3(
        \inq_ary[7][134] ), .A4(n3322), .Y(n3063) );
  AO22X1_RVT U3364 ( .A1(\inq_ary[0][134] ), .A2(n3315), .A3(\inq_ary[8][134] ), .A4(n3313), .Y(n3062) );
  AO22X1_RVT U3365 ( .A1(\inq_ary[9][134] ), .A2(n3314), .A3(
        \inq_ary[11][134] ), .A4(n3316), .Y(n3061) );
  NOR4X1_RVT U3366 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), .Y(n3065)
         );
  NAND2X0_RVT U3367 ( .A1(n3066), .A2(n3065), .Y(N396) );
  AO22X1_RVT U3368 ( .A1(\inq_ary[14][135] ), .A2(n3325), .A3(
        \inq_ary[11][135] ), .A4(n3316), .Y(n3070) );
  AO22X1_RVT U3369 ( .A1(\inq_ary[4][135] ), .A2(n3321), .A3(\inq_ary[9][135] ), .A4(n3314), .Y(n3069) );
  AO22X1_RVT U3370 ( .A1(\inq_ary[0][135] ), .A2(n3315), .A3(\inq_ary[7][135] ), .A4(n3322), .Y(n3068) );
  AO22X1_RVT U3371 ( .A1(\inq_ary[12][135] ), .A2(n3303), .A3(
        \inq_ary[5][135] ), .A4(n3298), .Y(n3067) );
  NOR4X1_RVT U3372 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .Y(n3076)
         );
  AO22X1_RVT U3373 ( .A1(\inq_ary[1][135] ), .A2(n3324), .A3(\inq_ary[8][135] ), .A4(n3313), .Y(n3074) );
  AO22X1_RVT U3374 ( .A1(\inq_ary[2][135] ), .A2(n3271), .A3(\inq_ary[6][135] ), .A4(n3311), .Y(n3073) );
  AO22X1_RVT U3375 ( .A1(\inq_ary[3][135] ), .A2(n3310), .A3(
        \inq_ary[15][135] ), .A4(n3312), .Y(n3072) );
  AO22X1_RVT U3376 ( .A1(\inq_ary[13][135] ), .A2(n3323), .A3(
        \inq_ary[10][135] ), .A4(n3326), .Y(n3071) );
  NOR4X1_RVT U3377 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .Y(n3075)
         );
  NAND2X0_RVT U3378 ( .A1(n3076), .A2(n3075), .Y(N397) );
  AO22X1_RVT U3379 ( .A1(\inq_ary[11][136] ), .A2(n3316), .A3(
        \inq_ary[15][136] ), .A4(n3312), .Y(n3080) );
  AO22X1_RVT U3380 ( .A1(\inq_ary[13][136] ), .A2(n3323), .A3(
        \inq_ary[12][136] ), .A4(n3303), .Y(n3079) );
  AO22X1_RVT U3381 ( .A1(\inq_ary[10][136] ), .A2(n3326), .A3(
        \inq_ary[4][136] ), .A4(n3321), .Y(n3078) );
  AO22X1_RVT U3382 ( .A1(\inq_ary[7][136] ), .A2(n3322), .A3(
        \inq_ary[14][136] ), .A4(n3325), .Y(n3077) );
  NOR4X1_RVT U3383 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), .Y(n3086)
         );
  AO22X1_RVT U3384 ( .A1(\inq_ary[0][136] ), .A2(n3315), .A3(\inq_ary[3][136] ), .A4(n3310), .Y(n3084) );
  AO22X1_RVT U3385 ( .A1(\inq_ary[2][136] ), .A2(n3271), .A3(\inq_ary[5][136] ), .A4(n3298), .Y(n3083) );
  AO22X1_RVT U3386 ( .A1(\inq_ary[6][136] ), .A2(n3311), .A3(\inq_ary[8][136] ), .A4(n3313), .Y(n3082) );
  AO22X1_RVT U3387 ( .A1(\inq_ary[9][136] ), .A2(n3314), .A3(\inq_ary[1][136] ), .A4(n3324), .Y(n3081) );
  NOR4X1_RVT U3388 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .Y(n3085)
         );
  NAND2X0_RVT U3389 ( .A1(n3086), .A2(n3085), .Y(N398) );
  AO22X1_RVT U3390 ( .A1(\inq_ary[0][137] ), .A2(n3315), .A3(
        \inq_ary[15][137] ), .A4(n3312), .Y(n3090) );
  AO22X1_RVT U3391 ( .A1(\inq_ary[14][137] ), .A2(n3325), .A3(
        \inq_ary[10][137] ), .A4(n3326), .Y(n3089) );
  AO22X1_RVT U3392 ( .A1(\inq_ary[6][137] ), .A2(n3311), .A3(\inq_ary[5][137] ), .A4(n3298), .Y(n3088) );
  AO22X1_RVT U3393 ( .A1(\inq_ary[2][137] ), .A2(n3271), .A3(
        \inq_ary[12][137] ), .A4(n3303), .Y(n3087) );
  NOR4X1_RVT U3394 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .Y(n3096)
         );
  AO22X1_RVT U3395 ( .A1(\inq_ary[1][137] ), .A2(n3324), .A3(\inq_ary[3][137] ), .A4(n3310), .Y(n3094) );
  AO22X1_RVT U3396 ( .A1(\inq_ary[8][137] ), .A2(n3313), .A3(\inq_ary[4][137] ), .A4(n3321), .Y(n3093) );
  AO22X1_RVT U3397 ( .A1(\inq_ary[9][137] ), .A2(n3314), .A3(
        \inq_ary[11][137] ), .A4(n3316), .Y(n3092) );
  AO22X1_RVT U3398 ( .A1(\inq_ary[13][137] ), .A2(n3323), .A3(
        \inq_ary[7][137] ), .A4(n3322), .Y(n3091) );
  NOR4X1_RVT U3399 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .Y(n3095)
         );
  NAND2X0_RVT U3400 ( .A1(n3096), .A2(n3095), .Y(N399) );
  AO22X1_RVT U3401 ( .A1(\inq_ary[10][138] ), .A2(n3326), .A3(
        \inq_ary[12][138] ), .A4(n3303), .Y(n3100) );
  AO22X1_RVT U3402 ( .A1(\inq_ary[9][138] ), .A2(n3314), .A3(\inq_ary[1][138] ), .A4(n3324), .Y(n3099) );
  AO22X1_RVT U3403 ( .A1(\inq_ary[2][138] ), .A2(n3271), .A3(
        \inq_ary[13][138] ), .A4(n3323), .Y(n3098) );
  AO22X1_RVT U3404 ( .A1(\inq_ary[5][138] ), .A2(n3298), .A3(\inq_ary[4][138] ), .A4(n3321), .Y(n3097) );
  NOR4X1_RVT U3405 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .Y(n3106)
         );
  AO22X1_RVT U3406 ( .A1(\inq_ary[3][138] ), .A2(n3310), .A3(\inq_ary[7][138] ), .A4(n3322), .Y(n3104) );
  AO22X1_RVT U3407 ( .A1(\inq_ary[6][138] ), .A2(n3311), .A3(
        \inq_ary[14][138] ), .A4(n3325), .Y(n3103) );
  AO22X1_RVT U3408 ( .A1(\inq_ary[0][138] ), .A2(n3315), .A3(
        \inq_ary[15][138] ), .A4(n3312), .Y(n3102) );
  AO22X1_RVT U3409 ( .A1(\inq_ary[11][138] ), .A2(n3316), .A3(
        \inq_ary[8][138] ), .A4(n3313), .Y(n3101) );
  NOR4X1_RVT U3410 ( .A1(n3104), .A2(n3103), .A3(n3102), .A4(n3101), .Y(n3105)
         );
  NAND2X0_RVT U3411 ( .A1(n3106), .A2(n3105), .Y(N400) );
  AO22X1_RVT U3412 ( .A1(\inq_ary[11][139] ), .A2(n3316), .A3(
        \inq_ary[13][139] ), .A4(n3323), .Y(n3110) );
  AO22X1_RVT U3413 ( .A1(\inq_ary[5][139] ), .A2(n3298), .A3(\inq_ary[7][139] ), .A4(n3322), .Y(n3109) );
  AO22X1_RVT U3414 ( .A1(\inq_ary[4][139] ), .A2(n3321), .A3(
        \inq_ary[10][139] ), .A4(n3326), .Y(n3108) );
  AO22X1_RVT U3415 ( .A1(\inq_ary[14][139] ), .A2(n3325), .A3(
        \inq_ary[8][139] ), .A4(n3313), .Y(n3107) );
  NOR4X1_RVT U3416 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .Y(n3116)
         );
  AO22X1_RVT U3417 ( .A1(\inq_ary[9][139] ), .A2(n3314), .A3(\inq_ary[1][139] ), .A4(n3324), .Y(n3114) );
  AO22X1_RVT U3418 ( .A1(\inq_ary[15][139] ), .A2(n3312), .A3(
        \inq_ary[2][139] ), .A4(n3271), .Y(n3113) );
  AO22X1_RVT U3419 ( .A1(\inq_ary[0][139] ), .A2(n3315), .A3(
        \inq_ary[12][139] ), .A4(n3303), .Y(n3112) );
  AO22X1_RVT U3420 ( .A1(\inq_ary[3][139] ), .A2(n3310), .A3(\inq_ary[6][139] ), .A4(n3311), .Y(n3111) );
  NOR4X1_RVT U3421 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .Y(n3115)
         );
  NAND2X0_RVT U3422 ( .A1(n3116), .A2(n3115), .Y(N401) );
  AO22X1_RVT U3423 ( .A1(\inq_ary[15][140] ), .A2(n3312), .A3(
        \inq_ary[6][140] ), .A4(n3311), .Y(n3120) );
  AO22X1_RVT U3424 ( .A1(\inq_ary[8][140] ), .A2(n3313), .A3(
        \inq_ary[13][140] ), .A4(n3323), .Y(n3119) );
  AO22X1_RVT U3425 ( .A1(\inq_ary[4][140] ), .A2(n3321), .A3(\inq_ary[1][140] ), .A4(n3324), .Y(n3118) );
  AO22X1_RVT U3426 ( .A1(\inq_ary[2][140] ), .A2(n3271), .A3(\inq_ary[5][140] ), .A4(n3298), .Y(n3117) );
  NOR4X1_RVT U3427 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .Y(n3126)
         );
  AO22X1_RVT U3428 ( .A1(\inq_ary[10][140] ), .A2(n3326), .A3(
        \inq_ary[3][140] ), .A4(n3310), .Y(n3124) );
  AO22X1_RVT U3429 ( .A1(\inq_ary[0][140] ), .A2(n3315), .A3(\inq_ary[9][140] ), .A4(n3314), .Y(n3123) );
  AO22X1_RVT U3430 ( .A1(\inq_ary[12][140] ), .A2(n3303), .A3(
        \inq_ary[11][140] ), .A4(n3316), .Y(n3122) );
  AO22X1_RVT U3431 ( .A1(\inq_ary[7][140] ), .A2(n3322), .A3(
        \inq_ary[14][140] ), .A4(n3325), .Y(n3121) );
  NOR4X1_RVT U3432 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .Y(n3125)
         );
  NAND2X0_RVT U3433 ( .A1(n3126), .A2(n3125), .Y(N402) );
  AO22X1_RVT U3434 ( .A1(\inq_ary[10][141] ), .A2(n3326), .A3(
        \inq_ary[11][141] ), .A4(n3316), .Y(n3130) );
  AO22X1_RVT U3435 ( .A1(\inq_ary[14][141] ), .A2(n3325), .A3(
        \inq_ary[12][141] ), .A4(n3303), .Y(n3129) );
  AO22X1_RVT U3436 ( .A1(\inq_ary[0][141] ), .A2(n3315), .A3(\inq_ary[7][141] ), .A4(n3322), .Y(n3128) );
  AO22X1_RVT U3437 ( .A1(\inq_ary[2][141] ), .A2(n3271), .A3(\inq_ary[9][141] ), .A4(n3314), .Y(n3127) );
  NOR4X1_RVT U3438 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .Y(n3136)
         );
  AO22X1_RVT U3439 ( .A1(\inq_ary[15][141] ), .A2(n3312), .A3(
        \inq_ary[13][141] ), .A4(n3323), .Y(n3134) );
  AO22X1_RVT U3440 ( .A1(\inq_ary[8][141] ), .A2(n3313), .A3(\inq_ary[6][141] ), .A4(n3311), .Y(n3133) );
  AO22X1_RVT U3441 ( .A1(\inq_ary[1][141] ), .A2(n3324), .A3(\inq_ary[5][141] ), .A4(n3298), .Y(n3132) );
  AO22X1_RVT U3442 ( .A1(\inq_ary[4][141] ), .A2(n3321), .A3(\inq_ary[3][141] ), .A4(n3310), .Y(n3131) );
  NOR4X1_RVT U3443 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .Y(n3135)
         );
  NAND2X0_RVT U3444 ( .A1(n3136), .A2(n3135), .Y(N403) );
  AO22X1_RVT U3445 ( .A1(\inq_ary[4][142] ), .A2(n3321), .A3(\inq_ary[0][142] ), .A4(n3315), .Y(n3140) );
  AO22X1_RVT U3446 ( .A1(\inq_ary[5][142] ), .A2(n3298), .A3(\inq_ary[7][142] ), .A4(n3322), .Y(n3139) );
  AO22X1_RVT U3447 ( .A1(\inq_ary[1][142] ), .A2(n3324), .A3(\inq_ary[6][142] ), .A4(n3311), .Y(n3138) );
  AO22X1_RVT U3448 ( .A1(\inq_ary[14][142] ), .A2(n3325), .A3(
        \inq_ary[11][142] ), .A4(n3316), .Y(n3137) );
  NOR4X1_RVT U3449 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .Y(n3146)
         );
  AO22X1_RVT U3450 ( .A1(\inq_ary[12][142] ), .A2(n3303), .A3(
        \inq_ary[3][142] ), .A4(n3310), .Y(n3144) );
  AO22X1_RVT U3451 ( .A1(\inq_ary[15][142] ), .A2(n3312), .A3(
        \inq_ary[13][142] ), .A4(n3323), .Y(n3143) );
  AO22X1_RVT U3452 ( .A1(\inq_ary[2][142] ), .A2(n3271), .A3(
        \inq_ary[10][142] ), .A4(n3326), .Y(n3142) );
  AO22X1_RVT U3453 ( .A1(\inq_ary[8][142] ), .A2(n3313), .A3(\inq_ary[9][142] ), .A4(n3314), .Y(n3141) );
  NOR4X1_RVT U3454 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .Y(n3145)
         );
  NAND2X0_RVT U3455 ( .A1(n3146), .A2(n3145), .Y(N404) );
  AO22X1_RVT U3456 ( .A1(\inq_ary[3][143] ), .A2(n3310), .A3(
        \inq_ary[10][143] ), .A4(n3326), .Y(n3150) );
  AO22X1_RVT U3457 ( .A1(\inq_ary[14][143] ), .A2(n3325), .A3(
        \inq_ary[5][143] ), .A4(n3298), .Y(n3149) );
  AO22X1_RVT U3458 ( .A1(\inq_ary[9][143] ), .A2(n3314), .A3(\inq_ary[1][143] ), .A4(n3324), .Y(n3148) );
  AO22X1_RVT U3459 ( .A1(\inq_ary[13][143] ), .A2(n3323), .A3(
        \inq_ary[8][143] ), .A4(n3313), .Y(n3147) );
  NOR4X1_RVT U3460 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .Y(n3156)
         );
  AO22X1_RVT U3461 ( .A1(\inq_ary[2][143] ), .A2(n3271), .A3(
        \inq_ary[12][143] ), .A4(n3303), .Y(n3154) );
  AO22X1_RVT U3462 ( .A1(\inq_ary[15][143] ), .A2(n3312), .A3(
        \inq_ary[7][143] ), .A4(n3322), .Y(n3153) );
  AO22X1_RVT U3463 ( .A1(\inq_ary[11][143] ), .A2(n3316), .A3(
        \inq_ary[0][143] ), .A4(n3315), .Y(n3152) );
  AO22X1_RVT U3464 ( .A1(\inq_ary[4][143] ), .A2(n3321), .A3(\inq_ary[6][143] ), .A4(n3311), .Y(n3151) );
  NOR4X1_RVT U3465 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .Y(n3155)
         );
  NAND2X0_RVT U3466 ( .A1(n3156), .A2(n3155), .Y(N405) );
  AO22X1_RVT U3467 ( .A1(\inq_ary[12][144] ), .A2(n3303), .A3(
        \inq_ary[8][144] ), .A4(n3313), .Y(n3160) );
  AO22X1_RVT U3468 ( .A1(\inq_ary[10][144] ), .A2(n3326), .A3(
        \inq_ary[9][144] ), .A4(n3314), .Y(n3159) );
  AO22X1_RVT U3469 ( .A1(\inq_ary[7][144] ), .A2(n3322), .A3(
        \inq_ary[15][144] ), .A4(n3312), .Y(n3158) );
  AO22X1_RVT U3470 ( .A1(\inq_ary[11][144] ), .A2(n3316), .A3(
        \inq_ary[13][144] ), .A4(n3323), .Y(n3157) );
  NOR4X1_RVT U3471 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .Y(n3166)
         );
  AO22X1_RVT U3472 ( .A1(\inq_ary[5][144] ), .A2(n3298), .A3(\inq_ary[6][144] ), .A4(n3311), .Y(n3164) );
  AO22X1_RVT U3473 ( .A1(\inq_ary[4][144] ), .A2(n3321), .A3(\inq_ary[2][144] ), .A4(n3271), .Y(n3163) );
  AO22X1_RVT U3474 ( .A1(\inq_ary[14][144] ), .A2(n3325), .A3(
        \inq_ary[3][144] ), .A4(n3310), .Y(n3162) );
  AO22X1_RVT U3475 ( .A1(\inq_ary[0][144] ), .A2(n3315), .A3(\inq_ary[1][144] ), .A4(n3324), .Y(n3161) );
  NOR4X1_RVT U3476 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .Y(n3165)
         );
  NAND2X0_RVT U3477 ( .A1(n3166), .A2(n3165), .Y(N406) );
  AO22X1_RVT U3478 ( .A1(\inq_ary[5][145] ), .A2(n3298), .A3(
        \inq_ary[13][145] ), .A4(n3323), .Y(n3170) );
  AO22X1_RVT U3479 ( .A1(\inq_ary[2][145] ), .A2(n3271), .A3(\inq_ary[6][145] ), .A4(n3311), .Y(n3169) );
  AO22X1_RVT U3480 ( .A1(\inq_ary[14][145] ), .A2(n3325), .A3(
        \inq_ary[15][145] ), .A4(n3312), .Y(n3168) );
  AO22X1_RVT U3481 ( .A1(\inq_ary[7][145] ), .A2(n3322), .A3(\inq_ary[3][145] ), .A4(n3310), .Y(n3167) );
  NOR4X1_RVT U3482 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .Y(n3176)
         );
  AO22X1_RVT U3483 ( .A1(\inq_ary[12][145] ), .A2(n3303), .A3(
        \inq_ary[10][145] ), .A4(n3326), .Y(n3174) );
  AO22X1_RVT U3484 ( .A1(\inq_ary[9][145] ), .A2(n3314), .A3(\inq_ary[8][145] ), .A4(n3313), .Y(n3173) );
  AO22X1_RVT U3485 ( .A1(\inq_ary[1][145] ), .A2(n3324), .A3(\inq_ary[4][145] ), .A4(n3321), .Y(n3172) );
  AO22X1_RVT U3486 ( .A1(\inq_ary[0][145] ), .A2(n3315), .A3(
        \inq_ary[11][145] ), .A4(n3316), .Y(n3171) );
  NOR4X1_RVT U3487 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .Y(n3175)
         );
  NAND2X0_RVT U3488 ( .A1(n3176), .A2(n3175), .Y(N407) );
  AO22X1_RVT U3489 ( .A1(\inq_ary[0][146] ), .A2(n3315), .A3(\inq_ary[2][146] ), .A4(n3271), .Y(n3180) );
  AO22X1_RVT U3490 ( .A1(\inq_ary[8][146] ), .A2(n3313), .A3(\inq_ary[3][146] ), .A4(n3310), .Y(n3179) );
  AO22X1_RVT U3491 ( .A1(\inq_ary[9][146] ), .A2(n3314), .A3(\inq_ary[1][146] ), .A4(n3324), .Y(n3178) );
  AO22X1_RVT U3492 ( .A1(\inq_ary[6][146] ), .A2(n3311), .A3(
        \inq_ary[10][146] ), .A4(n3326), .Y(n3177) );
  NOR4X1_RVT U3493 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .Y(n3186)
         );
  AO22X1_RVT U3494 ( .A1(\inq_ary[14][146] ), .A2(n3325), .A3(
        \inq_ary[15][146] ), .A4(n3312), .Y(n3184) );
  AO22X1_RVT U3495 ( .A1(\inq_ary[4][146] ), .A2(n3321), .A3(
        \inq_ary[11][146] ), .A4(n3316), .Y(n3183) );
  AO22X1_RVT U3496 ( .A1(\inq_ary[5][146] ), .A2(n3298), .A3(
        \inq_ary[12][146] ), .A4(n3303), .Y(n3182) );
  AO22X1_RVT U3497 ( .A1(\inq_ary[7][146] ), .A2(n3322), .A3(
        \inq_ary[13][146] ), .A4(n3323), .Y(n3181) );
  NOR4X1_RVT U3498 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .Y(n3185)
         );
  NAND2X0_RVT U3499 ( .A1(n3186), .A2(n3185), .Y(N408) );
  AO22X1_RVT U3500 ( .A1(\inq_ary[14][147] ), .A2(n3325), .A3(
        \inq_ary[13][147] ), .A4(n3323), .Y(n3190) );
  AO22X1_RVT U3501 ( .A1(\inq_ary[10][147] ), .A2(n3326), .A3(
        \inq_ary[2][147] ), .A4(n3271), .Y(n3189) );
  AO22X1_RVT U3502 ( .A1(\inq_ary[11][147] ), .A2(n3316), .A3(
        \inq_ary[0][147] ), .A4(n3315), .Y(n3188) );
  AO22X1_RVT U3503 ( .A1(\inq_ary[12][147] ), .A2(n3303), .A3(
        \inq_ary[8][147] ), .A4(n3313), .Y(n3187) );
  NOR4X1_RVT U3504 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .Y(n3196)
         );
  AO22X1_RVT U3505 ( .A1(\inq_ary[7][147] ), .A2(n3322), .A3(\inq_ary[3][147] ), .A4(n3310), .Y(n3194) );
  AO22X1_RVT U3506 ( .A1(\inq_ary[5][147] ), .A2(n3298), .A3(\inq_ary[4][147] ), .A4(n3321), .Y(n3193) );
  AO22X1_RVT U3507 ( .A1(\inq_ary[6][147] ), .A2(n3311), .A3(
        \inq_ary[15][147] ), .A4(n3312), .Y(n3192) );
  AO22X1_RVT U3508 ( .A1(\inq_ary[9][147] ), .A2(n3314), .A3(\inq_ary[1][147] ), .A4(n3324), .Y(n3191) );
  NOR4X1_RVT U3509 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .Y(n3195)
         );
  NAND2X0_RVT U3510 ( .A1(n3196), .A2(n3195), .Y(N409) );
  AO22X1_RVT U3511 ( .A1(\inq_ary[12][148] ), .A2(n3303), .A3(
        \inq_ary[3][148] ), .A4(n3310), .Y(n3200) );
  AO22X1_RVT U3512 ( .A1(\inq_ary[10][148] ), .A2(n3326), .A3(
        \inq_ary[1][148] ), .A4(n3324), .Y(n3199) );
  AO22X1_RVT U3513 ( .A1(\inq_ary[6][148] ), .A2(n3311), .A3(
        \inq_ary[14][148] ), .A4(n3325), .Y(n3198) );
  AO22X1_RVT U3514 ( .A1(\inq_ary[11][148] ), .A2(n3316), .A3(
        \inq_ary[15][148] ), .A4(n3312), .Y(n3197) );
  NOR4X1_RVT U3515 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .Y(n3206)
         );
  AO22X1_RVT U3516 ( .A1(\inq_ary[4][148] ), .A2(n3321), .A3(\inq_ary[5][148] ), .A4(n3298), .Y(n3204) );
  AO22X1_RVT U3517 ( .A1(\inq_ary[0][148] ), .A2(n3315), .A3(\inq_ary[9][148] ), .A4(n3314), .Y(n3203) );
  AO22X1_RVT U3518 ( .A1(\inq_ary[13][148] ), .A2(n3323), .A3(
        \inq_ary[2][148] ), .A4(n3271), .Y(n3202) );
  AO22X1_RVT U3519 ( .A1(\inq_ary[8][148] ), .A2(n3313), .A3(\inq_ary[7][148] ), .A4(n3322), .Y(n3201) );
  NOR4X1_RVT U3520 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .Y(n3205)
         );
  NAND2X0_RVT U3521 ( .A1(n3206), .A2(n3205), .Y(N410) );
  AO22X1_RVT U3522 ( .A1(\inq_ary[6][149] ), .A2(n3311), .A3(\inq_ary[7][149] ), .A4(n3322), .Y(n3210) );
  AO22X1_RVT U3523 ( .A1(\inq_ary[10][149] ), .A2(n3326), .A3(
        \inq_ary[14][149] ), .A4(n3325), .Y(n3209) );
  AO22X1_RVT U3524 ( .A1(\inq_ary[0][149] ), .A2(n3315), .A3(\inq_ary[5][149] ), .A4(n3298), .Y(n3208) );
  AO22X1_RVT U3525 ( .A1(\inq_ary[9][149] ), .A2(n3314), .A3(\inq_ary[8][149] ), .A4(n3313), .Y(n3207) );
  NOR4X1_RVT U3526 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .Y(n3216)
         );
  AO22X1_RVT U3527 ( .A1(\inq_ary[12][149] ), .A2(n3303), .A3(
        \inq_ary[13][149] ), .A4(n3323), .Y(n3214) );
  AO22X1_RVT U3528 ( .A1(\inq_ary[3][149] ), .A2(n3310), .A3(\inq_ary[4][149] ), .A4(n3321), .Y(n3213) );
  AO22X1_RVT U3529 ( .A1(\inq_ary[15][149] ), .A2(n3312), .A3(
        \inq_ary[2][149] ), .A4(n3271), .Y(n3212) );
  AO22X1_RVT U3530 ( .A1(\inq_ary[11][149] ), .A2(n3316), .A3(
        \inq_ary[1][149] ), .A4(n3324), .Y(n3211) );
  NOR4X1_RVT U3531 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .Y(n3215)
         );
  NAND2X0_RVT U3532 ( .A1(n3216), .A2(n3215), .Y(N411) );
  AO22X1_RVT U3533 ( .A1(\inq_ary[8][150] ), .A2(n3313), .A3(
        \inq_ary[12][150] ), .A4(n3303), .Y(n3220) );
  AO22X1_RVT U3534 ( .A1(\inq_ary[4][150] ), .A2(n3321), .A3(\inq_ary[0][150] ), .A4(n3315), .Y(n3219) );
  AO22X1_RVT U3535 ( .A1(\inq_ary[6][150] ), .A2(n3311), .A3(\inq_ary[3][150] ), .A4(n3310), .Y(n3218) );
  AO22X1_RVT U3536 ( .A1(\inq_ary[11][150] ), .A2(n3316), .A3(
        \inq_ary[5][150] ), .A4(n3298), .Y(n3217) );
  NOR4X1_RVT U3537 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .Y(n3226)
         );
  AO22X1_RVT U3538 ( .A1(\inq_ary[14][150] ), .A2(n3325), .A3(
        \inq_ary[9][150] ), .A4(n3314), .Y(n3224) );
  AO22X1_RVT U3539 ( .A1(\inq_ary[1][150] ), .A2(n3324), .A3(
        \inq_ary[10][150] ), .A4(n3326), .Y(n3223) );
  AO22X1_RVT U3540 ( .A1(\inq_ary[7][150] ), .A2(n3322), .A3(\inq_ary[2][150] ), .A4(n3271), .Y(n3222) );
  AO22X1_RVT U3541 ( .A1(\inq_ary[13][150] ), .A2(n3323), .A3(
        \inq_ary[15][150] ), .A4(n3312), .Y(n3221) );
  NOR4X1_RVT U3542 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .Y(n3225)
         );
  NAND2X0_RVT U3543 ( .A1(n3226), .A2(n3225), .Y(N412) );
  AO22X1_RVT U3544 ( .A1(\inq_ary[4][151] ), .A2(n3321), .A3(\inq_ary[6][151] ), .A4(n3311), .Y(n3230) );
  AO22X1_RVT U3545 ( .A1(\inq_ary[12][151] ), .A2(n3303), .A3(
        \inq_ary[0][151] ), .A4(n3315), .Y(n3229) );
  AO22X1_RVT U3546 ( .A1(\inq_ary[9][151] ), .A2(n3314), .A3(
        \inq_ary[11][151] ), .A4(n3316), .Y(n3228) );
  AO22X1_RVT U3547 ( .A1(\inq_ary[13][151] ), .A2(n3323), .A3(
        \inq_ary[8][151] ), .A4(n3313), .Y(n3227) );
  NOR4X1_RVT U3548 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .Y(n3236)
         );
  AO22X1_RVT U3549 ( .A1(\inq_ary[10][151] ), .A2(n3326), .A3(
        \inq_ary[1][151] ), .A4(n3324), .Y(n3234) );
  AO22X1_RVT U3550 ( .A1(\inq_ary[2][151] ), .A2(n3271), .A3(\inq_ary[3][151] ), .A4(n3310), .Y(n3233) );
  AO22X1_RVT U3551 ( .A1(\inq_ary[14][151] ), .A2(n3325), .A3(
        \inq_ary[7][151] ), .A4(n3322), .Y(n3232) );
  AO22X1_RVT U3552 ( .A1(\inq_ary[15][151] ), .A2(n3312), .A3(
        \inq_ary[5][151] ), .A4(n3298), .Y(n3231) );
  NOR4X1_RVT U3553 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .Y(n3235)
         );
  NAND2X0_RVT U3554 ( .A1(n3236), .A2(n3235), .Y(N413) );
  AO22X1_RVT U3555 ( .A1(\inq_ary[3][152] ), .A2(n3310), .A3(
        \inq_ary[11][152] ), .A4(n3316), .Y(n3240) );
  AO22X1_RVT U3556 ( .A1(\inq_ary[15][152] ), .A2(n3312), .A3(
        \inq_ary[2][152] ), .A4(n3271), .Y(n3239) );
  AO22X1_RVT U3557 ( .A1(\inq_ary[10][152] ), .A2(n3326), .A3(
        \inq_ary[7][152] ), .A4(n3322), .Y(n3238) );
  AO22X1_RVT U3558 ( .A1(\inq_ary[0][152] ), .A2(n3315), .A3(\inq_ary[5][152] ), .A4(n3298), .Y(n3237) );
  NOR4X1_RVT U3559 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .Y(n3246)
         );
  AO22X1_RVT U3560 ( .A1(\inq_ary[9][152] ), .A2(n3314), .A3(\inq_ary[6][152] ), .A4(n3311), .Y(n3244) );
  AO22X1_RVT U3561 ( .A1(\inq_ary[4][152] ), .A2(n3321), .A3(\inq_ary[8][152] ), .A4(n3313), .Y(n3243) );
  AO22X1_RVT U3562 ( .A1(\inq_ary[14][152] ), .A2(n3325), .A3(
        \inq_ary[13][152] ), .A4(n3323), .Y(n3242) );
  AO22X1_RVT U3563 ( .A1(\inq_ary[1][152] ), .A2(n3324), .A3(
        \inq_ary[12][152] ), .A4(n3303), .Y(n3241) );
  NOR4X1_RVT U3564 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .Y(n3245)
         );
  NAND2X0_RVT U3565 ( .A1(n3246), .A2(n3245), .Y(N414) );
  AO22X1_RVT U3566 ( .A1(\inq_ary[4][153] ), .A2(n3321), .A3(\inq_ary[8][153] ), .A4(n3313), .Y(n3250) );
  AO22X1_RVT U3567 ( .A1(\inq_ary[14][153] ), .A2(n3325), .A3(
        \inq_ary[6][153] ), .A4(n3311), .Y(n3249) );
  AO22X1_RVT U3568 ( .A1(\inq_ary[3][153] ), .A2(n3310), .A3(
        \inq_ary[13][153] ), .A4(n3323), .Y(n3248) );
  AO22X1_RVT U3569 ( .A1(\inq_ary[7][153] ), .A2(n3322), .A3(
        \inq_ary[12][153] ), .A4(n3303), .Y(n3247) );
  NOR4X1_RVT U3570 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .Y(n3256)
         );
  AO22X1_RVT U3571 ( .A1(\inq_ary[2][153] ), .A2(n3271), .A3(\inq_ary[1][153] ), .A4(n3324), .Y(n3254) );
  AO22X1_RVT U3572 ( .A1(\inq_ary[15][153] ), .A2(n3312), .A3(
        \inq_ary[0][153] ), .A4(n3315), .Y(n3253) );
  AO22X1_RVT U3573 ( .A1(\inq_ary[5][153] ), .A2(n3298), .A3(\inq_ary[9][153] ), .A4(n3314), .Y(n3252) );
  AO22X1_RVT U3574 ( .A1(\inq_ary[10][153] ), .A2(n3326), .A3(
        \inq_ary[11][153] ), .A4(n3316), .Y(n3251) );
  NOR4X1_RVT U3575 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .Y(n3255)
         );
  NAND2X0_RVT U3576 ( .A1(n3256), .A2(n3255), .Y(N415) );
  AO22X1_RVT U3577 ( .A1(\inq_ary[5][154] ), .A2(n3298), .A3(\inq_ary[4][154] ), .A4(n3321), .Y(n3260) );
  AO22X1_RVT U3578 ( .A1(\inq_ary[7][154] ), .A2(n3322), .A3(
        \inq_ary[14][154] ), .A4(n3325), .Y(n3259) );
  AO22X1_RVT U3579 ( .A1(\inq_ary[0][154] ), .A2(n3315), .A3(\inq_ary[1][154] ), .A4(n3324), .Y(n3258) );
  AO22X1_RVT U3580 ( .A1(\inq_ary[11][154] ), .A2(n3316), .A3(
        \inq_ary[2][154] ), .A4(n3271), .Y(n3257) );
  NOR4X1_RVT U3581 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .Y(n3266)
         );
  AO22X1_RVT U3582 ( .A1(\inq_ary[13][154] ), .A2(n3323), .A3(
        \inq_ary[6][154] ), .A4(n3311), .Y(n3264) );
  AO22X1_RVT U3583 ( .A1(\inq_ary[12][154] ), .A2(n3303), .A3(
        \inq_ary[9][154] ), .A4(n3314), .Y(n3263) );
  AO22X1_RVT U3584 ( .A1(\inq_ary[10][154] ), .A2(n3326), .A3(
        \inq_ary[8][154] ), .A4(n3313), .Y(n3262) );
  AO22X1_RVT U3585 ( .A1(\inq_ary[3][154] ), .A2(n3310), .A3(
        \inq_ary[15][154] ), .A4(n3312), .Y(n3261) );
  NOR4X1_RVT U3586 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .Y(n3265)
         );
  NAND2X0_RVT U3587 ( .A1(n3266), .A2(n3265), .Y(N416) );
  AO22X1_RVT U3588 ( .A1(\inq_ary[13][155] ), .A2(n3323), .A3(
        \inq_ary[15][155] ), .A4(n3312), .Y(n3270) );
  AO22X1_RVT U3589 ( .A1(\inq_ary[14][155] ), .A2(n3325), .A3(
        \inq_ary[11][155] ), .A4(n3316), .Y(n3269) );
  AO22X1_RVT U3590 ( .A1(\inq_ary[12][155] ), .A2(n3303), .A3(
        \inq_ary[4][155] ), .A4(n3321), .Y(n3268) );
  AO22X1_RVT U3591 ( .A1(\inq_ary[10][155] ), .A2(n3326), .A3(
        \inq_ary[6][155] ), .A4(n3311), .Y(n3267) );
  NOR4X1_RVT U3592 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .Y(n3277)
         );
  AO22X1_RVT U3593 ( .A1(\inq_ary[9][155] ), .A2(n3314), .A3(\inq_ary[0][155] ), .A4(n3315), .Y(n3275) );
  AO22X1_RVT U3594 ( .A1(\inq_ary[7][155] ), .A2(n3322), .A3(\inq_ary[2][155] ), .A4(n3271), .Y(n3274) );
  AO22X1_RVT U3595 ( .A1(\inq_ary[1][155] ), .A2(n3324), .A3(\inq_ary[8][155] ), .A4(n3313), .Y(n3273) );
  AO22X1_RVT U3596 ( .A1(\inq_ary[5][155] ), .A2(n3298), .A3(\inq_ary[3][155] ), .A4(n3310), .Y(n3272) );
  NOR4X1_RVT U3597 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .Y(n3276)
         );
  NAND2X0_RVT U3598 ( .A1(n3277), .A2(n3276), .Y(N417) );
  AO22X1_RVT U3599 ( .A1(\inq_ary[5][156] ), .A2(n3298), .A3(
        \inq_ary[12][156] ), .A4(n3303), .Y(n3281) );
  AO22X1_RVT U3600 ( .A1(\inq_ary[2][156] ), .A2(n3271), .A3(\inq_ary[0][156] ), .A4(n3315), .Y(n3280) );
  AO22X1_RVT U3601 ( .A1(\inq_ary[13][156] ), .A2(n3323), .A3(
        \inq_ary[6][156] ), .A4(n3311), .Y(n3279) );
  AO22X1_RVT U3602 ( .A1(\inq_ary[3][156] ), .A2(n3310), .A3(\inq_ary[9][156] ), .A4(n3314), .Y(n3278) );
  NOR4X1_RVT U3603 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .Y(n3287)
         );
  AO22X1_RVT U3604 ( .A1(\inq_ary[14][156] ), .A2(n3325), .A3(
        \inq_ary[7][156] ), .A4(n3322), .Y(n3285) );
  AO22X1_RVT U3605 ( .A1(\inq_ary[11][156] ), .A2(n3316), .A3(
        \inq_ary[8][156] ), .A4(n3313), .Y(n3284) );
  AO22X1_RVT U3606 ( .A1(\inq_ary[4][156] ), .A2(n3321), .A3(
        \inq_ary[10][156] ), .A4(n3326), .Y(n3283) );
  AO22X1_RVT U3607 ( .A1(\inq_ary[15][156] ), .A2(n3312), .A3(
        \inq_ary[1][156] ), .A4(n3324), .Y(n3282) );
  NOR4X1_RVT U3608 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .Y(n3286)
         );
  NAND2X0_RVT U3609 ( .A1(n3287), .A2(n3286), .Y(N418) );
  AO22X1_RVT U3610 ( .A1(\inq_ary[13][157] ), .A2(n3323), .A3(
        \inq_ary[10][157] ), .A4(n3326), .Y(n3291) );
  AO22X1_RVT U3611 ( .A1(\inq_ary[11][157] ), .A2(n3316), .A3(
        \inq_ary[5][157] ), .A4(n3298), .Y(n3290) );
  AO22X1_RVT U3612 ( .A1(\inq_ary[9][157] ), .A2(n3314), .A3(\inq_ary[6][157] ), .A4(n3311), .Y(n3289) );
  AO22X1_RVT U3613 ( .A1(\inq_ary[15][157] ), .A2(n3312), .A3(
        \inq_ary[0][157] ), .A4(n3315), .Y(n3288) );
  NOR4X1_RVT U3614 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .Y(n3297)
         );
  AO22X1_RVT U3615 ( .A1(\inq_ary[8][157] ), .A2(n3313), .A3(\inq_ary[4][157] ), .A4(n3321), .Y(n3295) );
  AO22X1_RVT U3616 ( .A1(\inq_ary[3][157] ), .A2(n3310), .A3(\inq_ary[1][157] ), .A4(n3324), .Y(n3294) );
  AO22X1_RVT U3617 ( .A1(\inq_ary[14][157] ), .A2(n3325), .A3(
        \inq_ary[7][157] ), .A4(n3322), .Y(n3293) );
  AO22X1_RVT U3618 ( .A1(\inq_ary[2][157] ), .A2(n3271), .A3(
        \inq_ary[12][157] ), .A4(n3303), .Y(n3292) );
  NOR4X1_RVT U3619 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .Y(n3296)
         );
  NAND2X0_RVT U3620 ( .A1(n3297), .A2(n3296), .Y(N419) );
  AO22X1_RVT U3621 ( .A1(\inq_ary[10][158] ), .A2(n3326), .A3(
        \inq_ary[2][158] ), .A4(n3271), .Y(n3302) );
  AO22X1_RVT U3622 ( .A1(\inq_ary[7][158] ), .A2(n3322), .A3(
        \inq_ary[14][158] ), .A4(n3325), .Y(n3301) );
  AO22X1_RVT U3623 ( .A1(\inq_ary[5][158] ), .A2(n3298), .A3(\inq_ary[4][158] ), .A4(n3321), .Y(n3300) );
  AO22X1_RVT U3624 ( .A1(\inq_ary[6][158] ), .A2(n3311), .A3(\inq_ary[8][158] ), .A4(n3313), .Y(n3299) );
  NOR4X1_RVT U3625 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .Y(n3309)
         );
  AO22X1_RVT U3626 ( .A1(\inq_ary[1][158] ), .A2(n3324), .A3(
        \inq_ary[13][158] ), .A4(n3323), .Y(n3307) );
  AO22X1_RVT U3627 ( .A1(\inq_ary[11][158] ), .A2(n3316), .A3(
        \inq_ary[15][158] ), .A4(n3312), .Y(n3306) );
  AO22X1_RVT U3628 ( .A1(\inq_ary[0][158] ), .A2(n3315), .A3(\inq_ary[3][158] ), .A4(n3310), .Y(n3305) );
  AO22X1_RVT U3629 ( .A1(\inq_ary[9][158] ), .A2(n3314), .A3(
        \inq_ary[12][158] ), .A4(n3303), .Y(n3304) );
  NOR4X1_RVT U3630 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .Y(n3308)
         );
  NAND2X0_RVT U3631 ( .A1(n3309), .A2(n3308), .Y(N420) );
  AO22X1_RVT U3632 ( .A1(\inq_ary[5][159] ), .A2(n3298), .A3(\inq_ary[3][159] ), .A4(n3310), .Y(n3320) );
  AO22X1_RVT U3633 ( .A1(\inq_ary[15][159] ), .A2(n3312), .A3(
        \inq_ary[6][159] ), .A4(n3311), .Y(n3319) );
  AO22X1_RVT U3634 ( .A1(\inq_ary[9][159] ), .A2(n3314), .A3(\inq_ary[8][159] ), .A4(n3313), .Y(n3318) );
  AO22X1_RVT U3635 ( .A1(\inq_ary[11][159] ), .A2(n3316), .A3(
        \inq_ary[0][159] ), .A4(n3315), .Y(n3317) );
  NOR4X1_RVT U3636 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .Y(n3332)
         );
  AO22X1_RVT U3637 ( .A1(\inq_ary[12][159] ), .A2(n3303), .A3(
        \inq_ary[2][159] ), .A4(n3271), .Y(n3330) );
  AO22X1_RVT U3638 ( .A1(\inq_ary[7][159] ), .A2(n3322), .A3(\inq_ary[4][159] ), .A4(n3321), .Y(n3329) );
  AO22X1_RVT U3639 ( .A1(\inq_ary[1][159] ), .A2(n3324), .A3(
        \inq_ary[13][159] ), .A4(n3323), .Y(n3328) );
  AO22X1_RVT U3640 ( .A1(\inq_ary[10][159] ), .A2(n3326), .A3(
        \inq_ary[14][159] ), .A4(n3325), .Y(n3327) );
  NOR4X1_RVT U3641 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .Y(n3331)
         );
  NAND2X0_RVT U3642 ( .A1(n3332), .A2(n3331), .Y(N421) );
endmodule


module fpu ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, arst_l, grst_l, gclk, 
        cluster_cken, fp_cpx_req_cq, fp_cpx_data_ca, ctu_tst_pre_grst_l, 
        global_shift_enable, ctu_tst_scan_disable, ctu_tst_scanmode, 
        ctu_tst_macrotest, ctu_tst_short_chain, si, so );
  input [123:0] pcx_fpio_data_px2;
  output [7:0] fp_cpx_req_cq;
  output [144:0] fp_cpx_data_ca;
  input pcx_fpio_data_rdy_px2, arst_l, grst_l, gclk, cluster_cken,
         ctu_tst_pre_grst_l, global_shift_enable, ctu_tst_scan_disable,
         ctu_tst_scanmode, ctu_tst_macrotest, ctu_tst_short_chain, si;
  output so;
  wire   pcx_fpio_data_rdy_px2_buf1, a1stg_step, m1stg_step, d1stg_step,
         add_pipe_active, mul_pipe_active, div_pipe_active, sehold,
         arst_l_in_buf3, fpu_grst_l_in_buf2, rclk, fadd_clken_l, fmul_clken_l,
         fdiv_clken_l, inq_add, inq_mul, inq_div, inq_in1_exp_neq_ffs,
         inq_in1_exp_eq_0, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in2_exp_neq_ffs, inq_in2_exp_eq_0,
         inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0,
         inq_read_en, inq_we, se_in_buf3, se, rst_tri_en,
         inq_in1_50_0_neq_0_add_buf1, inq_in1_53_32_neq_0_add_buf1,
         inq_in1_exp_eq_0_add_buf1, inq_in1_exp_neq_ffs_add_buf1,
         inq_in2_50_0_neq_0_add_buf1, inq_in2_53_32_neq_0_add_buf1,
         inq_in2_exp_eq_0_add_buf1, inq_in2_exp_neq_ffs_add_buf1, add_dest_rdy,
         arst_l_add_buf4, fpu_grst_l_add_buf3, a6stg_fadd_in, a6stg_fcmpop,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         add_sign_out, se_add_exp_buf2, se_add_frac_buf2,
         inq_in1_50_0_neq_0_mul_buf1, inq_in1_53_32_neq_0_mul_buf1,
         inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_neq_ffs_mul_buf1,
         inq_in2_50_0_neq_0_mul_buf1, inq_in2_53_32_neq_0_mul_buf1,
         inq_in2_exp_eq_0_mul_buf1, inq_in2_exp_neq_ffs_mul_buf1, mul_dest_rdy,
         fmul_clken_l_buf1, arst_l_mul_buf2, fpu_grst_l_mul_buf1,
         m6stg_fmul_in, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out,
         se_mul_buf4, se_mul64_buf2, inq_in1_53_0_neq_0_div_buf1,
         inq_in1_50_0_neq_0_div_buf1, inq_in1_53_32_neq_0_div_buf1,
         inq_in1_exp_eq_0_div_buf1, inq_in1_exp_neq_ffs_div_buf1,
         inq_in2_53_0_neq_0_div_buf1, inq_in2_50_0_neq_0_div_buf1,
         inq_in2_53_32_neq_0_div_buf1, inq_in2_exp_eq_0_div_buf1,
         inq_in2_exp_neq_ffs_div_buf1, div_dest_rdy,
         fdiv_clken_l_div_frac_buf1, fdiv_clken_l_div_exp_buf1,
         arst_l_div_buf2, fpu_grst_l, d8stg_fdiv_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, se_div_buf5, arst_l_out_buf3, se_out_buf2,
         ctu_tst_pre_grst_l_buf1, global_shift_enable_buf1,
         ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1,
         ctu_tst_macrotest_buf1, ctu_tst_short_chain_buf1, scan_manual_6_buf1,
         so_unbuf, cluster_cken_buf1, arst_l_cluster_header_buf2, grst_l_buf1,
         se_cluster_header_buf2, scan_manual_6, net211169, net211170,
         net211171, net211172, net211173, net211174, net211175, net211176,
         net211177, net211178, net211179, net211180, net211181, net211182,
         net211183, net211184, net211185, net211186, net211187, net211188,
         net211189, net211190, net211191, net211192, net211193, net211194,
         net211195, net211196, net211197, net211198, net211199, net211200,
         net211201, net211202, net211203, net211204, net211205, net211206,
         net211207, net211208, net211209, net211210, net211211, net211212,
         net211213, net211214, net211215, net211216, net211217, net211218,
         net211219, net211220, net211221, net211222, net211223, net211224,
         net211225, net211226, net211227, net211228, net211229, net211230,
         net211231, net211232, net211233, net211234, net211235, net211236,
         net211237, net211238, net211239, net211240, net211241, net211242,
         net211243, net211244, net211245, net211246, net211247, net211248,
         net211249, net211250, net211251, net211252, net211253, net211254,
         net211255, net211256, net211257, net211258, net211259, net211260,
         net211261, net211262, net211263, net211264, net211265, net211266,
         net211267, net211268, net211269, net211270, net211271, net211272,
         net211273, net211274, net211275, net211276, net211277, net211278,
         net211279, net211280, net211281, net211282, net211283, net211284,
         net211285, net211286, net211287, net211288, net211289, net211290,
         net211291, net211292, net211293, net211294, net211295, net211296,
         net211297, net211298, net211299, net211300, net211301, net211302,
         net211303, net211304, net211305, net211306, net211307, net211308,
         net211309, net211310, net211311, net211312, net211313, net211314,
         net211315, net211316, net211317, net211318, net211319, net211320,
         net211321, net211322;
  wire   [123:0] pcx_fpio_data_px2_buf1;
  wire   [154:0] inq_dout;
  wire   [4:0] inq_id;
  wire   [1:0] inq_rnd_mode;
  wire   [1:0] inq_fcc;
  wire   [7:0] inq_op;
  wire   [63:0] inq_in1;
  wire   [63:0] inq_in2;
  wire   [4:0] fp_id_in;
  wire   [1:0] fp_rnd_mode_in;
  wire   [1:0] fp_fcc_in;
  wire   [7:0] fp_op_in;
  wire   [68:0] fp_src1_in;
  wire   [68:0] fp_src2_in;
  wire   [3:0] inq_rdaddr;
  wire   [3:0] inq_wraddr;
  wire   [155:0] inq_sram_din_buf1;
  wire   [7:0] inq_op_add_buf1;
  wire   [1:0] inq_rnd_mode_add_buf1;
  wire   [4:0] inq_id_add_buf1;
  wire   [63:0] inq_in1_add_buf1;
  wire   [63:0] inq_in2_add_buf1;
  wire   [9:0] add_id_out_in;
  wire   [4:0] add_exc_out;
  wire   [10:0] add_exp_out;
  wire   [63:0] add_frac_out;
  wire   [1:0] add_cc_out;
  wire   [1:0] add_fcc_out;
  wire   [7:0] inq_op_mul_buf1;
  wire   [1:0] inq_rnd_mode_mul_buf1;
  wire   [4:0] inq_id_mul_buf1;
  wire   [63:0] inq_in1_mul_buf1;
  wire   [63:0] inq_in2_mul_buf1;
  wire   [9:0] m6stg_id_in;
  wire   [4:0] mul_exc_out;
  wire   [10:0] mul_exp_out;
  wire   [51:0] mul_frac_out;
  wire   [7:0] inq_op_div_buf1;
  wire   [1:0] inq_rnd_mode_div_buf1;
  wire   [4:0] inq_id_div_buf1;
  wire   [63:0] inq_in1_div_buf1;
  wire   [63:0] inq_in2_div_buf1;
  wire   [9:0] div_id_out_in;
  wire   [4:0] div_exc_out;
  wire   [10:0] div_exp_out;
  wire   [51:0] div_frac_out;
  wire   [7:0] fp_cpx_req_cq_unbuf;
  wire   [144:0] fp_cpx_data_ca_unbuf;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178;
  assign fp_cpx_data_ca[71] = 1'b0;
  assign fp_cpx_data_ca[70] = 1'b0;
  assign fp_cpx_data_ca[64] = 1'b0;
  assign fp_cpx_data_ca[142] = 1'b0;
  assign fp_cpx_data_ca[141] = 1'b0;
  assign fp_cpx_data_ca[140] = 1'b0;
  assign fp_cpx_data_ca[136] = 1'b0;
  assign fp_cpx_data_ca[77] = 1'b0;
  assign fp_cpx_data_ca[78] = 1'b0;
  assign fp_cpx_data_ca[79] = 1'b0;
  assign fp_cpx_data_ca[80] = 1'b0;
  assign fp_cpx_data_ca[81] = 1'b0;
  assign fp_cpx_data_ca[82] = 1'b0;
  assign fp_cpx_data_ca[83] = 1'b0;
  assign fp_cpx_data_ca[84] = 1'b0;
  assign fp_cpx_data_ca[85] = 1'b0;
  assign fp_cpx_data_ca[86] = 1'b0;
  assign fp_cpx_data_ca[87] = 1'b0;
  assign fp_cpx_data_ca[88] = 1'b0;
  assign fp_cpx_data_ca[89] = 1'b0;
  assign fp_cpx_data_ca[90] = 1'b0;
  assign fp_cpx_data_ca[91] = 1'b0;
  assign fp_cpx_data_ca[92] = 1'b0;
  assign fp_cpx_data_ca[93] = 1'b0;
  assign fp_cpx_data_ca[94] = 1'b0;
  assign fp_cpx_data_ca[95] = 1'b0;
  assign fp_cpx_data_ca[96] = 1'b0;
  assign fp_cpx_data_ca[97] = 1'b0;
  assign fp_cpx_data_ca[98] = 1'b0;
  assign fp_cpx_data_ca[99] = 1'b0;
  assign fp_cpx_data_ca[100] = 1'b0;
  assign fp_cpx_data_ca[101] = 1'b0;
  assign fp_cpx_data_ca[102] = 1'b0;
  assign fp_cpx_data_ca[103] = 1'b0;
  assign fp_cpx_data_ca[104] = 1'b0;
  assign fp_cpx_data_ca[105] = 1'b0;
  assign fp_cpx_data_ca[106] = 1'b0;
  assign fp_cpx_data_ca[107] = 1'b0;
  assign fp_cpx_data_ca[108] = 1'b0;
  assign fp_cpx_data_ca[109] = 1'b0;
  assign fp_cpx_data_ca[110] = 1'b0;
  assign fp_cpx_data_ca[111] = 1'b0;
  assign fp_cpx_data_ca[112] = 1'b0;
  assign fp_cpx_data_ca[113] = 1'b0;
  assign fp_cpx_data_ca[114] = 1'b0;
  assign fp_cpx_data_ca[115] = 1'b0;
  assign fp_cpx_data_ca[116] = 1'b0;
  assign fp_cpx_data_ca[117] = 1'b0;
  assign fp_cpx_data_ca[118] = 1'b0;
  assign fp_cpx_data_ca[119] = 1'b0;
  assign fp_cpx_data_ca[120] = 1'b0;
  assign fp_cpx_data_ca[121] = 1'b0;
  assign fp_cpx_data_ca[122] = 1'b0;
  assign fp_cpx_data_ca[123] = 1'b0;
  assign fp_cpx_data_ca[124] = 1'b0;
  assign fp_cpx_data_ca[125] = 1'b0;
  assign fp_cpx_data_ca[126] = 1'b0;
  assign fp_cpx_data_ca[127] = 1'b0;
  assign fp_cpx_data_ca[128] = 1'b0;
  assign fp_cpx_data_ca[129] = 1'b0;
  assign fp_cpx_data_ca[130] = 1'b0;
  assign fp_cpx_data_ca[131] = 1'b0;
  assign fp_cpx_data_ca[132] = 1'b0;
  assign fp_cpx_data_ca[133] = 1'b0;
  assign fp_cpx_data_ca[137] = 1'b0;
  assign fp_cpx_data_ca[138] = 1'b0;
  assign fp_cpx_data_ca[139] = 1'b0;

  fpu_in fpu_in ( .pcx_fpio_data_rdy_px2(pcx_fpio_data_rdy_px2_buf1), 
        .pcx_fpio_data_px2({pcx_fpio_data_px2_buf1[123:118], net211285, 
        pcx_fpio_data_px2_buf1[116:112], net211286, net211287, net211288, 
        net211289, net211290, net211291, net211292, net211293, net211294, 
        net211295, net211296, net211297, net211298, net211299, net211300, 
        net211301, net211302, net211303, net211304, net211305, net211306, 
        net211307, net211308, net211309, net211310, net211311, net211312, 
        net211313, net211314, net211315, net211316, net211317, 
        pcx_fpio_data_px2_buf1[79:72], net211318, net211319, net211320, 
        net211321, pcx_fpio_data_px2_buf1[67:0]}), .a1stg_step(a1stg_step), 
        .m1stg_step(m1stg_step), .d1stg_step(d1stg_step), .add_pipe_active(
        add_pipe_active), .mul_pipe_active(mul_pipe_active), .div_pipe_active(
        div_pipe_active), .inq_dout(inq_dout), .sehold(sehold), .arst_l(
        arst_l_in_buf3), .grst_l(fpu_grst_l_in_buf2), .rclk(rclk), 
        .fadd_clken_l(fadd_clken_l), .fmul_clken_l(fmul_clken_l), 
        .fdiv_clken_l(fdiv_clken_l), .inq_add(inq_add), .inq_mul(inq_mul), 
        .inq_div(inq_div), .inq_id(inq_id), .inq_rnd_mode(inq_rnd_mode), 
        .inq_fcc(inq_fcc), .inq_op(inq_op), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in1_exp_eq_0(inq_in1_exp_eq_0), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1(inq_in1), .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), 
        .inq_in2_exp_eq_0(inq_in2_exp_eq_0), .inq_in2_53_0_neq_0(
        inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), .inq_in2(inq_in2), 
        .fp_id_in(fp_id_in), .fp_rnd_mode_in(fp_rnd_mode_in), .fp_fcc_in(
        fp_fcc_in), .fp_op_in(fp_op_in), .fp_src1_in(fp_src1_in), .fp_src2_in(
        fp_src2_in), .inq_rdaddr(inq_rdaddr), .inq_wraddr(inq_wraddr), 
        .inq_read_en(inq_read_en), .inq_we(inq_we), .se(se_in_buf3), .si(
        net211322) );
  bw_r_rf16x160 bw_r_rf16x160 ( .dout({inq_dout, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4}), .din({
        inq_sram_din_buf1[155:1], net211282, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .rd_adr(inq_rdaddr), .wr_adr(inq_wraddr), .read_en(inq_read_en), 
        .wr_en(inq_we), .rst_tri_en(rst_tri_en), .word_wen({1'b1, 1'b1, 1'b1, 
        1'b1}), .byte_wen({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .rd_clk(rclk), .wr_clk(rclk), .se(se), .si_r(net211283), .si_w(net211284), 
        .reset_l(arst_l_in_buf3), .sehold(sehold) );
  fpu_add fpu_add ( .inq_op(inq_op_add_buf1), .inq_rnd_mode(
        inq_rnd_mode_add_buf1), .inq_id(inq_id_add_buf1), .inq_fcc(inq_fcc), 
        .inq_in1(inq_in1_add_buf1), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0_add_buf1), .inq_in1_53_32_neq_0(
        inq_in1_53_32_neq_0_add_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_add_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_add_buf1), .inq_in2(inq_in2_add_buf1), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0_add_buf1), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0_add_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_add_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_add_buf1), .inq_add(inq_add), .fadd_clken_l(
        fadd_clken_l), .arst_l(arst_l_add_buf4), .grst_l(fpu_grst_l_add_buf3), 
        .rclk(rclk), .add_pipe_active(add_pipe_active), .a1stg_step(a1stg_step), .a6stg_fadd_in(a6stg_fadd_in), .add_id_out_in(add_id_out_in), .a6stg_fcmpop(
        a6stg_fcmpop), .add_exc_out({add_exc_out[4:2], SYNOPSYS_UNCONNECTED__5, 
        add_exc_out[0]}), .a6stg_dbl_dst(a6stg_dbl_dst), .a6stg_sng_dst(
        a6stg_sng_dst), .a6stg_long_dst(a6stg_long_dst), .a6stg_int_dst(
        a6stg_int_dst), .add_sign_out(add_sign_out), .add_exp_out(add_exp_out), 
        .add_frac_out(add_frac_out), .add_cc_out(add_cc_out), .add_fcc_out(
        add_fcc_out), .se_add_exp(se_add_exp_buf2), .se_add_frac(
        se_add_frac_buf2), .si(net211281), .add_dest_rdy_BAR(add_dest_rdy) );
  fpu_mul fpu_mul ( .inq_op(inq_op_mul_buf1), .inq_rnd_mode(
        inq_rnd_mode_mul_buf1), .inq_id(inq_id_mul_buf1), .inq_in1(
        inq_in1_mul_buf1), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0_mul_buf1), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0_mul_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_mul_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_mul_buf1), .inq_in2(inq_in2_mul_buf1), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0_mul_buf1), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0_mul_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_mul_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_mul_buf1), .inq_mul(inq_mul), .fmul_clken_l(
        fmul_clken_l), .fmul_clken_l_buf1(fmul_clken_l_buf1), .arst_l(
        arst_l_mul_buf2), .grst_l(fpu_grst_l_mul_buf1), .rclk(rclk), 
        .mul_pipe_active(mul_pipe_active), .m1stg_step(m1stg_step), 
        .m6stg_fmul_in(m6stg_fmul_in), .m6stg_id_in(m6stg_id_in), 
        .mul_exc_out({mul_exc_out[4:2], SYNOPSYS_UNCONNECTED__6, 
        mul_exc_out[0]}), .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), 
        .m6stg_fmuls(m6stg_fmuls), .mul_sign_out(mul_sign_out), .mul_exp_out(
        mul_exp_out), .mul_frac_out(mul_frac_out), .se_mul(se_mul_buf4), 
        .se_mul64(se_mul64_buf2), .si(net211280), .mul_dest_rdy_BAR(
        mul_dest_rdy), .mul_dest_rdya_BAR(mul_dest_rdy) );
  fpu_div fpu_div ( .inq_op(inq_op_div_buf1), .inq_rnd_mode(
        inq_rnd_mode_div_buf1), .inq_id(inq_id_div_buf1), .inq_in1(
        inq_in1_div_buf1), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0_div_buf1), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0_div_buf1), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0_div_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_div_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_div_buf1), .inq_in2(inq_in2_div_buf1), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0_div_buf1), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0_div_buf1), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0_div_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_div_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_div_buf1), .inq_div(inq_div), .fdiv_clken_l(
        fdiv_clken_l_div_frac_buf1), .fdiv_clken_l_div_exp_buf1(
        fdiv_clken_l_div_exp_buf1), .arst_l(arst_l_div_buf2), .grst_l(
        fpu_grst_l), .rclk(rclk), .div_pipe_active(div_pipe_active), 
        .d1stg_step(d1stg_step), .d8stg_fdiv_in(d8stg_fdiv_in), 
        .div_id_out_in(div_id_out_in), .div_exc_out(div_exc_out), 
        .d8stg_fdivd(d8stg_fdivd), .d8stg_fdivs(d8stg_fdivs), .div_sign_out(
        div_sign_out), .div_exp_outa(div_exp_out), .div_frac_outa(div_frac_out), .se(se_div_buf5), .si(net211279), .div_dest_rdy_BAR(div_dest_rdy) );
  fpu_out fpu_out ( .d8stg_fdiv_in(d8stg_fdiv_in), .m6stg_fmul_in(
        m6stg_fmul_in), .a6stg_fadd_in(a6stg_fadd_in), .div_id_out_in(
        div_id_out_in), .m6stg_id_in(m6stg_id_in), .add_id_out_in(
        add_id_out_in), .div_exc_out(div_exc_out), .d8stg_fdivd(d8stg_fdivd), 
        .d8stg_fdivs(d8stg_fdivs), .div_sign_out(div_sign_out), .div_exp_out(
        div_exp_out), .div_frac_out(div_frac_out), .mul_exc_out({
        mul_exc_out[4:2], net211276, mul_exc_out[0]}), .m6stg_fmul_dbl_dst(
        m6stg_fmul_dbl_dst), .m6stg_fmuls(m6stg_fmuls), .mul_sign_out(
        mul_sign_out), .mul_exp_out(mul_exp_out), .mul_frac_out(mul_frac_out), 
        .add_exc_out({add_exc_out[4:2], net211277, add_exc_out[0]}), 
        .a6stg_fcmpop(a6stg_fcmpop), .add_cc_out(add_cc_out), .add_fcc_out(
        add_fcc_out), .a6stg_dbl_dst(a6stg_dbl_dst), .a6stg_sng_dst(
        a6stg_sng_dst), .a6stg_long_dst(a6stg_long_dst), .a6stg_int_dst(
        a6stg_int_dst), .add_sign_out(add_sign_out), .add_exp_out(add_exp_out), 
        .add_frac_out(add_frac_out), .arst_l(arst_l_out_buf3), .grst_l(
        fpu_grst_l_add_buf3), .rclk(rclk), .fp_cpx_req_cq(fp_cpx_req_cq_unbuf), 
        .fp_cpx_data_ca({fp_cpx_data_ca_unbuf[144:143], 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, fp_cpx_data_ca_unbuf[135:134], 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, fp_cpx_data_ca_unbuf[76:72], 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        fp_cpx_data_ca_unbuf[69:65], SYNOPSYS_UNCONNECTED__73, 
        fp_cpx_data_ca_unbuf[63:0]}), .se(se_out_buf2), .si(net211278), 
        .add_dest_rdy_BAR(add_dest_rdy), .div_dest_rdy_BAR(div_dest_rdy), 
        .mul_dest_rdy_BAR(mul_dest_rdy) );
  test_stub_scan test_stub_scan ( .mem_write_disable(rst_tri_en), .sehold(
        sehold), .se(se), .so_0(so_unbuf), .ctu_tst_pre_grst_l(
        ctu_tst_pre_grst_l_buf1), .arst_l(arst_l_add_buf4), 
        .global_shift_enable(global_shift_enable_buf1), .ctu_tst_scan_disable(
        ctu_tst_scan_disable_buf1), .ctu_tst_scanmode(ctu_tst_scanmode_buf1), 
        .ctu_tst_macrotest(ctu_tst_macrotest_buf1), .ctu_tst_short_chain(
        ctu_tst_short_chain_buf1), .long_chain_so_0(scan_manual_6_buf1), 
        .short_chain_so_0(net211275), .long_chain_so_1(1'b0), 
        .short_chain_so_1(1'b0), .long_chain_so_2(1'b0), .short_chain_so_2(
        1'b0) );
  bw_clk_cl_fpu_cmp cluster_header ( .so(scan_manual_6), .cluster_grst_l(
        fpu_grst_l), .rclk(rclk), .si(net211274), .se(se_cluster_header_buf2), 
        .adbginit_l(1'b1), .gdbginit_l(1'b1), .arst_l(
        arst_l_cluster_header_buf2), .grst_l(grst_l_buf1), .cluster_cken(
        cluster_cken_buf1), .gclk(gclk) );
  fpu_rptr_groups fpu_rptr_groups ( .inq_in1(inq_in1), .inq_in2(inq_in2), 
        .inq_id(inq_id), .inq_op(inq_op), .inq_rnd_mode(inq_rnd_mode), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), .inq_in1_53_0_neq_0(
        inq_in1_53_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .ctu_tst_macrotest(
        ctu_tst_macrotest), .ctu_tst_pre_grst_l(ctu_tst_pre_grst_l), 
        .ctu_tst_scan_disable(ctu_tst_scan_disable), .ctu_tst_scanmode(
        ctu_tst_scanmode), .ctu_tst_short_chain(ctu_tst_short_chain), 
        .global_shift_enable(global_shift_enable), .grst_l(grst_l), 
        .cluster_cken(cluster_cken), .se(se), .arst_l(arst_l), .fpu_grst_l(
        fpu_grst_l), .fmul_clken_l(fmul_clken_l), .fdiv_clken_l(fdiv_clken_l), 
        .scan_manual_6(scan_manual_6), .si(net211169), .so_unbuf(so_unbuf), 
        .pcx_fpio_data_px2({pcx_fpio_data_px2[123:118], net211170, 
        pcx_fpio_data_px2[116:112], net211171, net211172, net211173, net211174, 
        net211175, net211176, net211177, net211178, net211179, net211180, 
        net211181, net211182, net211183, net211184, net211185, net211186, 
        net211187, net211188, net211189, net211190, net211191, net211192, 
        net211193, net211194, net211195, net211196, net211197, net211198, 
        net211199, net211200, net211201, net211202, pcx_fpio_data_px2[79:72], 
        net211203, net211204, net211205, net211206, pcx_fpio_data_px2[67:0]}), 
        .pcx_fpio_data_rdy_px2(pcx_fpio_data_rdy_px2), .fp_cpx_req_cq(
        fp_cpx_req_cq_unbuf), .fp_cpx_data_ca({fp_cpx_data_ca_unbuf[144:143], 
        net211207, net211208, net211209, net211210, net211211, net211212, 
        net211213, fp_cpx_data_ca_unbuf[135:134], net211214, net211215, 
        net211216, net211217, net211218, net211219, net211220, net211221, 
        net211222, net211223, net211224, net211225, net211226, net211227, 
        net211228, net211229, net211230, net211231, net211232, net211233, 
        net211234, net211235, net211236, net211237, net211238, net211239, 
        net211240, net211241, net211242, net211243, net211244, net211245, 
        net211246, net211247, net211248, net211249, net211250, net211251, 
        net211252, net211253, net211254, net211255, net211256, net211257, 
        net211258, net211259, net211260, net211261, net211262, net211263, 
        net211264, net211265, net211266, net211267, net211268, net211269, 
        net211270, fp_cpx_data_ca_unbuf[76:72], net211271, net211272, 
        fp_cpx_data_ca_unbuf[69:65], net211273, fp_cpx_data_ca_unbuf[63:0]}), 
        .inq_sram_din_unbuf({fp_id_in, fp_rnd_mode_in, fp_fcc_in, fp_op_in, 
        fp_src1_in, fp_src2_in, 1'b0}), .inq_in1_add_buf1(inq_in1_add_buf1), 
        .inq_in1_mul_buf1(inq_in1_mul_buf1), .inq_in1_div_buf1(
        inq_in1_div_buf1), .inq_in2_add_buf1(inq_in2_add_buf1), 
        .inq_in2_mul_buf1(inq_in2_mul_buf1), .inq_in2_div_buf1(
        inq_in2_div_buf1), .inq_id_add_buf1(inq_id_add_buf1), 
        .inq_id_mul_buf1(inq_id_mul_buf1), .inq_id_div_buf1(inq_id_div_buf1), 
        .inq_op_add_buf1(inq_op_add_buf1), .inq_op_div_buf1(inq_op_div_buf1), 
        .inq_op_mul_buf1(inq_op_mul_buf1), .inq_rnd_mode_add_buf1(
        inq_rnd_mode_add_buf1), .inq_rnd_mode_div_buf1(inq_rnd_mode_div_buf1), 
        .inq_rnd_mode_mul_buf1(inq_rnd_mode_mul_buf1), 
        .inq_in1_50_0_neq_0_add_buf1(inq_in1_50_0_neq_0_add_buf1), 
        .inq_in1_50_0_neq_0_mul_buf1(inq_in1_50_0_neq_0_mul_buf1), 
        .inq_in1_50_0_neq_0_div_buf1(inq_in1_50_0_neq_0_div_buf1), 
        .inq_in1_53_0_neq_0_div_buf1(inq_in1_53_0_neq_0_div_buf1), 
        .inq_in1_53_32_neq_0_add_buf1(inq_in1_53_32_neq_0_add_buf1), 
        .inq_in1_53_32_neq_0_mul_buf1(inq_in1_53_32_neq_0_mul_buf1), 
        .inq_in1_53_32_neq_0_div_buf1(inq_in1_53_32_neq_0_div_buf1), 
        .inq_in1_exp_eq_0_add_buf1(inq_in1_exp_eq_0_add_buf1), 
        .inq_in1_exp_eq_0_mul_buf1(inq_in1_exp_eq_0_mul_buf1), 
        .inq_in1_exp_eq_0_div_buf1(inq_in1_exp_eq_0_div_buf1), 
        .inq_in1_exp_neq_ffs_add_buf1(inq_in1_exp_neq_ffs_add_buf1), 
        .inq_in1_exp_neq_ffs_mul_buf1(inq_in1_exp_neq_ffs_mul_buf1), 
        .inq_in1_exp_neq_ffs_div_buf1(inq_in1_exp_neq_ffs_div_buf1), 
        .inq_in2_50_0_neq_0_add_buf1(inq_in2_50_0_neq_0_add_buf1), 
        .inq_in2_50_0_neq_0_mul_buf1(inq_in2_50_0_neq_0_mul_buf1), 
        .inq_in2_50_0_neq_0_div_buf1(inq_in2_50_0_neq_0_div_buf1), 
        .inq_in2_53_0_neq_0_div_buf1(inq_in2_53_0_neq_0_div_buf1), 
        .inq_in2_53_32_neq_0_add_buf1(inq_in2_53_32_neq_0_add_buf1), 
        .inq_in2_53_32_neq_0_mul_buf1(inq_in2_53_32_neq_0_mul_buf1), 
        .inq_in2_53_32_neq_0_div_buf1(inq_in2_53_32_neq_0_div_buf1), 
        .inq_in2_exp_eq_0_add_buf1(inq_in2_exp_eq_0_add_buf1), 
        .inq_in2_exp_eq_0_mul_buf1(inq_in2_exp_eq_0_mul_buf1), 
        .inq_in2_exp_eq_0_div_buf1(inq_in2_exp_eq_0_div_buf1), 
        .inq_in2_exp_neq_ffs_add_buf1(inq_in2_exp_neq_ffs_add_buf1), 
        .inq_in2_exp_neq_ffs_mul_buf1(inq_in2_exp_neq_ffs_mul_buf1), 
        .inq_in2_exp_neq_ffs_div_buf1(inq_in2_exp_neq_ffs_div_buf1), 
        .ctu_tst_macrotest_buf1(ctu_tst_macrotest_buf1), 
        .ctu_tst_pre_grst_l_buf1(ctu_tst_pre_grst_l_buf1), 
        .ctu_tst_scan_disable_buf1(ctu_tst_scan_disable_buf1), 
        .ctu_tst_scanmode_buf1(ctu_tst_scanmode_buf1), 
        .ctu_tst_short_chain_buf1(ctu_tst_short_chain_buf1), 
        .global_shift_enable_buf1(global_shift_enable_buf1), .grst_l_buf1(
        grst_l_buf1), .cluster_cken_buf1(cluster_cken_buf1), .se_add_exp_buf2(
        se_add_exp_buf2), .se_add_frac_buf2(se_add_frac_buf2), .se_out_buf2(
        se_out_buf2), .se_mul64_buf2(se_mul64_buf2), .se_cluster_header_buf2(
        se_cluster_header_buf2), .se_in_buf3(se_in_buf3), .se_mul_buf4(
        se_mul_buf4), .se_div_buf5(se_div_buf5), .arst_l_div_buf2(
        arst_l_div_buf2), .arst_l_mul_buf2(arst_l_mul_buf2), 
        .arst_l_cluster_header_buf2(arst_l_cluster_header_buf2), 
        .arst_l_in_buf3(arst_l_in_buf3), .arst_l_out_buf3(arst_l_out_buf3), 
        .arst_l_add_buf4(arst_l_add_buf4), .fpu_grst_l_mul_buf1(
        fpu_grst_l_mul_buf1), .fpu_grst_l_in_buf2(fpu_grst_l_in_buf2), 
        .fpu_grst_l_add_buf3(fpu_grst_l_add_buf3), .fmul_clken_l_buf1(
        fmul_clken_l_buf1), .fdiv_clken_l_div_exp_buf1(
        fdiv_clken_l_div_exp_buf1), .fdiv_clken_l_div_frac_buf1(
        fdiv_clken_l_div_frac_buf1), .scan_manual_6_buf1(scan_manual_6_buf1), 
        .so(so), .pcx_fpio_data_px2_buf1({pcx_fpio_data_px2_buf1[123:118], 
        SYNOPSYS_UNCONNECTED__74, pcx_fpio_data_px2_buf1[116:112], 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        pcx_fpio_data_px2_buf1[79:72], SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, pcx_fpio_data_px2_buf1[67:0]}), 
        .pcx_fpio_data_rdy_px2_buf1(pcx_fpio_data_rdy_px2_buf1), 
        .fp_cpx_req_cq_buf1(fp_cpx_req_cq), .fp_cpx_data_ca_buf1({
        fp_cpx_data_ca[144:143], SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        fp_cpx_data_ca[135:134], SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        fp_cpx_data_ca[76:72], SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, fp_cpx_data_ca[69:65], 
        SYNOPSYS_UNCONNECTED__177, fp_cpx_data_ca[63:0]}), .inq_sram_din_buf1(
        {inq_sram_din_buf1[155:1], SYNOPSYS_UNCONNECTED__178}) );
endmodule

