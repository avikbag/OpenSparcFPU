
module dffrl_async_SIZE1 ( din, clk, rst_l, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst_l, se;
  wire   N0, N1, N2, N3, N4;
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[0]  ( .clear(N2), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C18 ( .DATA1(si[0]), .DATA2(din[0]), .CONTROL1(N0), .CONTROL2(N1), 
        .Z(N4) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N3), .Z(N1) );
  GTECH_NOT I_0 ( .A(rst_l), .Z(N2) );
  GTECH_NOT I_1 ( .A(se), .Z(N3) );
endmodule


module dffr_SIZE1 ( din, clk, rst, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, rst, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7;
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C17 ( .DATA1(1'b0), .DATA2(din[0]), .CONTROL1(N0), .CONTROL2(N1), 
        .Z(N6) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  GTECH_BUF B_1 ( .A(N5), .Z(N1) );
  SELECT_OP C18 ( .DATA1(si[0]), .DATA2(N6), .CONTROL1(N2), .CONTROL2(N3), .Z(
        N7) );
  GTECH_BUF B_2 ( .A(se), .Z(N2) );
  GTECH_BUF B_3 ( .A(N4), .Z(N3) );
  GTECH_NOT I_0 ( .A(se), .Z(N4) );
  GTECH_NOT I_1 ( .A(rst), .Z(N5) );
endmodule


module dff_SIZE1 ( din, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input clk, se;
  wire   N0, N1, N2, N3;
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C11 ( .DATA1(si[0]), .DATA2(din[0]), .CONTROL1(N0), .CONTROL2(N1), 
        .Z(N3) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE5 ( din, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7;
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C15 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dffre_SIZE4 ( din, rst, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17;
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  SELECT_OP C42 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(din), .CONTROL1(N0), 
        .CONTROL2(N15), .Z({N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C43 ( .DATA1(si), .DATA2({N9, N8, N7, N6}), .CONTROL1(N1), 
        .CONTROL2(N2), .Z({N13, N12, N11, N10}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C51 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N14) );
  GTECH_AND2 C54 ( .A(en), .B(N14), .Z(N15) );
  GTECH_AND2 C55 ( .A(N5), .B(N3), .Z(N16) );
  GTECH_NOT I_3 ( .A(N16), .Z(N17) );
endmodule


module dff_SIZE4 ( din, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6;
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C14 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dffre_SIZE1 ( din, rst, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11;
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  SELECT_OP C27 ( .DATA1(1'b0), .DATA2(din[0]), .CONTROL1(N0), .CONTROL2(N9), 
        .Z(N6) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C28 ( .DATA1(si[0]), .DATA2(N6), .CONTROL1(N1), .CONTROL2(N2), .Z(
        N7) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C36 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N8) );
  GTECH_AND2 C39 ( .A(en), .B(N8), .Z(N9) );
  GTECH_AND2 C40 ( .A(N5), .B(N3), .Z(N10) );
  GTECH_NOT I_3 ( .A(N10), .Z(N11) );
endmodule


module dff_SIZE8 ( din, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10;
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C18 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE16 ( din, clk, q, se, si, so );
  input [15:0] din;
  output [15:0] q;
  input [15:0] si;
  output [15:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18;
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C26 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, 
        N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dffre_SIZE3 ( din, rst, en, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15;
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  SELECT_OP C37 ( .DATA1({1'b0, 1'b0, 1'b0}), .DATA2(din), .CONTROL1(N0), 
        .CONTROL2(N13), .Z({N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C38 ( .DATA1(si), .DATA2({N8, N7, N6}), .CONTROL1(N1), .CONTROL2(
        N2), .Z({N11, N10, N9}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C46 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N12) );
  GTECH_AND2 C49 ( .A(en), .B(N12), .Z(N13) );
  GTECH_AND2 C50 ( .A(N5), .B(N3), .Z(N14) );
  GTECH_NOT I_3 ( .A(N14), .Z(N15) );
endmodule


module fpu_in_ctl ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, fp_op_in, 
        fp_op_in_7in, a1stg_step, m1stg_step, d1stg_step, add_pipe_active, 
        mul_pipe_active, div_pipe_active, sehold, arst_l, grst_l, rclk, 
        fp_data_rdy, fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_we, 
        inq_wraddr, inq_read_en, inq_rdaddr, inq_bp, inq_bp_inv, inq_fwrd, 
        inq_fwrd_inv, inq_add, inq_mul, inq_div, se, si, so );
  input [123:118] pcx_fpio_data_px2;
  input [3:2] fp_op_in;
  output [3:0] inq_wraddr;
  output [3:0] inq_rdaddr;
  input pcx_fpio_data_rdy_px2, fp_op_in_7in, a1stg_step, m1stg_step,
         d1stg_step, add_pipe_active, mul_pipe_active, div_pipe_active, sehold,
         arst_l, grst_l, rclk, se, si;
  output fp_data_rdy, fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_we,
         inq_read_en, inq_bp, inq_bp_inv, inq_fwrd, inq_fwrd_inv, inq_add,
         inq_mul, inq_div, so;
  wire   in_ctl_rst_l, reset, fp_vld_in, fp_op_in_7_inv, inq_wrptr_step,
         inq_div_wrptr_step, inq_empty, inq_div_empty, inq_re, N0, inq_div_re,
         N1, inq_div_rd, valid_packet, valid_packet_dly, sehold_inv, N2,
         fp_add_in, fp_mul_in, N3, N4, N5, inq_pipe0_we, inq_pipe1_we,
         inq_pipe2_we, inq_pipe3_we, inq_pipe4_we, inq_pipe5_we, inq_pipe6_we,
         inq_pipe7_we, inq_pipe8_we, inq_pipe9_we, inq_pipe10_we,
         inq_pipe11_we, inq_pipe12_we, inq_pipe13_we, inq_pipe14_we,
         inq_pipe15_we, tag_sel, d1stg_step_dly, inq_diva_dly, inq_adda_dly,
         inq_mula_dly, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, net16642,
         net16643, net16644, net16645, net16646, net16647, net16648, net16649,
         net16650, net16651, net16652, net16653, net16654, net16655, net16656,
         net16657, net16658, net16659, net16660, net16661, net16662, net16663,
         net16664, net16665, net16666, net16667, net16668, net16669, net16670,
         net16671, net16672, net16673, net16674, net16675, net16676, net16677,
         net16678, net16679, net16680, net16681, net16682, net16683, net16684,
         net16685, net16686, net16687, net16688, net16689, net16690, net16691,
         net16692, net16693, net16694, net16695, net16696, net16697, net16698,
         net16699, net16700, net16701, net16702, net16703, net16704, net16705,
         net16706, net16707, net16708, net16709, net16710, net16711, net16712,
         net16713, net16714, net16715, net16716, net16717, net16718, net16719,
         net16720, net16721, net16722, net16723, net16724, net16725, net16726,
         net16727, net16728, net16729, net16730, net16731, net16732, net16733,
         net16734, net16735, net16736, net16737, net16738, net16739, net16740,
         net16741, net16742, net16743, net16744, net16745, net16746, net16747,
         net16748, net16749, net16750, net16751, net16752, net16753, net16754,
         net16755, net16756, net16757, net16758, net16759, net16760;
  wire   [4:0] fp_type_in;
  wire   [3:0] inq_wrptr;
  wire   [3:0] inq_wrptr_plus1;
  wire   [3:0] inq_div_wrptr;
  wire   [3:0] inq_div_wrptr_plus1;
  wire   [3:0] inq_wraddr_del;
  wire   [3:0] inq_rdptr;
  wire   [3:0] inq_rdptr_plus1;
  wire   [3:0] inq_rdptr_in;
  wire   [3:0] inq_div_rdptr;
  wire   [3:0] inq_div_rdptr_plus1;
  wire   [3:0] inq_div_rdptr_in;
  wire   [3:0] inq_rdaddr_del;
  wire   [7:0] inq_rdptr_dec;
  wire   [7:0] inq_rdptr_dec_in;
  wire   [7:0] inq_div_rdptr_dec;
  wire   [7:0] inq_div_rdptr_dec_in;
  wire   [15:0] inq_rdaddr_del_dec_in;
  wire   [15:0] inq_rdaddr_del_dec;
  wire   [2:0] inq_pipe0;
  wire   [2:0] inq_pipe1;
  wire   [2:0] inq_pipe2;
  wire   [2:0] inq_pipe3;
  wire   [2:0] inq_pipe4;
  wire   [2:0] inq_pipe5;
  wire   [2:0] inq_pipe6;
  wire   [2:0] inq_pipe7;
  wire   [2:0] inq_pipe8;
  wire   [2:0] inq_pipe9;
  wire   [2:0] inq_pipe10;
  wire   [2:0] inq_pipe11;
  wire   [2:0] inq_pipe12;
  wire   [2:0] inq_pipe13;
  wire   [2:0] inq_pipe14;
  wire   [2:0] inq_pipe15;

  dffrl_async_SIZE1 dffrl_in_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(in_ctl_rst_l), .se(se), .si(net16760) );
  dffr_SIZE1 i_fp_data_rdy ( .din(pcx_fpio_data_rdy_px2), .clk(rclk), .rst(
        reset), .q(fp_data_rdy), .se(se), .si(net16759) );
  dff_SIZE1 i_fp_vld_in ( .din(pcx_fpio_data_px2[123]), .clk(rclk), .q(
        fp_vld_in), .se(se), .si(net16758) );
  dff_SIZE5 i_fp_type_in ( .din(pcx_fpio_data_px2[122:118]), .clk(rclk), .q(
        fp_type_in), .se(se), .si({net16753, net16754, net16755, net16756, 
        net16757}) );
  dffre_SIZE4 i_inq_wrptr ( .din(inq_wrptr_plus1), .rst(reset), .en(
        inq_wrptr_step), .clk(rclk), .q(inq_wrptr), .se(se), .si({net16749, 
        net16750, net16751, net16752}) );
  dffre_SIZE4 i_inq_div_wrptr ( .din(inq_div_wrptr_plus1), .rst(reset), .en(
        inq_div_wrptr_step), .clk(rclk), .q(inq_div_wrptr), .se(se), .si({
        net16745, net16746, net16747, net16748}) );
  dff_SIZE4 i_inq_wraddr_del ( .din(inq_wraddr), .clk(rclk), .q(inq_wraddr_del), .se(se), .si({net16741, net16742, net16743, net16744}) );
  dff_SIZE4 i_inq_rdptr ( .din(inq_rdptr_in), .clk(rclk), .q(inq_rdptr), .se(
        se), .si({net16737, net16738, net16739, net16740}) );
  dff_SIZE4 i_inq_div_rdptr ( .din(inq_div_rdptr_in), .clk(rclk), .q(
        inq_div_rdptr), .se(se), .si({net16733, net16734, net16735, net16736})
         );
  dff_SIZE1 i_inq_div_rd ( .din(inq_rdaddr[3]), .clk(rclk), .q(inq_div_rd), 
        .se(se), .si(net16732) );
  dff_SIZE4 i_inq_rdaddr_del ( .din(inq_rdaddr), .clk(rclk), .q(inq_rdaddr_del), .se(se), .si({net16728, net16729, net16730, net16731}) );
  dffre_SIZE1 i_valid_packet_dly ( .din(valid_packet), .rst(reset), .en(1'b1), 
        .clk(rclk), .q(valid_packet_dly), .se(se), .si(net16727) );
  EQ_UNS_OP eq_433 ( .A(inq_wraddr_del), .B(inq_rdaddr_del), .Z(N2) );
  EQ_UNS_OP eq_437 ( .A(inq_wrptr), .B(inq_rdptr), .Z(inq_empty) );
  EQ_UNS_OP eq_439 ( .A(inq_div_wrptr), .B(inq_div_rdptr), .Z(inq_div_empty)
         );
  dff_SIZE8 i_inq_rdptr_dec ( .din(inq_rdptr_dec_in), .clk(rclk), .q(
        inq_rdptr_dec), .se(se), .si({net16719, net16720, net16721, net16722, 
        net16723, net16724, net16725, net16726}) );
  dff_SIZE8 i_inq_div_rdptr_dec ( .din(inq_div_rdptr_dec_in), .clk(rclk), .q(
        inq_div_rdptr_dec), .se(se), .si({net16711, net16712, net16713, 
        net16714, net16715, net16716, net16717, net16718}) );
  dff_SIZE16 i_inq_rdaddr_del_dec ( .din(inq_rdaddr_del_dec_in), .clk(rclk), 
        .q(inq_rdaddr_del_dec), .se(se), .si({net16695, net16696, net16697, 
        net16698, net16699, net16700, net16701, net16702, net16703, net16704, 
        net16705, net16706, net16707, net16708, net16709, net16710}) );
  dffre_SIZE3 i_inq_pipe0 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe0_we), .clk(rclk), .q(inq_pipe0), .se(se), .si({
        net16692, net16693, net16694}) );
  dffre_SIZE3 i_inq_pipe1 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe1_we), .clk(rclk), .q(inq_pipe1), .se(se), .si({
        net16689, net16690, net16691}) );
  dffre_SIZE3 i_inq_pipe2 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe2_we), .clk(rclk), .q(inq_pipe2), .se(se), .si({
        net16686, net16687, net16688}) );
  dffre_SIZE3 i_inq_pipe3 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe3_we), .clk(rclk), .q(inq_pipe3), .se(se), .si({
        net16683, net16684, net16685}) );
  dffre_SIZE3 i_inq_pipe4 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe4_we), .clk(rclk), .q(inq_pipe4), .se(se), .si({
        net16680, net16681, net16682}) );
  dffre_SIZE3 i_inq_pipe5 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe5_we), .clk(rclk), .q(inq_pipe5), .se(se), .si({
        net16677, net16678, net16679}) );
  dffre_SIZE3 i_inq_pipe6 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe6_we), .clk(rclk), .q(inq_pipe6), .se(se), .si({
        net16674, net16675, net16676}) );
  dffre_SIZE3 i_inq_pipe7 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe7_we), .clk(rclk), .q(inq_pipe7), .se(se), .si({
        net16671, net16672, net16673}) );
  dffre_SIZE3 i_inq_pipe8 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe8_we), .clk(rclk), .q(inq_pipe8), .se(se), .si({
        net16668, net16669, net16670}) );
  dffre_SIZE3 i_inq_pipe9 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), .rst(
        reset), .en(inq_pipe9_we), .clk(rclk), .q(inq_pipe9), .se(se), .si({
        net16665, net16666, net16667}) );
  dffre_SIZE3 i_inq_pipe10 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe10_we), .clk(rclk), .q(inq_pipe10), .se(se), 
        .si({net16662, net16663, net16664}) );
  dffre_SIZE3 i_inq_pipe11 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe11_we), .clk(rclk), .q(inq_pipe11), .se(se), 
        .si({net16659, net16660, net16661}) );
  dffre_SIZE3 i_inq_pipe12 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe12_we), .clk(rclk), .q(inq_pipe12), .se(se), 
        .si({net16656, net16657, net16658}) );
  dffre_SIZE3 i_inq_pipe13 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe13_we), .clk(rclk), .q(inq_pipe13), .se(se), 
        .si({net16653, net16654, net16655}) );
  dffre_SIZE3 i_inq_pipe14 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe14_we), .clk(rclk), .q(inq_pipe14), .se(se), 
        .si({net16650, net16651, net16652}) );
  dffre_SIZE3 i_inq_pipe15 ( .din({inq_wraddr[3], fp_mul_in, fp_add_in}), 
        .rst(reset), .en(inq_pipe15_we), .clk(rclk), .q(inq_pipe15), .se(se), 
        .si({net16647, net16648, net16649}) );
  dffre_SIZE1 i_inq_adda_dly ( .din(inq_add), .rst(reset), .en(1'b1), .clk(
        rclk), .q(inq_adda_dly), .se(se), .si(net16646) );
  dffre_SIZE1 i_inq_mula_dly ( .din(inq_mul), .rst(reset), .en(1'b1), .clk(
        rclk), .q(inq_mula_dly), .se(se), .si(net16645) );
  dffre_SIZE1 i_inq_diva_dly ( .din(inq_div), .rst(reset), .en(1'b1), .clk(
        rclk), .q(inq_diva_dly), .se(se), .si(net16644) );
  dffre_SIZE1 i_d1stg_step_dly ( .din(d1stg_step), .rst(reset), .en(1'b1), 
        .clk(rclk), .q(d1stg_step_dly), .se(se), .si(net16643) );
  GTECH_OR2 C97 ( .A(inq_wrptr[1]), .B(inq_wrptr[2]), .Z(N6) );
  GTECH_OR2 C98 ( .A(inq_wrptr[0]), .B(N6), .Z(N7) );
  GTECH_NOT I_0 ( .A(N7), .Z(N8) );
  GTECH_NOT I_1 ( .A(inq_wrptr[0]), .Z(N9) );
  GTECH_OR2 C101 ( .A(inq_wrptr[1]), .B(inq_wrptr[2]), .Z(N10) );
  GTECH_OR2 C102 ( .A(N9), .B(N10), .Z(N11) );
  GTECH_NOT I_2 ( .A(N11), .Z(N12) );
  GTECH_NOT I_3 ( .A(inq_wrptr[1]), .Z(N13) );
  GTECH_OR2 C105 ( .A(N13), .B(inq_wrptr[2]), .Z(N14) );
  GTECH_OR2 C106 ( .A(inq_wrptr[0]), .B(N14), .Z(N15) );
  GTECH_NOT I_4 ( .A(N15), .Z(N16) );
  GTECH_OR2 C110 ( .A(N13), .B(inq_wrptr[2]), .Z(N17) );
  GTECH_OR2 C111 ( .A(N9), .B(N17), .Z(N18) );
  GTECH_NOT I_5 ( .A(N18), .Z(N19) );
  GTECH_NOT I_6 ( .A(inq_wrptr[2]), .Z(N20) );
  GTECH_OR2 C114 ( .A(inq_wrptr[1]), .B(N20), .Z(N21) );
  GTECH_OR2 C115 ( .A(inq_wrptr[0]), .B(N21), .Z(N22) );
  GTECH_NOT I_7 ( .A(N22), .Z(N23) );
  GTECH_OR2 C119 ( .A(inq_wrptr[1]), .B(N20), .Z(N24) );
  GTECH_OR2 C120 ( .A(N9), .B(N24), .Z(N25) );
  GTECH_NOT I_8 ( .A(N25), .Z(N26) );
  GTECH_OR2 C124 ( .A(N13), .B(N20), .Z(N27) );
  GTECH_OR2 C125 ( .A(inq_wrptr[0]), .B(N27), .Z(N28) );
  GTECH_NOT I_9 ( .A(N28), .Z(N29) );
  GTECH_AND2 C127 ( .A(inq_wrptr[1]), .B(inq_wrptr[2]), .Z(N30) );
  GTECH_AND2 C128 ( .A(inq_wrptr[0]), .B(N30), .Z(N31) );
  GTECH_OR2 C129 ( .A(inq_div_wrptr[1]), .B(inq_div_wrptr[2]), .Z(N32) );
  GTECH_OR2 C130 ( .A(inq_div_wrptr[0]), .B(N32), .Z(N33) );
  GTECH_NOT I_10 ( .A(N33), .Z(N34) );
  GTECH_NOT I_11 ( .A(inq_div_wrptr[0]), .Z(N35) );
  GTECH_OR2 C133 ( .A(inq_div_wrptr[1]), .B(inq_div_wrptr[2]), .Z(N36) );
  GTECH_OR2 C134 ( .A(N35), .B(N36), .Z(N37) );
  GTECH_NOT I_12 ( .A(N37), .Z(N38) );
  GTECH_NOT I_13 ( .A(inq_div_wrptr[1]), .Z(N39) );
  GTECH_OR2 C137 ( .A(N39), .B(inq_div_wrptr[2]), .Z(N40) );
  GTECH_OR2 C138 ( .A(inq_div_wrptr[0]), .B(N40), .Z(N41) );
  GTECH_NOT I_14 ( .A(N41), .Z(N42) );
  GTECH_OR2 C142 ( .A(N39), .B(inq_div_wrptr[2]), .Z(N43) );
  GTECH_OR2 C143 ( .A(N35), .B(N43), .Z(N44) );
  GTECH_NOT I_15 ( .A(N44), .Z(N45) );
  GTECH_NOT I_16 ( .A(inq_div_wrptr[2]), .Z(N46) );
  GTECH_OR2 C146 ( .A(inq_div_wrptr[1]), .B(N46), .Z(N47) );
  GTECH_OR2 C147 ( .A(inq_div_wrptr[0]), .B(N47), .Z(N48) );
  GTECH_NOT I_17 ( .A(N48), .Z(N49) );
  GTECH_OR2 C151 ( .A(inq_div_wrptr[1]), .B(N46), .Z(N50) );
  GTECH_OR2 C152 ( .A(N35), .B(N50), .Z(N51) );
  GTECH_NOT I_18 ( .A(N51), .Z(N52) );
  GTECH_OR2 C156 ( .A(N39), .B(N46), .Z(N53) );
  GTECH_OR2 C157 ( .A(inq_div_wrptr[0]), .B(N53), .Z(N54) );
  GTECH_NOT I_19 ( .A(N54), .Z(N55) );
  GTECH_AND2 C159 ( .A(inq_div_wrptr[1]), .B(inq_div_wrptr[2]), .Z(N56) );
  GTECH_AND2 C160 ( .A(inq_div_wrptr[0]), .B(N56), .Z(N57) );
  GTECH_NOT I_20 ( .A(fp_type_in[3]), .Z(N58) );
  GTECH_NOT I_21 ( .A(fp_type_in[1]), .Z(N59) );
  GTECH_OR2 C163 ( .A(N58), .B(fp_type_in[4]), .Z(N60) );
  GTECH_OR2 C164 ( .A(fp_type_in[2]), .B(N60), .Z(N61) );
  GTECH_OR2 C165 ( .A(N59), .B(N61), .Z(N62) );
  GTECH_OR2 C166 ( .A(fp_type_in[0]), .B(N62), .Z(N63) );
  GTECH_NOT I_22 ( .A(N63), .Z(N64) );
  GTECH_NOT I_23 ( .A(fp_type_in[0]), .Z(N65) );
  GTECH_OR2 C171 ( .A(N58), .B(fp_type_in[4]), .Z(N66) );
  GTECH_OR2 C172 ( .A(fp_type_in[2]), .B(N66), .Z(N67) );
  GTECH_OR2 C173 ( .A(N59), .B(N67), .Z(N68) );
  GTECH_OR2 C174 ( .A(N65), .B(N68), .Z(N69) );
  GTECH_NOT I_24 ( .A(N69), .Z(N70) );
  GTECH_OR2 C178 ( .A(N58), .B(fp_type_in[4]), .Z(N71) );
  GTECH_OR2 C179 ( .A(fp_type_in[2]), .B(N71), .Z(N72) );
  GTECH_OR2 C180 ( .A(N59), .B(N72), .Z(N73) );
  GTECH_OR2 C181 ( .A(fp_type_in[0]), .B(N73), .Z(N74) );
  GTECH_NOT I_25 ( .A(N74), .Z(N75) );
  GTECH_OR2 C186 ( .A(N58), .B(fp_type_in[4]), .Z(N76) );
  GTECH_OR2 C187 ( .A(fp_type_in[2]), .B(N76), .Z(N77) );
  GTECH_OR2 C188 ( .A(N59), .B(N77), .Z(N78) );
  GTECH_OR2 C189 ( .A(N65), .B(N78), .Z(N79) );
  GTECH_NOT I_26 ( .A(N79), .Z(N80) );
  GTECH_OR2 C193 ( .A(N58), .B(fp_type_in[4]), .Z(N81) );
  GTECH_OR2 C194 ( .A(fp_type_in[2]), .B(N81), .Z(N82) );
  GTECH_OR2 C195 ( .A(N59), .B(N82), .Z(N83) );
  GTECH_NOT I_27 ( .A(N83), .Z(N84) );
  GTECH_OR2 C200 ( .A(N58), .B(fp_type_in[4]), .Z(N85) );
  GTECH_OR2 C201 ( .A(fp_type_in[2]), .B(N85), .Z(N86) );
  GTECH_OR2 C202 ( .A(N59), .B(N86), .Z(N87) );
  GTECH_OR2 C203 ( .A(N65), .B(N87), .Z(N88) );
  GTECH_NOT I_28 ( .A(N88), .Z(N89) );
  GTECH_NOT I_29 ( .A(fp_op_in[3]), .Z(N90) );
  GTECH_OR2 C206 ( .A(fp_op_in[2]), .B(N90), .Z(N91) );
  GTECH_NOT I_30 ( .A(N91), .Z(N92) );
  GTECH_OR2 C211 ( .A(N58), .B(fp_type_in[4]), .Z(N93) );
  GTECH_OR2 C212 ( .A(fp_type_in[2]), .B(N93), .Z(N94) );
  GTECH_OR2 C213 ( .A(N59), .B(N94), .Z(N95) );
  GTECH_OR2 C214 ( .A(N65), .B(N95), .Z(N96) );
  GTECH_NOT I_31 ( .A(N96), .Z(N97) );
  GTECH_AND2 C216 ( .A(fp_op_in[2]), .B(fp_op_in[3]), .Z(N98) );
  ADD_UNS_OP add_278 ( .A(inq_wrptr), .B(1'b1), .Z(inq_wrptr_plus1) );
  ADD_UNS_OP add_295 ( .A(inq_div_wrptr), .B(1'b1), .Z(inq_div_wrptr_plus1) );
  ADD_UNS_OP add_334 ( .A(inq_rdptr), .B(1'b1), .Z(inq_rdptr_plus1) );
  ADD_UNS_OP add_354 ( .A(inq_div_rdptr), .B(1'b1), .Z(inq_div_rdptr_plus1) );
  GTECH_NOT I_32 ( .A(in_ctl_rst_l), .Z(reset) );
  GTECH_NOT I_33 ( .A(fp_op_in_7in), .Z(fp_op_in_7_inv) );
  GTECH_AND2 C220 ( .A(N99), .B(N102), .Z(inq_we) );
  GTECH_AND2 C221 ( .A(fp_data_rdy), .B(fp_vld_in), .Z(N99) );
  GTECH_OR2 C222 ( .A(N100), .B(N101), .Z(N102) );
  GTECH_AND2 C223 ( .A(N64), .B(fp_op_in_7in), .Z(N100) );
  GTECH_AND2 C224 ( .A(N70), .B(fp_op_in_7_inv), .Z(N101) );
  GTECH_AND2 C225 ( .A(inq_we), .B(N103), .Z(inq_wrptr_step) );
  GTECH_NOT I_34 ( .A(inq_wraddr[3]), .Z(N103) );
  GTECH_AND2 C227 ( .A(inq_we), .B(inq_wraddr[3]), .Z(inq_div_wrptr_step) );
  GTECH_OR2 C228 ( .A(N104), .B(N106), .Z(inq_wraddr[2]) );
  GTECH_AND2 C229 ( .A(inq_wraddr[3]), .B(inq_div_wrptr[2]), .Z(N104) );
  GTECH_AND2 C230 ( .A(N105), .B(inq_wrptr[2]), .Z(N106) );
  GTECH_NOT I_35 ( .A(inq_wraddr[3]), .Z(N105) );
  GTECH_OR2 C232 ( .A(N107), .B(N109), .Z(inq_wraddr[1]) );
  GTECH_AND2 C233 ( .A(inq_wraddr[3]), .B(inq_div_wrptr[1]), .Z(N107) );
  GTECH_AND2 C234 ( .A(N108), .B(inq_wrptr[1]), .Z(N109) );
  GTECH_NOT I_36 ( .A(inq_wraddr[3]), .Z(N108) );
  GTECH_OR2 C236 ( .A(N110), .B(N112), .Z(inq_wraddr[0]) );
  GTECH_AND2 C237 ( .A(inq_wraddr[3]), .B(inq_div_wrptr[0]), .Z(N110) );
  GTECH_AND2 C238 ( .A(N111), .B(inq_wrptr[0]), .Z(N112) );
  GTECH_NOT I_37 ( .A(inq_wraddr[3]), .Z(N111) );
  GTECH_OR2 C240 ( .A(N113), .B(N114), .Z(inq_read_en) );
  GTECH_NOT I_38 ( .A(inq_empty), .Z(N113) );
  GTECH_NOT I_39 ( .A(inq_div_empty), .Z(N114) );
  GTECH_OR2 C243 ( .A(N115), .B(N116), .Z(inq_re) );
  GTECH_AND2 C244 ( .A(inq_add), .B(a1stg_step), .Z(N115) );
  GTECH_AND2 C245 ( .A(inq_mul), .B(m1stg_step), .Z(N116) );
  GTECH_NOT I_40 ( .A(reset), .Z(N0) );
  GTECH_OR2 C247 ( .A(N118), .B(N121), .Z(inq_rdptr_in[3]) );
  GTECH_AND2 C248 ( .A(N117), .B(inq_rdptr_plus1[3]), .Z(N118) );
  GTECH_AND2 C249 ( .A(inq_re), .B(N0), .Z(N117) );
  GTECH_AND2 C250 ( .A(N120), .B(inq_rdptr[3]), .Z(N121) );
  GTECH_AND2 C251 ( .A(N119), .B(N0), .Z(N120) );
  GTECH_NOT I_41 ( .A(inq_re), .Z(N119) );
  GTECH_OR2 C253 ( .A(N123), .B(N125), .Z(inq_rdptr_in[2]) );
  GTECH_AND2 C254 ( .A(N122), .B(inq_rdptr_plus1[2]), .Z(N123) );
  GTECH_AND2 C255 ( .A(inq_re), .B(N0), .Z(N122) );
  GTECH_AND2 C256 ( .A(N124), .B(inq_rdptr[2]), .Z(N125) );
  GTECH_AND2 C257 ( .A(N119), .B(N0), .Z(N124) );
  GTECH_OR2 C259 ( .A(N127), .B(N129), .Z(inq_rdptr_in[1]) );
  GTECH_AND2 C260 ( .A(N126), .B(inq_rdptr_plus1[1]), .Z(N127) );
  GTECH_AND2 C261 ( .A(inq_re), .B(N0), .Z(N126) );
  GTECH_AND2 C262 ( .A(N128), .B(inq_rdptr[1]), .Z(N129) );
  GTECH_AND2 C263 ( .A(N119), .B(N0), .Z(N128) );
  GTECH_OR2 C265 ( .A(N131), .B(N133), .Z(inq_rdptr_in[0]) );
  GTECH_AND2 C266 ( .A(N130), .B(inq_rdptr_plus1[0]), .Z(N131) );
  GTECH_AND2 C267 ( .A(inq_re), .B(N0), .Z(N130) );
  GTECH_AND2 C268 ( .A(N132), .B(inq_rdptr[0]), .Z(N133) );
  GTECH_AND2 C269 ( .A(N119), .B(N0), .Z(N132) );
  GTECH_AND2 C271 ( .A(inq_div), .B(d1stg_step), .Z(inq_div_re) );
  GTECH_NOT I_42 ( .A(reset), .Z(N1) );
  GTECH_OR2 C273 ( .A(N135), .B(N138), .Z(inq_div_rdptr_in[3]) );
  GTECH_AND2 C274 ( .A(N134), .B(inq_div_rdptr_plus1[3]), .Z(N135) );
  GTECH_AND2 C275 ( .A(inq_div_re), .B(N1), .Z(N134) );
  GTECH_AND2 C276 ( .A(N137), .B(inq_div_rdptr[3]), .Z(N138) );
  GTECH_AND2 C277 ( .A(N136), .B(N1), .Z(N137) );
  GTECH_NOT I_43 ( .A(inq_div_re), .Z(N136) );
  GTECH_OR2 C279 ( .A(N140), .B(N142), .Z(inq_div_rdptr_in[2]) );
  GTECH_AND2 C280 ( .A(N139), .B(inq_div_rdptr_plus1[2]), .Z(N140) );
  GTECH_AND2 C281 ( .A(inq_div_re), .B(N1), .Z(N139) );
  GTECH_AND2 C282 ( .A(N141), .B(inq_div_rdptr[2]), .Z(N142) );
  GTECH_AND2 C283 ( .A(N136), .B(N1), .Z(N141) );
  GTECH_OR2 C285 ( .A(N144), .B(N146), .Z(inq_div_rdptr_in[1]) );
  GTECH_AND2 C286 ( .A(N143), .B(inq_div_rdptr_plus1[1]), .Z(N144) );
  GTECH_AND2 C287 ( .A(inq_div_re), .B(N1), .Z(N143) );
  GTECH_AND2 C288 ( .A(N145), .B(inq_div_rdptr[1]), .Z(N146) );
  GTECH_AND2 C289 ( .A(N136), .B(N1), .Z(N145) );
  GTECH_OR2 C291 ( .A(N148), .B(N150), .Z(inq_div_rdptr_in[0]) );
  GTECH_AND2 C292 ( .A(N147), .B(inq_div_rdptr_plus1[0]), .Z(N148) );
  GTECH_AND2 C293 ( .A(inq_div_re), .B(N1), .Z(N147) );
  GTECH_AND2 C294 ( .A(N149), .B(inq_div_rdptr[0]), .Z(N150) );
  GTECH_AND2 C295 ( .A(N136), .B(N1), .Z(N149) );
  GTECH_AND2 C297 ( .A(N151), .B(N152), .Z(inq_rdaddr[3]) );
  GTECH_AND2 C298 ( .A(N114), .B(d1stg_step), .Z(N151) );
  GTECH_NOT I_44 ( .A(inq_div), .Z(N152) );
  GTECH_OR2 C301 ( .A(N155), .B(N157), .Z(inq_rdaddr[2]) );
  GTECH_AND2 C302 ( .A(inq_rdaddr[3]), .B(N154), .Z(N155) );
  GTECH_AND2 C303 ( .A(inq_div_rdptr[2]), .B(N153), .Z(N154) );
  GTECH_NOT I_45 ( .A(reset), .Z(N153) );
  GTECH_AND2 C305 ( .A(N156), .B(inq_rdptr_in[2]), .Z(N157) );
  GTECH_NOT I_46 ( .A(inq_rdaddr[3]), .Z(N156) );
  GTECH_OR2 C307 ( .A(N160), .B(N162), .Z(inq_rdaddr[1]) );
  GTECH_AND2 C308 ( .A(inq_rdaddr[3]), .B(N159), .Z(N160) );
  GTECH_AND2 C309 ( .A(inq_div_rdptr[1]), .B(N158), .Z(N159) );
  GTECH_NOT I_47 ( .A(reset), .Z(N158) );
  GTECH_AND2 C311 ( .A(N161), .B(inq_rdptr_in[1]), .Z(N162) );
  GTECH_NOT I_48 ( .A(inq_rdaddr[3]), .Z(N161) );
  GTECH_OR2 C313 ( .A(N165), .B(N167), .Z(inq_rdaddr[0]) );
  GTECH_AND2 C314 ( .A(inq_rdaddr[3]), .B(N164), .Z(N165) );
  GTECH_AND2 C315 ( .A(inq_div_rdptr[0]), .B(N163), .Z(N164) );
  GTECH_NOT I_49 ( .A(reset), .Z(N163) );
  GTECH_AND2 C317 ( .A(N166), .B(inq_rdptr_in[0]), .Z(N167) );
  GTECH_NOT I_50 ( .A(inq_rdaddr[3]), .Z(N166) );
  GTECH_AND2 C319 ( .A(N168), .B(N169), .Z(valid_packet) );
  GTECH_AND2 C320 ( .A(fp_data_rdy), .B(fp_vld_in), .Z(N168) );
  GTECH_OR2 C321 ( .A(N75), .B(N80), .Z(N169) );
  GTECH_NOT I_51 ( .A(sehold), .Z(sehold_inv) );
  GTECH_AND2 C323 ( .A(N170), .B(sehold_inv), .Z(inq_bp) );
  GTECH_AND2 C324 ( .A(N2), .B(valid_packet_dly), .Z(N170) );
  GTECH_NOT I_52 ( .A(inq_bp), .Z(inq_bp_inv) );
  GTECH_AND2 C326 ( .A(N176), .B(sehold_inv), .Z(inq_fwrd) );
  GTECH_AND2 C327 ( .A(N175), .B(valid_packet), .Z(N176) );
  GTECH_OR2 C328 ( .A(N172), .B(N174), .Z(N175) );
  GTECH_AND2 C329 ( .A(inq_empty), .B(N171), .Z(N172) );
  GTECH_NOT I_53 ( .A(inq_div_rd), .Z(N171) );
  GTECH_AND2 C331 ( .A(N173), .B(d1stg_step), .Z(N174) );
  GTECH_AND2 C332 ( .A(inq_div_empty), .B(inq_wraddr[3]), .Z(N173) );
  GTECH_NOT I_54 ( .A(inq_fwrd), .Z(inq_fwrd_inv) );
  GTECH_AND2 C334 ( .A(N178), .B(N182), .Z(fp_add_in) );
  GTECH_AND2 C335 ( .A(N177), .B(N84), .Z(N178) );
  GTECH_AND2 C336 ( .A(fp_data_rdy), .B(fp_vld_in), .Z(N177) );
  GTECH_OR2 C337 ( .A(N179), .B(N181), .Z(N182) );
  GTECH_AND2 C338 ( .A(fp_op_in_7in), .B(N65), .Z(N179) );
  GTECH_AND2 C340 ( .A(N180), .B(fp_type_in[0]), .Z(N181) );
  GTECH_AND2 C341 ( .A(fp_op_in_7_inv), .B(N90), .Z(N180) );
  GTECH_AND2 C343 ( .A(N185), .B(N92), .Z(fp_mul_in) );
  GTECH_AND2 C344 ( .A(N184), .B(fp_op_in_7_inv), .Z(N185) );
  GTECH_AND2 C345 ( .A(N183), .B(N89), .Z(N184) );
  GTECH_AND2 C346 ( .A(fp_data_rdy), .B(fp_vld_in), .Z(N183) );
  GTECH_AND2 C347 ( .A(N188), .B(N98), .Z(inq_wraddr[3]) );
  GTECH_AND2 C348 ( .A(N187), .B(fp_op_in_7_inv), .Z(N188) );
  GTECH_AND2 C349 ( .A(N186), .B(N97), .Z(N187) );
  GTECH_AND2 C350 ( .A(fp_data_rdy), .B(fp_vld_in), .Z(N186) );
  GTECH_NOT I_55 ( .A(reset), .Z(N3) );
  GTECH_OR2 C352 ( .A(N190), .B(N192), .Z(inq_rdptr_dec_in[7]) );
  GTECH_AND2 C353 ( .A(N189), .B(inq_rdptr_dec[6]), .Z(N190) );
  GTECH_AND2 C354 ( .A(inq_re), .B(N3), .Z(N189) );
  GTECH_AND2 C355 ( .A(N191), .B(inq_rdptr_dec[7]), .Z(N192) );
  GTECH_AND2 C356 ( .A(N119), .B(N3), .Z(N191) );
  GTECH_OR2 C358 ( .A(N194), .B(N196), .Z(inq_rdptr_dec_in[6]) );
  GTECH_AND2 C359 ( .A(N193), .B(inq_rdptr_dec[5]), .Z(N194) );
  GTECH_AND2 C360 ( .A(inq_re), .B(N3), .Z(N193) );
  GTECH_AND2 C361 ( .A(N195), .B(inq_rdptr_dec[6]), .Z(N196) );
  GTECH_AND2 C362 ( .A(N119), .B(N3), .Z(N195) );
  GTECH_OR2 C364 ( .A(N198), .B(N200), .Z(inq_rdptr_dec_in[5]) );
  GTECH_AND2 C365 ( .A(N197), .B(inq_rdptr_dec[4]), .Z(N198) );
  GTECH_AND2 C366 ( .A(inq_re), .B(N3), .Z(N197) );
  GTECH_AND2 C367 ( .A(N199), .B(inq_rdptr_dec[5]), .Z(N200) );
  GTECH_AND2 C368 ( .A(N119), .B(N3), .Z(N199) );
  GTECH_OR2 C370 ( .A(N202), .B(N204), .Z(inq_rdptr_dec_in[4]) );
  GTECH_AND2 C371 ( .A(N201), .B(inq_rdptr_dec[3]), .Z(N202) );
  GTECH_AND2 C372 ( .A(inq_re), .B(N3), .Z(N201) );
  GTECH_AND2 C373 ( .A(N203), .B(inq_rdptr_dec[4]), .Z(N204) );
  GTECH_AND2 C374 ( .A(N119), .B(N3), .Z(N203) );
  GTECH_OR2 C376 ( .A(N206), .B(N208), .Z(inq_rdptr_dec_in[3]) );
  GTECH_AND2 C377 ( .A(N205), .B(inq_rdptr_dec[2]), .Z(N206) );
  GTECH_AND2 C378 ( .A(inq_re), .B(N3), .Z(N205) );
  GTECH_AND2 C379 ( .A(N207), .B(inq_rdptr_dec[3]), .Z(N208) );
  GTECH_AND2 C380 ( .A(N119), .B(N3), .Z(N207) );
  GTECH_OR2 C382 ( .A(N210), .B(N212), .Z(inq_rdptr_dec_in[2]) );
  GTECH_AND2 C383 ( .A(N209), .B(inq_rdptr_dec[1]), .Z(N210) );
  GTECH_AND2 C384 ( .A(inq_re), .B(N3), .Z(N209) );
  GTECH_AND2 C385 ( .A(N211), .B(inq_rdptr_dec[2]), .Z(N212) );
  GTECH_AND2 C386 ( .A(N119), .B(N3), .Z(N211) );
  GTECH_OR2 C388 ( .A(N214), .B(N216), .Z(inq_rdptr_dec_in[1]) );
  GTECH_AND2 C389 ( .A(N213), .B(inq_rdptr_dec[0]), .Z(N214) );
  GTECH_AND2 C390 ( .A(inq_re), .B(N3), .Z(N213) );
  GTECH_AND2 C391 ( .A(N215), .B(inq_rdptr_dec[1]), .Z(N216) );
  GTECH_AND2 C392 ( .A(N119), .B(N3), .Z(N215) );
  GTECH_OR2 C394 ( .A(N219), .B(N221), .Z(inq_rdptr_dec_in[0]) );
  GTECH_OR2 C395 ( .A(reset), .B(N218), .Z(N219) );
  GTECH_AND2 C396 ( .A(N217), .B(inq_rdptr_dec[7]), .Z(N218) );
  GTECH_AND2 C397 ( .A(inq_re), .B(N3), .Z(N217) );
  GTECH_AND2 C398 ( .A(N220), .B(inq_rdptr_dec[0]), .Z(N221) );
  GTECH_AND2 C399 ( .A(N119), .B(N3), .Z(N220) );
  GTECH_NOT I_56 ( .A(reset), .Z(N4) );
  GTECH_OR2 C402 ( .A(N223), .B(N225), .Z(inq_div_rdptr_dec_in[7]) );
  GTECH_AND2 C403 ( .A(N222), .B(inq_div_rdptr_dec[6]), .Z(N223) );
  GTECH_AND2 C404 ( .A(inq_div_re), .B(N4), .Z(N222) );
  GTECH_AND2 C405 ( .A(N224), .B(inq_div_rdptr_dec[7]), .Z(N225) );
  GTECH_AND2 C406 ( .A(N136), .B(N4), .Z(N224) );
  GTECH_OR2 C408 ( .A(N227), .B(N229), .Z(inq_div_rdptr_dec_in[6]) );
  GTECH_AND2 C409 ( .A(N226), .B(inq_div_rdptr_dec[5]), .Z(N227) );
  GTECH_AND2 C410 ( .A(inq_div_re), .B(N4), .Z(N226) );
  GTECH_AND2 C411 ( .A(N228), .B(inq_div_rdptr_dec[6]), .Z(N229) );
  GTECH_AND2 C412 ( .A(N136), .B(N4), .Z(N228) );
  GTECH_OR2 C414 ( .A(N231), .B(N233), .Z(inq_div_rdptr_dec_in[5]) );
  GTECH_AND2 C415 ( .A(N230), .B(inq_div_rdptr_dec[4]), .Z(N231) );
  GTECH_AND2 C416 ( .A(inq_div_re), .B(N4), .Z(N230) );
  GTECH_AND2 C417 ( .A(N232), .B(inq_div_rdptr_dec[5]), .Z(N233) );
  GTECH_AND2 C418 ( .A(N136), .B(N4), .Z(N232) );
  GTECH_OR2 C420 ( .A(N235), .B(N237), .Z(inq_div_rdptr_dec_in[4]) );
  GTECH_AND2 C421 ( .A(N234), .B(inq_div_rdptr_dec[3]), .Z(N235) );
  GTECH_AND2 C422 ( .A(inq_div_re), .B(N4), .Z(N234) );
  GTECH_AND2 C423 ( .A(N236), .B(inq_div_rdptr_dec[4]), .Z(N237) );
  GTECH_AND2 C424 ( .A(N136), .B(N4), .Z(N236) );
  GTECH_OR2 C426 ( .A(N239), .B(N241), .Z(inq_div_rdptr_dec_in[3]) );
  GTECH_AND2 C427 ( .A(N238), .B(inq_div_rdptr_dec[2]), .Z(N239) );
  GTECH_AND2 C428 ( .A(inq_div_re), .B(N4), .Z(N238) );
  GTECH_AND2 C429 ( .A(N240), .B(inq_div_rdptr_dec[3]), .Z(N241) );
  GTECH_AND2 C430 ( .A(N136), .B(N4), .Z(N240) );
  GTECH_OR2 C432 ( .A(N243), .B(N245), .Z(inq_div_rdptr_dec_in[2]) );
  GTECH_AND2 C433 ( .A(N242), .B(inq_div_rdptr_dec[1]), .Z(N243) );
  GTECH_AND2 C434 ( .A(inq_div_re), .B(N4), .Z(N242) );
  GTECH_AND2 C435 ( .A(N244), .B(inq_div_rdptr_dec[2]), .Z(N245) );
  GTECH_AND2 C436 ( .A(N136), .B(N4), .Z(N244) );
  GTECH_OR2 C438 ( .A(N247), .B(N249), .Z(inq_div_rdptr_dec_in[1]) );
  GTECH_AND2 C439 ( .A(N246), .B(inq_div_rdptr_dec[0]), .Z(N247) );
  GTECH_AND2 C440 ( .A(inq_div_re), .B(N4), .Z(N246) );
  GTECH_AND2 C441 ( .A(N248), .B(inq_div_rdptr_dec[1]), .Z(N249) );
  GTECH_AND2 C442 ( .A(N136), .B(N4), .Z(N248) );
  GTECH_OR2 C444 ( .A(N252), .B(N254), .Z(inq_div_rdptr_dec_in[0]) );
  GTECH_OR2 C445 ( .A(reset), .B(N251), .Z(N252) );
  GTECH_AND2 C446 ( .A(N250), .B(inq_div_rdptr_dec[7]), .Z(N251) );
  GTECH_AND2 C447 ( .A(inq_div_re), .B(N4), .Z(N250) );
  GTECH_AND2 C448 ( .A(N253), .B(inq_div_rdptr_dec[0]), .Z(N254) );
  GTECH_AND2 C449 ( .A(N136), .B(N4), .Z(N253) );
  GTECH_AND2 C451 ( .A(N255), .B(N256), .Z(N5) );
  GTECH_AND2 C452 ( .A(N114), .B(d1stg_step), .Z(N255) );
  GTECH_NOT I_57 ( .A(inq_div), .Z(N256) );
  GTECH_AND2 C455 ( .A(N5), .B(N258), .Z(inq_rdaddr_del_dec_in[15]) );
  GTECH_AND2 C456 ( .A(inq_div_rdptr_dec[7]), .B(N257), .Z(N258) );
  GTECH_NOT I_58 ( .A(reset), .Z(N257) );
  GTECH_AND2 C458 ( .A(N5), .B(N260), .Z(inq_rdaddr_del_dec_in[14]) );
  GTECH_AND2 C459 ( .A(inq_div_rdptr_dec[6]), .B(N259), .Z(N260) );
  GTECH_NOT I_59 ( .A(reset), .Z(N259) );
  GTECH_AND2 C461 ( .A(N5), .B(N262), .Z(inq_rdaddr_del_dec_in[13]) );
  GTECH_AND2 C462 ( .A(inq_div_rdptr_dec[5]), .B(N261), .Z(N262) );
  GTECH_NOT I_60 ( .A(reset), .Z(N261) );
  GTECH_AND2 C464 ( .A(N5), .B(N264), .Z(inq_rdaddr_del_dec_in[12]) );
  GTECH_AND2 C465 ( .A(inq_div_rdptr_dec[4]), .B(N263), .Z(N264) );
  GTECH_NOT I_61 ( .A(reset), .Z(N263) );
  GTECH_AND2 C467 ( .A(N5), .B(N266), .Z(inq_rdaddr_del_dec_in[11]) );
  GTECH_AND2 C468 ( .A(inq_div_rdptr_dec[3]), .B(N265), .Z(N266) );
  GTECH_NOT I_62 ( .A(reset), .Z(N265) );
  GTECH_AND2 C470 ( .A(N5), .B(N268), .Z(inq_rdaddr_del_dec_in[10]) );
  GTECH_AND2 C471 ( .A(inq_div_rdptr_dec[2]), .B(N267), .Z(N268) );
  GTECH_NOT I_63 ( .A(reset), .Z(N267) );
  GTECH_AND2 C473 ( .A(N5), .B(N270), .Z(inq_rdaddr_del_dec_in[9]) );
  GTECH_AND2 C474 ( .A(inq_div_rdptr_dec[1]), .B(N269), .Z(N270) );
  GTECH_NOT I_64 ( .A(reset), .Z(N269) );
  GTECH_AND2 C476 ( .A(N5), .B(N271), .Z(inq_rdaddr_del_dec_in[8]) );
  GTECH_OR2 C477 ( .A(inq_div_rdptr_dec[0]), .B(reset), .Z(N271) );
  GTECH_AND2 C478 ( .A(N272), .B(inq_rdptr_dec_in[7]), .Z(
        inq_rdaddr_del_dec_in[7]) );
  GTECH_NOT I_65 ( .A(N5), .Z(N272) );
  GTECH_AND2 C480 ( .A(N272), .B(inq_rdptr_dec_in[6]), .Z(
        inq_rdaddr_del_dec_in[6]) );
  GTECH_AND2 C482 ( .A(N272), .B(inq_rdptr_dec_in[5]), .Z(
        inq_rdaddr_del_dec_in[5]) );
  GTECH_AND2 C484 ( .A(N272), .B(inq_rdptr_dec_in[4]), .Z(
        inq_rdaddr_del_dec_in[4]) );
  GTECH_AND2 C486 ( .A(N272), .B(inq_rdptr_dec_in[3]), .Z(
        inq_rdaddr_del_dec_in[3]) );
  GTECH_AND2 C488 ( .A(N272), .B(inq_rdptr_dec_in[2]), .Z(
        inq_rdaddr_del_dec_in[2]) );
  GTECH_AND2 C490 ( .A(N272), .B(inq_rdptr_dec_in[1]), .Z(
        inq_rdaddr_del_dec_in[1]) );
  GTECH_AND2 C492 ( .A(N272), .B(inq_rdptr_dec_in[0]), .Z(
        inq_rdaddr_del_dec_in[0]) );
  GTECH_AND2 C494 ( .A(N274), .B(N8), .Z(inq_pipe0_we) );
  GTECH_AND2 C495 ( .A(inq_we), .B(N273), .Z(N274) );
  GTECH_NOT I_66 ( .A(inq_wraddr[3]), .Z(N273) );
  GTECH_AND2 C497 ( .A(N276), .B(N12), .Z(inq_pipe1_we) );
  GTECH_AND2 C498 ( .A(inq_we), .B(N275), .Z(N276) );
  GTECH_NOT I_67 ( .A(inq_wraddr[3]), .Z(N275) );
  GTECH_AND2 C500 ( .A(N278), .B(N16), .Z(inq_pipe2_we) );
  GTECH_AND2 C501 ( .A(inq_we), .B(N277), .Z(N278) );
  GTECH_NOT I_68 ( .A(inq_wraddr[3]), .Z(N277) );
  GTECH_AND2 C503 ( .A(N280), .B(N19), .Z(inq_pipe3_we) );
  GTECH_AND2 C504 ( .A(inq_we), .B(N279), .Z(N280) );
  GTECH_NOT I_69 ( .A(inq_wraddr[3]), .Z(N279) );
  GTECH_AND2 C506 ( .A(N282), .B(N23), .Z(inq_pipe4_we) );
  GTECH_AND2 C507 ( .A(inq_we), .B(N281), .Z(N282) );
  GTECH_NOT I_70 ( .A(inq_wraddr[3]), .Z(N281) );
  GTECH_AND2 C509 ( .A(N284), .B(N26), .Z(inq_pipe5_we) );
  GTECH_AND2 C510 ( .A(inq_we), .B(N283), .Z(N284) );
  GTECH_NOT I_71 ( .A(inq_wraddr[3]), .Z(N283) );
  GTECH_AND2 C512 ( .A(N286), .B(N29), .Z(inq_pipe6_we) );
  GTECH_AND2 C513 ( .A(inq_we), .B(N285), .Z(N286) );
  GTECH_NOT I_72 ( .A(inq_wraddr[3]), .Z(N285) );
  GTECH_AND2 C515 ( .A(N288), .B(N31), .Z(inq_pipe7_we) );
  GTECH_AND2 C516 ( .A(inq_we), .B(N287), .Z(N288) );
  GTECH_NOT I_73 ( .A(inq_wraddr[3]), .Z(N287) );
  GTECH_AND2 C518 ( .A(N289), .B(N34), .Z(inq_pipe8_we) );
  GTECH_AND2 C519 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N289) );
  GTECH_AND2 C520 ( .A(N290), .B(N38), .Z(inq_pipe9_we) );
  GTECH_AND2 C521 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N290) );
  GTECH_AND2 C522 ( .A(N291), .B(N42), .Z(inq_pipe10_we) );
  GTECH_AND2 C523 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N291) );
  GTECH_AND2 C524 ( .A(N292), .B(N45), .Z(inq_pipe11_we) );
  GTECH_AND2 C525 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N292) );
  GTECH_AND2 C526 ( .A(N293), .B(N49), .Z(inq_pipe12_we) );
  GTECH_AND2 C527 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N293) );
  GTECH_AND2 C528 ( .A(N294), .B(N52), .Z(inq_pipe13_we) );
  GTECH_AND2 C529 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N294) );
  GTECH_AND2 C530 ( .A(N295), .B(N55), .Z(inq_pipe14_we) );
  GTECH_AND2 C531 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N295) );
  GTECH_AND2 C532 ( .A(N296), .B(N57), .Z(inq_pipe15_we) );
  GTECH_AND2 C533 ( .A(inq_we), .B(inq_wraddr[3]), .Z(N296) );
  GTECH_OR2 C534 ( .A(N297), .B(N301), .Z(tag_sel) );
  GTECH_AND2 C535 ( .A(inq_empty), .B(N171), .Z(N297) );
  GTECH_AND2 C537 ( .A(N300), .B(d1stg_step), .Z(N301) );
  GTECH_AND2 C538 ( .A(N299), .B(fp_vld_in), .Z(N300) );
  GTECH_AND2 C539 ( .A(N298), .B(fp_data_rdy), .Z(N299) );
  GTECH_AND2 C540 ( .A(inq_div_empty), .B(inq_wraddr[3]), .Z(N298) );
  GTECH_OR2 C541 ( .A(N309), .B(N342), .Z(inq_div) );
  GTECH_AND2 C542 ( .A(tag_sel), .B(N308), .Z(N309) );
  GTECH_AND2 C543 ( .A(N306), .B(N307), .Z(N308) );
  GTECH_AND2 C544 ( .A(N305), .B(d1stg_step_dly), .Z(N306) );
  GTECH_AND2 C545 ( .A(N304), .B(d1stg_step), .Z(N305) );
  GTECH_AND2 C546 ( .A(N303), .B(fp_vld_in), .Z(N304) );
  GTECH_AND2 C547 ( .A(N302), .B(fp_data_rdy), .Z(N303) );
  GTECH_AND2 C548 ( .A(inq_div_empty), .B(inq_wraddr[3]), .Z(N302) );
  GTECH_NOT I_74 ( .A(inq_diva_dly), .Z(N307) );
  GTECH_AND2 C550 ( .A(N310), .B(N341), .Z(N342) );
  GTECH_NOT I_75 ( .A(tag_sel), .Z(N310) );
  GTECH_OR2 C552 ( .A(N339), .B(N340), .Z(N341) );
  GTECH_OR2 C553 ( .A(N337), .B(N338), .Z(N339) );
  GTECH_OR2 C554 ( .A(N335), .B(N336), .Z(N337) );
  GTECH_OR2 C555 ( .A(N333), .B(N334), .Z(N335) );
  GTECH_OR2 C556 ( .A(N331), .B(N332), .Z(N333) );
  GTECH_OR2 C557 ( .A(N329), .B(N330), .Z(N331) );
  GTECH_OR2 C558 ( .A(N327), .B(N328), .Z(N329) );
  GTECH_OR2 C559 ( .A(N325), .B(N326), .Z(N327) );
  GTECH_OR2 C560 ( .A(N323), .B(N324), .Z(N325) );
  GTECH_OR2 C561 ( .A(N321), .B(N322), .Z(N323) );
  GTECH_OR2 C562 ( .A(N319), .B(N320), .Z(N321) );
  GTECH_OR2 C563 ( .A(N317), .B(N318), .Z(N319) );
  GTECH_OR2 C564 ( .A(N315), .B(N316), .Z(N317) );
  GTECH_OR2 C565 ( .A(N313), .B(N314), .Z(N315) );
  GTECH_OR2 C566 ( .A(N311), .B(N312), .Z(N313) );
  GTECH_AND2 C567 ( .A(inq_rdaddr_del_dec[0]), .B(inq_pipe0[2]), .Z(N311) );
  GTECH_AND2 C568 ( .A(inq_rdaddr_del_dec[1]), .B(inq_pipe1[2]), .Z(N312) );
  GTECH_AND2 C569 ( .A(inq_rdaddr_del_dec[2]), .B(inq_pipe2[2]), .Z(N314) );
  GTECH_AND2 C570 ( .A(inq_rdaddr_del_dec[3]), .B(inq_pipe3[2]), .Z(N316) );
  GTECH_AND2 C571 ( .A(inq_rdaddr_del_dec[4]), .B(inq_pipe4[2]), .Z(N318) );
  GTECH_AND2 C572 ( .A(inq_rdaddr_del_dec[5]), .B(inq_pipe5[2]), .Z(N320) );
  GTECH_AND2 C573 ( .A(inq_rdaddr_del_dec[6]), .B(inq_pipe6[2]), .Z(N322) );
  GTECH_AND2 C574 ( .A(inq_rdaddr_del_dec[7]), .B(inq_pipe7[2]), .Z(N324) );
  GTECH_AND2 C575 ( .A(inq_rdaddr_del_dec[8]), .B(inq_pipe8[2]), .Z(N326) );
  GTECH_AND2 C576 ( .A(inq_rdaddr_del_dec[9]), .B(inq_pipe9[2]), .Z(N328) );
  GTECH_AND2 C577 ( .A(inq_rdaddr_del_dec[10]), .B(inq_pipe10[2]), .Z(N330) );
  GTECH_AND2 C578 ( .A(inq_rdaddr_del_dec[11]), .B(inq_pipe11[2]), .Z(N332) );
  GTECH_AND2 C579 ( .A(inq_rdaddr_del_dec[12]), .B(inq_pipe12[2]), .Z(N334) );
  GTECH_AND2 C580 ( .A(inq_rdaddr_del_dec[13]), .B(inq_pipe13[2]), .Z(N336) );
  GTECH_AND2 C581 ( .A(inq_rdaddr_del_dec[14]), .B(inq_pipe14[2]), .Z(N338) );
  GTECH_AND2 C582 ( .A(inq_rdaddr_del_dec[15]), .B(inq_pipe15[2]), .Z(N340) );
  GTECH_OR2 C583 ( .A(N343), .B(N375), .Z(inq_mul) );
  GTECH_AND2 C584 ( .A(tag_sel), .B(fp_mul_in), .Z(N343) );
  GTECH_AND2 C585 ( .A(N310), .B(N374), .Z(N375) );
  GTECH_OR2 C587 ( .A(N372), .B(N373), .Z(N374) );
  GTECH_OR2 C588 ( .A(N370), .B(N371), .Z(N372) );
  GTECH_OR2 C589 ( .A(N368), .B(N369), .Z(N370) );
  GTECH_OR2 C590 ( .A(N366), .B(N367), .Z(N368) );
  GTECH_OR2 C591 ( .A(N364), .B(N365), .Z(N366) );
  GTECH_OR2 C592 ( .A(N362), .B(N363), .Z(N364) );
  GTECH_OR2 C593 ( .A(N360), .B(N361), .Z(N362) );
  GTECH_OR2 C594 ( .A(N358), .B(N359), .Z(N360) );
  GTECH_OR2 C595 ( .A(N356), .B(N357), .Z(N358) );
  GTECH_OR2 C596 ( .A(N354), .B(N355), .Z(N356) );
  GTECH_OR2 C597 ( .A(N352), .B(N353), .Z(N354) );
  GTECH_OR2 C598 ( .A(N350), .B(N351), .Z(N352) );
  GTECH_OR2 C599 ( .A(N348), .B(N349), .Z(N350) );
  GTECH_OR2 C600 ( .A(N346), .B(N347), .Z(N348) );
  GTECH_OR2 C601 ( .A(N344), .B(N345), .Z(N346) );
  GTECH_AND2 C602 ( .A(inq_rdaddr_del_dec[0]), .B(inq_pipe0[1]), .Z(N344) );
  GTECH_AND2 C603 ( .A(inq_rdaddr_del_dec[1]), .B(inq_pipe1[1]), .Z(N345) );
  GTECH_AND2 C604 ( .A(inq_rdaddr_del_dec[2]), .B(inq_pipe2[1]), .Z(N347) );
  GTECH_AND2 C605 ( .A(inq_rdaddr_del_dec[3]), .B(inq_pipe3[1]), .Z(N349) );
  GTECH_AND2 C606 ( .A(inq_rdaddr_del_dec[4]), .B(inq_pipe4[1]), .Z(N351) );
  GTECH_AND2 C607 ( .A(inq_rdaddr_del_dec[5]), .B(inq_pipe5[1]), .Z(N353) );
  GTECH_AND2 C608 ( .A(inq_rdaddr_del_dec[6]), .B(inq_pipe6[1]), .Z(N355) );
  GTECH_AND2 C609 ( .A(inq_rdaddr_del_dec[7]), .B(inq_pipe7[1]), .Z(N357) );
  GTECH_AND2 C610 ( .A(inq_rdaddr_del_dec[8]), .B(inq_pipe8[1]), .Z(N359) );
  GTECH_AND2 C611 ( .A(inq_rdaddr_del_dec[9]), .B(inq_pipe9[1]), .Z(N361) );
  GTECH_AND2 C612 ( .A(inq_rdaddr_del_dec[10]), .B(inq_pipe10[1]), .Z(N363) );
  GTECH_AND2 C613 ( .A(inq_rdaddr_del_dec[11]), .B(inq_pipe11[1]), .Z(N365) );
  GTECH_AND2 C614 ( .A(inq_rdaddr_del_dec[12]), .B(inq_pipe12[1]), .Z(N367) );
  GTECH_AND2 C615 ( .A(inq_rdaddr_del_dec[13]), .B(inq_pipe13[1]), .Z(N369) );
  GTECH_AND2 C616 ( .A(inq_rdaddr_del_dec[14]), .B(inq_pipe14[1]), .Z(N371) );
  GTECH_AND2 C617 ( .A(inq_rdaddr_del_dec[15]), .B(inq_pipe15[1]), .Z(N373) );
  GTECH_OR2 C618 ( .A(N376), .B(N408), .Z(inq_add) );
  GTECH_AND2 C619 ( .A(tag_sel), .B(fp_add_in), .Z(N376) );
  GTECH_AND2 C620 ( .A(N310), .B(N407), .Z(N408) );
  GTECH_OR2 C622 ( .A(N405), .B(N406), .Z(N407) );
  GTECH_OR2 C623 ( .A(N403), .B(N404), .Z(N405) );
  GTECH_OR2 C624 ( .A(N401), .B(N402), .Z(N403) );
  GTECH_OR2 C625 ( .A(N399), .B(N400), .Z(N401) );
  GTECH_OR2 C626 ( .A(N397), .B(N398), .Z(N399) );
  GTECH_OR2 C627 ( .A(N395), .B(N396), .Z(N397) );
  GTECH_OR2 C628 ( .A(N393), .B(N394), .Z(N395) );
  GTECH_OR2 C629 ( .A(N391), .B(N392), .Z(N393) );
  GTECH_OR2 C630 ( .A(N389), .B(N390), .Z(N391) );
  GTECH_OR2 C631 ( .A(N387), .B(N388), .Z(N389) );
  GTECH_OR2 C632 ( .A(N385), .B(N386), .Z(N387) );
  GTECH_OR2 C633 ( .A(N383), .B(N384), .Z(N385) );
  GTECH_OR2 C634 ( .A(N381), .B(N382), .Z(N383) );
  GTECH_OR2 C635 ( .A(N379), .B(N380), .Z(N381) );
  GTECH_OR2 C636 ( .A(N377), .B(N378), .Z(N379) );
  GTECH_AND2 C637 ( .A(inq_rdaddr_del_dec[0]), .B(inq_pipe0[0]), .Z(N377) );
  GTECH_AND2 C638 ( .A(inq_rdaddr_del_dec[1]), .B(inq_pipe1[0]), .Z(N378) );
  GTECH_AND2 C639 ( .A(inq_rdaddr_del_dec[2]), .B(inq_pipe2[0]), .Z(N380) );
  GTECH_AND2 C640 ( .A(inq_rdaddr_del_dec[3]), .B(inq_pipe3[0]), .Z(N382) );
  GTECH_AND2 C641 ( .A(inq_rdaddr_del_dec[4]), .B(inq_pipe4[0]), .Z(N384) );
  GTECH_AND2 C642 ( .A(inq_rdaddr_del_dec[5]), .B(inq_pipe5[0]), .Z(N386) );
  GTECH_AND2 C643 ( .A(inq_rdaddr_del_dec[6]), .B(inq_pipe6[0]), .Z(N388) );
  GTECH_AND2 C644 ( .A(inq_rdaddr_del_dec[7]), .B(inq_pipe7[0]), .Z(N390) );
  GTECH_AND2 C645 ( .A(inq_rdaddr_del_dec[8]), .B(inq_pipe8[0]), .Z(N392) );
  GTECH_AND2 C646 ( .A(inq_rdaddr_del_dec[9]), .B(inq_pipe9[0]), .Z(N394) );
  GTECH_AND2 C647 ( .A(inq_rdaddr_del_dec[10]), .B(inq_pipe10[0]), .Z(N396) );
  GTECH_AND2 C648 ( .A(inq_rdaddr_del_dec[11]), .B(inq_pipe11[0]), .Z(N398) );
  GTECH_AND2 C649 ( .A(inq_rdaddr_del_dec[12]), .B(inq_pipe12[0]), .Z(N400) );
  GTECH_AND2 C650 ( .A(inq_rdaddr_del_dec[13]), .B(inq_pipe13[0]), .Z(N402) );
  GTECH_AND2 C651 ( .A(inq_rdaddr_del_dec[14]), .B(inq_pipe14[0]), .Z(N404) );
  GTECH_AND2 C652 ( .A(inq_rdaddr_del_dec[15]), .B(inq_pipe15[0]), .Z(N406) );
  GTECH_NOT I_76 ( .A(N411), .Z(fadd_clken_l) );
  GTECH_OR2 C654 ( .A(N410), .B(reset), .Z(N411) );
  GTECH_OR2 C655 ( .A(N409), .B(inq_adda_dly), .Z(N410) );
  GTECH_OR2 C656 ( .A(add_pipe_active), .B(inq_add), .Z(N409) );
  GTECH_NOT I_77 ( .A(N414), .Z(fmul_clken_l) );
  GTECH_OR2 C658 ( .A(N413), .B(reset), .Z(N414) );
  GTECH_OR2 C659 ( .A(N412), .B(inq_mula_dly), .Z(N413) );
  GTECH_OR2 C660 ( .A(mul_pipe_active), .B(inq_mul), .Z(N412) );
  GTECH_NOT I_78 ( .A(N417), .Z(fdiv_clken_l) );
  GTECH_OR2 C662 ( .A(N416), .B(reset), .Z(N417) );
  GTECH_OR2 C663 ( .A(N415), .B(inq_diva_dly), .Z(N416) );
  GTECH_OR2 C664 ( .A(div_pipe_active), .B(inq_div), .Z(N415) );
endmodule


module clken_buf ( clk, rclk, enb_l, tmb_l );
  input rclk, enb_l, tmb_l;
  output clk;
  wire   N0, N1, clken, N2, N3;

  \**SEQGEN**  clken_reg ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N1), .enable(N0), .Q(clken), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b0)
         );
  GTECH_NOT I_0 ( .A(rclk), .Z(N0) );
  GTECH_OR2 C18 ( .A(N2), .B(N3), .Z(N1) );
  GTECH_NOT I_1 ( .A(enb_l), .Z(N2) );
  GTECH_NOT I_2 ( .A(tmb_l), .Z(N3) );
  GTECH_AND2 C21 ( .A(clken), .B(rclk), .Z(clk) );
endmodule


module dff_SIZE2 ( din, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4;
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C12 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE64 ( din, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66;
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C74 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dffe_SIZE69 ( din, en, clk, q, se, si, so );
  input [68:0] din;
  output [68:0] q;
  input [68:0] si;
  output [68:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74;
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N74) );
  SELECT_OP C291 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C299 ( .A(N3), .B(N2), .Z(N73) );
  GTECH_NOT I_2 ( .A(N73), .Z(N74) );
endmodule


module dff_SIZE155 ( din, clk, q, se, si, so );
  input [154:0] din;
  output [154:0] q;
  input [154:0] si;
  output [154:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157;
  assign so[154] = q[154];
  assign so[153] = q[153];
  assign so[152] = q[152];
  assign so[151] = q[151];
  assign so[150] = q[150];
  assign so[149] = q[149];
  assign so[148] = q[148];
  assign so[147] = q[147];
  assign so[146] = q[146];
  assign so[145] = q[145];
  assign so[144] = q[144];
  assign so[143] = q[143];
  assign so[142] = q[142];
  assign so[141] = q[141];
  assign so[140] = q[140];
  assign so[139] = q[139];
  assign so[138] = q[138];
  assign so[137] = q[137];
  assign so[136] = q[136];
  assign so[135] = q[135];
  assign so[134] = q[134];
  assign so[133] = q[133];
  assign so[132] = q[132];
  assign so[131] = q[131];
  assign so[130] = q[130];
  assign so[129] = q[129];
  assign so[128] = q[128];
  assign so[127] = q[127];
  assign so[126] = q[126];
  assign so[125] = q[125];
  assign so[124] = q[124];
  assign so[123] = q[123];
  assign so[122] = q[122];
  assign so[121] = q[121];
  assign so[120] = q[120];
  assign so[119] = q[119];
  assign so[118] = q[118];
  assign so[117] = q[117];
  assign so[116] = q[116];
  assign so[115] = q[115];
  assign so[114] = q[114];
  assign so[113] = q[113];
  assign so[112] = q[112];
  assign so[111] = q[111];
  assign so[110] = q[110];
  assign so[109] = q[109];
  assign so[108] = q[108];
  assign so[107] = q[107];
  assign so[106] = q[106];
  assign so[105] = q[105];
  assign so[104] = q[104];
  assign so[103] = q[103];
  assign so[102] = q[102];
  assign so[101] = q[101];
  assign so[100] = q[100];
  assign so[99] = q[99];
  assign so[98] = q[98];
  assign so[97] = q[97];
  assign so[96] = q[96];
  assign so[95] = q[95];
  assign so[94] = q[94];
  assign so[93] = q[93];
  assign so[92] = q[92];
  assign so[91] = q[91];
  assign so[90] = q[90];
  assign so[89] = q[89];
  assign so[88] = q[88];
  assign so[87] = q[87];
  assign so[86] = q[86];
  assign so[85] = q[85];
  assign so[84] = q[84];
  assign so[83] = q[83];
  assign so[82] = q[82];
  assign so[81] = q[81];
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[154]  ( .clear(1'b0), .preset(1'b0), .next_state(N157), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[154]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[153]  ( .clear(1'b0), .preset(1'b0), .next_state(N156), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[153]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[152]  ( .clear(1'b0), .preset(1'b0), .next_state(N155), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[152]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[151]  ( .clear(1'b0), .preset(1'b0), .next_state(N154), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[151]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[150]  ( .clear(1'b0), .preset(1'b0), .next_state(N153), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[150]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[149]  ( .clear(1'b0), .preset(1'b0), .next_state(N152), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[149]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[148]  ( .clear(1'b0), .preset(1'b0), .next_state(N151), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[148]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[147]  ( .clear(1'b0), .preset(1'b0), .next_state(N150), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[147]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[146]  ( .clear(1'b0), .preset(1'b0), .next_state(N149), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[146]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[145]  ( .clear(1'b0), .preset(1'b0), .next_state(N148), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[145]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[144]  ( .clear(1'b0), .preset(1'b0), .next_state(N147), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[144]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[143]  ( .clear(1'b0), .preset(1'b0), .next_state(N146), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[143]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[142]  ( .clear(1'b0), .preset(1'b0), .next_state(N145), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[142]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[141]  ( .clear(1'b0), .preset(1'b0), .next_state(N144), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[141]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[140]  ( .clear(1'b0), .preset(1'b0), .next_state(N143), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[140]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[139]  ( .clear(1'b0), .preset(1'b0), .next_state(N142), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[139]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[138]  ( .clear(1'b0), .preset(1'b0), .next_state(N141), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[138]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[137]  ( .clear(1'b0), .preset(1'b0), .next_state(N140), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[137]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[136]  ( .clear(1'b0), .preset(1'b0), .next_state(N139), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[136]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[135]  ( .clear(1'b0), .preset(1'b0), .next_state(N138), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[135]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[134]  ( .clear(1'b0), .preset(1'b0), .next_state(N137), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[134]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[133]  ( .clear(1'b0), .preset(1'b0), .next_state(N136), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[133]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[132]  ( .clear(1'b0), .preset(1'b0), .next_state(N135), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[132]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[131]  ( .clear(1'b0), .preset(1'b0), .next_state(N134), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[131]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[130]  ( .clear(1'b0), .preset(1'b0), .next_state(N133), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[130]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[129]  ( .clear(1'b0), .preset(1'b0), .next_state(N132), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[129]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[128]  ( .clear(1'b0), .preset(1'b0), .next_state(N131), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[128]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[127]  ( .clear(1'b0), .preset(1'b0), .next_state(N130), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[127]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[126]  ( .clear(1'b0), .preset(1'b0), .next_state(N129), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[126]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[125]  ( .clear(1'b0), .preset(1'b0), .next_state(N128), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[125]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[124]  ( .clear(1'b0), .preset(1'b0), .next_state(N127), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[124]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[123]  ( .clear(1'b0), .preset(1'b0), .next_state(N126), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[123]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[122]  ( .clear(1'b0), .preset(1'b0), .next_state(N125), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[122]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[121]  ( .clear(1'b0), .preset(1'b0), .next_state(N124), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[121]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[120]  ( .clear(1'b0), .preset(1'b0), .next_state(N123), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[120]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[119]  ( .clear(1'b0), .preset(1'b0), .next_state(N122), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[119]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[118]  ( .clear(1'b0), .preset(1'b0), .next_state(N121), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[118]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[117]  ( .clear(1'b0), .preset(1'b0), .next_state(N120), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[117]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[116]  ( .clear(1'b0), .preset(1'b0), .next_state(N119), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[116]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[115]  ( .clear(1'b0), .preset(1'b0), .next_state(N118), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[115]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[114]  ( .clear(1'b0), .preset(1'b0), .next_state(N117), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[114]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[113]  ( .clear(1'b0), .preset(1'b0), .next_state(N116), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[113]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[112]  ( .clear(1'b0), .preset(1'b0), .next_state(N115), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[112]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[111]  ( .clear(1'b0), .preset(1'b0), .next_state(N114), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[111]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[110]  ( .clear(1'b0), .preset(1'b0), .next_state(N113), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[110]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[109]  ( .clear(1'b0), .preset(1'b0), .next_state(N112), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[109]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[108]  ( .clear(1'b0), .preset(1'b0), .next_state(N111), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[108]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[107]  ( .clear(1'b0), .preset(1'b0), .next_state(N110), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[107]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[106]  ( .clear(1'b0), .preset(1'b0), .next_state(N109), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[106]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[105]  ( .clear(1'b0), .preset(1'b0), .next_state(N108), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[105]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[104]  ( .clear(1'b0), .preset(1'b0), .next_state(N107), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[104]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[103]  ( .clear(1'b0), .preset(1'b0), .next_state(N106), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[103]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[102]  ( .clear(1'b0), .preset(1'b0), .next_state(N105), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[102]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[101]  ( .clear(1'b0), .preset(1'b0), .next_state(N104), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[101]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[100]  ( .clear(1'b0), .preset(1'b0), .next_state(N103), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[100]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[99]  ( .clear(1'b0), .preset(1'b0), .next_state(N102), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[98]  ( .clear(1'b0), .preset(1'b0), .next_state(N101), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[97]  ( .clear(1'b0), .preset(1'b0), .next_state(N100), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(N99), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(N98), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(N97), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(N96), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(N95), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(N94), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(N93), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(N92), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(N91), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(N90), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(N89), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(N88), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(N87), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(N86), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(N85), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C165 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module fpu_in_dp ( fp_data_rdy, fpio_data_px2_116_112, fpio_data_px2_79_72, 
        fpio_data_px2_67_0, inq_fwrd, inq_fwrd_inv, inq_bp, inq_bp_inv, 
        inq_dout, rclk, fp_op_in_7in, inq_id, inq_rnd_mode, inq_fcc, inq_op, 
        inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1, inq_in2_exp_neq_ffs, 
        inq_in2_exp_eq_0, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2, fp_id_in, fp_rnd_mode_in, fp_fcc_in, 
        fp_op_in, fp_src1_in, fp_src2_in, se, si, so );
  input [116:112] fpio_data_px2_116_112;
  input [79:72] fpio_data_px2_79_72;
  input [67:0] fpio_data_px2_67_0;
  input [154:0] inq_dout;
  output [4:0] inq_id;
  output [1:0] inq_rnd_mode;
  output [1:0] inq_fcc;
  output [7:0] inq_op;
  output [63:0] inq_in1;
  output [63:0] inq_in2;
  output [4:0] fp_id_in;
  output [1:0] fp_rnd_mode_in;
  output [1:0] fp_fcc_in;
  output [7:0] fp_op_in;
  output [68:0] fp_src1_in;
  output [68:0] fp_src2_in;
  input fp_data_rdy, inq_fwrd, inq_fwrd_inv, inq_bp, inq_bp_inv, rclk, se, si;
  output fp_op_in_7in, inq_in1_exp_neq_ffs, inq_in1_exp_eq_0,
         inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in2_exp_neq_ffs, inq_in2_exp_eq_0, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, so;
  wire   se_l, clk, fp_op_in_7_inv, fp_srca_53_0_neq_0, fp_srca_50_0_neq_0,
         fp_srca_53_32_neq_0, fp_srca_exp_eq_0, fp_srca_exp_neq_ffs, N0, N1,
         N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694,
         N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705,
         N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716,
         N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936,
         N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947,
         N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980,
         N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991,
         N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002,
         N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012,
         N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022,
         N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032,
         N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042,
         N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052,
         N1053, N1054, N1055, N1056, N1057, net16336, net16337, net16338,
         net16339, net16340, net16341, net16342, net16343, net16344, net16345,
         net16346, net16347, net16348, net16349, net16350, net16351, net16352,
         net16353, net16354, net16355, net16356, net16357, net16358, net16359,
         net16360, net16361, net16362, net16363, net16364, net16365, net16366,
         net16367, net16368, net16369, net16370, net16371, net16372, net16373,
         net16374, net16375, net16376, net16377, net16378, net16379, net16380,
         net16381, net16382, net16383, net16384, net16385, net16386, net16387,
         net16388, net16389, net16390, net16391, net16392, net16393, net16394,
         net16395, net16396, net16397, net16398, net16399, net16400, net16401,
         net16402, net16403, net16404, net16405, net16406, net16407, net16408,
         net16409, net16410, net16411, net16412, net16413, net16414, net16415,
         net16416, net16417, net16418, net16419, net16420, net16421, net16422,
         net16423, net16424, net16425, net16426, net16427, net16428, net16429,
         net16430, net16431, net16432, net16433, net16434, net16435, net16436,
         net16437, net16438, net16439, net16440, net16441, net16442, net16443,
         net16444, net16445, net16446, net16447, net16448, net16449, net16450,
         net16451, net16452, net16453, net16454, net16455, net16456, net16457,
         net16458, net16459, net16460, net16461, net16462, net16463, net16464,
         net16465, net16466, net16467, net16468, net16469, net16470, net16471,
         net16472, net16473, net16474, net16475, net16476, net16477, net16478,
         net16479, net16480, net16481, net16482, net16483, net16484, net16485,
         net16486, net16487, net16488, net16489, net16490, net16491, net16492,
         net16493, net16494, net16495, net16496, net16497, net16498, net16499,
         net16500, net16501, net16502, net16503, net16504, net16505, net16506,
         net16507, net16508, net16509, net16510, net16511, net16512, net16513,
         net16514, net16515, net16516, net16517, net16518, net16519, net16520,
         net16521, net16522, net16523, net16524, net16525, net16526, net16527,
         net16528, net16529, net16530, net16531, net16532, net16533, net16534,
         net16535, net16536, net16537, net16538, net16539, net16540, net16541,
         net16542, net16543, net16544, net16545, net16546, net16547, net16548,
         net16549, net16550, net16551, net16552, net16553, net16554, net16555,
         net16556, net16557, net16558, net16559, net16560, net16561, net16562,
         net16563, net16564, net16565, net16566, net16567, net16568, net16569,
         net16570, net16571, net16572, net16573, net16574, net16575, net16576,
         net16577, net16578, net16579, net16580, net16581, net16582, net16583,
         net16584, net16585, net16586, net16587, net16588, net16589, net16590,
         net16591, net16592, net16593, net16594, net16595, net16596, net16597,
         net16598, net16599, net16600, net16601, net16602, net16603, net16604,
         net16605, net16606, net16607, net16608, net16609, net16610, net16611,
         net16612, net16613, net16614, net16615, net16616, net16617, net16618,
         net16619, net16620, net16621, net16622, net16623, net16624, net16625,
         net16626, net16627, net16628, net16629, net16630, net16631, net16632,
         net16633, net16634, net16635, net16636, net16637, net16638, net16639,
         net16640, net16641;
  wire   [63:0] fp_srca_in;
  wire   [68:0] fp_srcb_in;
  wire   [154:0] inq_din_d1;
  assign fp_op_in_7in = fp_op_in[7];

  clken_buf ckbuf_in_dp ( .clk(clk), .rclk(rclk), .enb_l(1'b0), .tmb_l(se_l)
         );
  dff_SIZE5 i_fp_id_in ( .din(fpio_data_px2_116_112), .clk(clk), .q(fp_id_in), 
        .se(se), .si({net16637, net16638, net16639, net16640, net16641}) );
  dff_SIZE8 i_fp_op_in ( .din(fpio_data_px2_79_72), .clk(clk), .q(fp_op_in), 
        .se(se), .si({net16629, net16630, net16631, net16632, net16633, 
        net16634, net16635, net16636}) );
  dff_SIZE2 i_fp_fcc_in ( .din(fpio_data_px2_67_0[67:66]), .clk(clk), .q(
        fp_fcc_in), .se(se), .si({net16627, net16628}) );
  dff_SIZE2 i_fp_rnd_mode_in ( .din(fpio_data_px2_67_0[65:64]), .clk(clk), .q(
        fp_rnd_mode_in), .se(se), .si({net16625, net16626}) );
  dff_SIZE64 i_fp_srca_in ( .din(fpio_data_px2_67_0[63:0]), .clk(clk), .q(
        fp_srca_in), .se(se), .si({net16561, net16562, net16563, net16564, 
        net16565, net16566, net16567, net16568, net16569, net16570, net16571, 
        net16572, net16573, net16574, net16575, net16576, net16577, net16578, 
        net16579, net16580, net16581, net16582, net16583, net16584, net16585, 
        net16586, net16587, net16588, net16589, net16590, net16591, net16592, 
        net16593, net16594, net16595, net16596, net16597, net16598, net16599, 
        net16600, net16601, net16602, net16603, net16604, net16605, net16606, 
        net16607, net16608, net16609, net16610, net16611, net16612, net16613, 
        net16614, net16615, net16616, net16617, net16618, net16619, net16620, 
        net16621, net16622, net16623, net16624}) );
  dffe_SIZE69 i_fp_srcb_in ( .din({fp_srca_exp_neq_ffs, fp_srca_exp_eq_0, 
        fp_srca_53_0_neq_0, fp_srca_50_0_neq_0, fp_srca_53_32_neq_0, 
        fp_srca_in}), .en(fp_data_rdy), .clk(clk), .q(fp_srcb_in), .se(se), 
        .si({net16492, net16493, net16494, net16495, net16496, net16497, 
        net16498, net16499, net16500, net16501, net16502, net16503, net16504, 
        net16505, net16506, net16507, net16508, net16509, net16510, net16511, 
        net16512, net16513, net16514, net16515, net16516, net16517, net16518, 
        net16519, net16520, net16521, net16522, net16523, net16524, net16525, 
        net16526, net16527, net16528, net16529, net16530, net16531, net16532, 
        net16533, net16534, net16535, net16536, net16537, net16538, net16539, 
        net16540, net16541, net16542, net16543, net16544, net16545, net16546, 
        net16547, net16548, net16549, net16550, net16551, net16552, net16553, 
        net16554, net16555, net16556, net16557, net16558, net16559, net16560})
         );
  dff_SIZE155 i_inq_din_d1 ( .din({fp_id_in, fp_rnd_mode_in, fp_fcc_in, 
        fp_op_in, fp_src1_in, fp_src2_in}), .clk(clk), .q(inq_din_d1), .se(se), 
        .si({net16337, net16338, net16339, net16340, net16341, net16342, 
        net16343, net16344, net16345, net16346, net16347, net16348, net16349, 
        net16350, net16351, net16352, net16353, net16354, net16355, net16356, 
        net16357, net16358, net16359, net16360, net16361, net16362, net16363, 
        net16364, net16365, net16366, net16367, net16368, net16369, net16370, 
        net16371, net16372, net16373, net16374, net16375, net16376, net16377, 
        net16378, net16379, net16380, net16381, net16382, net16383, net16384, 
        net16385, net16386, net16387, net16388, net16389, net16390, net16391, 
        net16392, net16393, net16394, net16395, net16396, net16397, net16398, 
        net16399, net16400, net16401, net16402, net16403, net16404, net16405, 
        net16406, net16407, net16408, net16409, net16410, net16411, net16412, 
        net16413, net16414, net16415, net16416, net16417, net16418, net16419, 
        net16420, net16421, net16422, net16423, net16424, net16425, net16426, 
        net16427, net16428, net16429, net16430, net16431, net16432, net16433, 
        net16434, net16435, net16436, net16437, net16438, net16439, net16440, 
        net16441, net16442, net16443, net16444, net16445, net16446, net16447, 
        net16448, net16449, net16450, net16451, net16452, net16453, net16454, 
        net16455, net16456, net16457, net16458, net16459, net16460, net16461, 
        net16462, net16463, net16464, net16465, net16466, net16467, net16468, 
        net16469, net16470, net16471, net16472, net16473, net16474, net16475, 
        net16476, net16477, net16478, net16479, net16480, net16481, net16482, 
        net16483, net16484, net16485, net16486, net16487, net16488, net16489, 
        net16490, net16491}) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_NOT I_1 ( .A(fp_op_in[7]), .Z(fp_op_in_7_inv) );
  GTECH_OR2 C309 ( .A(N51), .B(fp_srca_in[0]), .Z(fp_srca_53_0_neq_0) );
  GTECH_OR2 C310 ( .A(N50), .B(fp_srca_in[1]), .Z(N51) );
  GTECH_OR2 C311 ( .A(N49), .B(fp_srca_in[2]), .Z(N50) );
  GTECH_OR2 C312 ( .A(N48), .B(fp_srca_in[3]), .Z(N49) );
  GTECH_OR2 C313 ( .A(N47), .B(fp_srca_in[4]), .Z(N48) );
  GTECH_OR2 C314 ( .A(N46), .B(fp_srca_in[5]), .Z(N47) );
  GTECH_OR2 C315 ( .A(N45), .B(fp_srca_in[6]), .Z(N46) );
  GTECH_OR2 C316 ( .A(N44), .B(fp_srca_in[7]), .Z(N45) );
  GTECH_OR2 C317 ( .A(N43), .B(fp_srca_in[8]), .Z(N44) );
  GTECH_OR2 C318 ( .A(N42), .B(fp_srca_in[9]), .Z(N43) );
  GTECH_OR2 C319 ( .A(N41), .B(fp_srca_in[10]), .Z(N42) );
  GTECH_OR2 C320 ( .A(N40), .B(fp_srca_in[11]), .Z(N41) );
  GTECH_OR2 C321 ( .A(N39), .B(fp_srca_in[12]), .Z(N40) );
  GTECH_OR2 C322 ( .A(N38), .B(fp_srca_in[13]), .Z(N39) );
  GTECH_OR2 C323 ( .A(N37), .B(fp_srca_in[14]), .Z(N38) );
  GTECH_OR2 C324 ( .A(N36), .B(fp_srca_in[15]), .Z(N37) );
  GTECH_OR2 C325 ( .A(N35), .B(fp_srca_in[16]), .Z(N36) );
  GTECH_OR2 C326 ( .A(N34), .B(fp_srca_in[17]), .Z(N35) );
  GTECH_OR2 C327 ( .A(N33), .B(fp_srca_in[18]), .Z(N34) );
  GTECH_OR2 C328 ( .A(N32), .B(fp_srca_in[19]), .Z(N33) );
  GTECH_OR2 C329 ( .A(N31), .B(fp_srca_in[20]), .Z(N32) );
  GTECH_OR2 C330 ( .A(N30), .B(fp_srca_in[21]), .Z(N31) );
  GTECH_OR2 C331 ( .A(N29), .B(fp_srca_in[22]), .Z(N30) );
  GTECH_OR2 C332 ( .A(N28), .B(fp_srca_in[23]), .Z(N29) );
  GTECH_OR2 C333 ( .A(N27), .B(fp_srca_in[24]), .Z(N28) );
  GTECH_OR2 C334 ( .A(N26), .B(fp_srca_in[25]), .Z(N27) );
  GTECH_OR2 C335 ( .A(N25), .B(fp_srca_in[26]), .Z(N26) );
  GTECH_OR2 C336 ( .A(N24), .B(fp_srca_in[27]), .Z(N25) );
  GTECH_OR2 C337 ( .A(N23), .B(fp_srca_in[28]), .Z(N24) );
  GTECH_OR2 C338 ( .A(N22), .B(fp_srca_in[29]), .Z(N23) );
  GTECH_OR2 C339 ( .A(N21), .B(fp_srca_in[30]), .Z(N22) );
  GTECH_OR2 C340 ( .A(N20), .B(fp_srca_in[31]), .Z(N21) );
  GTECH_OR2 C341 ( .A(N19), .B(fp_srca_in[32]), .Z(N20) );
  GTECH_OR2 C342 ( .A(N18), .B(fp_srca_in[33]), .Z(N19) );
  GTECH_OR2 C343 ( .A(N17), .B(fp_srca_in[34]), .Z(N18) );
  GTECH_OR2 C344 ( .A(N16), .B(fp_srca_in[35]), .Z(N17) );
  GTECH_OR2 C345 ( .A(N15), .B(fp_srca_in[36]), .Z(N16) );
  GTECH_OR2 C346 ( .A(N14), .B(fp_srca_in[37]), .Z(N15) );
  GTECH_OR2 C347 ( .A(N13), .B(fp_srca_in[38]), .Z(N14) );
  GTECH_OR2 C348 ( .A(N12), .B(fp_srca_in[39]), .Z(N13) );
  GTECH_OR2 C349 ( .A(N11), .B(fp_srca_in[40]), .Z(N12) );
  GTECH_OR2 C350 ( .A(N10), .B(fp_srca_in[41]), .Z(N11) );
  GTECH_OR2 C351 ( .A(N9), .B(fp_srca_in[42]), .Z(N10) );
  GTECH_OR2 C352 ( .A(N8), .B(fp_srca_in[43]), .Z(N9) );
  GTECH_OR2 C353 ( .A(N7), .B(fp_srca_in[44]), .Z(N8) );
  GTECH_OR2 C354 ( .A(N6), .B(fp_srca_in[45]), .Z(N7) );
  GTECH_OR2 C355 ( .A(N5), .B(fp_srca_in[46]), .Z(N6) );
  GTECH_OR2 C356 ( .A(N4), .B(fp_srca_in[47]), .Z(N5) );
  GTECH_OR2 C357 ( .A(N3), .B(fp_srca_in[48]), .Z(N4) );
  GTECH_OR2 C358 ( .A(N2), .B(fp_srca_in[49]), .Z(N3) );
  GTECH_OR2 C359 ( .A(N1), .B(fp_srca_in[50]), .Z(N2) );
  GTECH_OR2 C360 ( .A(N0), .B(fp_srca_in[51]), .Z(N1) );
  GTECH_OR2 C361 ( .A(fp_srca_in[53]), .B(fp_srca_in[52]), .Z(N0) );
  GTECH_OR2 C362 ( .A(N100), .B(fp_srca_in[0]), .Z(fp_srca_50_0_neq_0) );
  GTECH_OR2 C363 ( .A(N99), .B(fp_srca_in[1]), .Z(N100) );
  GTECH_OR2 C364 ( .A(N98), .B(fp_srca_in[2]), .Z(N99) );
  GTECH_OR2 C365 ( .A(N97), .B(fp_srca_in[3]), .Z(N98) );
  GTECH_OR2 C366 ( .A(N96), .B(fp_srca_in[4]), .Z(N97) );
  GTECH_OR2 C367 ( .A(N95), .B(fp_srca_in[5]), .Z(N96) );
  GTECH_OR2 C368 ( .A(N94), .B(fp_srca_in[6]), .Z(N95) );
  GTECH_OR2 C369 ( .A(N93), .B(fp_srca_in[7]), .Z(N94) );
  GTECH_OR2 C370 ( .A(N92), .B(fp_srca_in[8]), .Z(N93) );
  GTECH_OR2 C371 ( .A(N91), .B(fp_srca_in[9]), .Z(N92) );
  GTECH_OR2 C372 ( .A(N90), .B(fp_srca_in[10]), .Z(N91) );
  GTECH_OR2 C373 ( .A(N89), .B(fp_srca_in[11]), .Z(N90) );
  GTECH_OR2 C374 ( .A(N88), .B(fp_srca_in[12]), .Z(N89) );
  GTECH_OR2 C375 ( .A(N87), .B(fp_srca_in[13]), .Z(N88) );
  GTECH_OR2 C376 ( .A(N86), .B(fp_srca_in[14]), .Z(N87) );
  GTECH_OR2 C377 ( .A(N85), .B(fp_srca_in[15]), .Z(N86) );
  GTECH_OR2 C378 ( .A(N84), .B(fp_srca_in[16]), .Z(N85) );
  GTECH_OR2 C379 ( .A(N83), .B(fp_srca_in[17]), .Z(N84) );
  GTECH_OR2 C380 ( .A(N82), .B(fp_srca_in[18]), .Z(N83) );
  GTECH_OR2 C381 ( .A(N81), .B(fp_srca_in[19]), .Z(N82) );
  GTECH_OR2 C382 ( .A(N80), .B(fp_srca_in[20]), .Z(N81) );
  GTECH_OR2 C383 ( .A(N79), .B(fp_srca_in[21]), .Z(N80) );
  GTECH_OR2 C384 ( .A(N78), .B(fp_srca_in[22]), .Z(N79) );
  GTECH_OR2 C385 ( .A(N77), .B(fp_srca_in[23]), .Z(N78) );
  GTECH_OR2 C386 ( .A(N76), .B(fp_srca_in[24]), .Z(N77) );
  GTECH_OR2 C387 ( .A(N75), .B(fp_srca_in[25]), .Z(N76) );
  GTECH_OR2 C388 ( .A(N74), .B(fp_srca_in[26]), .Z(N75) );
  GTECH_OR2 C389 ( .A(N73), .B(fp_srca_in[27]), .Z(N74) );
  GTECH_OR2 C390 ( .A(N72), .B(fp_srca_in[28]), .Z(N73) );
  GTECH_OR2 C391 ( .A(N71), .B(fp_srca_in[29]), .Z(N72) );
  GTECH_OR2 C392 ( .A(N70), .B(fp_srca_in[30]), .Z(N71) );
  GTECH_OR2 C393 ( .A(N69), .B(fp_srca_in[31]), .Z(N70) );
  GTECH_OR2 C394 ( .A(N68), .B(fp_srca_in[32]), .Z(N69) );
  GTECH_OR2 C395 ( .A(N67), .B(fp_srca_in[33]), .Z(N68) );
  GTECH_OR2 C396 ( .A(N66), .B(fp_srca_in[34]), .Z(N67) );
  GTECH_OR2 C397 ( .A(N65), .B(fp_srca_in[35]), .Z(N66) );
  GTECH_OR2 C398 ( .A(N64), .B(fp_srca_in[36]), .Z(N65) );
  GTECH_OR2 C399 ( .A(N63), .B(fp_srca_in[37]), .Z(N64) );
  GTECH_OR2 C400 ( .A(N62), .B(fp_srca_in[38]), .Z(N63) );
  GTECH_OR2 C401 ( .A(N61), .B(fp_srca_in[39]), .Z(N62) );
  GTECH_OR2 C402 ( .A(N60), .B(fp_srca_in[40]), .Z(N61) );
  GTECH_OR2 C403 ( .A(N59), .B(fp_srca_in[41]), .Z(N60) );
  GTECH_OR2 C404 ( .A(N58), .B(fp_srca_in[42]), .Z(N59) );
  GTECH_OR2 C405 ( .A(N57), .B(fp_srca_in[43]), .Z(N58) );
  GTECH_OR2 C406 ( .A(N56), .B(fp_srca_in[44]), .Z(N57) );
  GTECH_OR2 C407 ( .A(N55), .B(fp_srca_in[45]), .Z(N56) );
  GTECH_OR2 C408 ( .A(N54), .B(fp_srca_in[46]), .Z(N55) );
  GTECH_OR2 C409 ( .A(N53), .B(fp_srca_in[47]), .Z(N54) );
  GTECH_OR2 C410 ( .A(N52), .B(fp_srca_in[48]), .Z(N53) );
  GTECH_OR2 C411 ( .A(fp_srca_in[50]), .B(fp_srca_in[49]), .Z(N52) );
  GTECH_OR2 C412 ( .A(N120), .B(fp_srca_in[32]), .Z(fp_srca_53_32_neq_0) );
  GTECH_OR2 C413 ( .A(N119), .B(fp_srca_in[33]), .Z(N120) );
  GTECH_OR2 C414 ( .A(N118), .B(fp_srca_in[34]), .Z(N119) );
  GTECH_OR2 C415 ( .A(N117), .B(fp_srca_in[35]), .Z(N118) );
  GTECH_OR2 C416 ( .A(N116), .B(fp_srca_in[36]), .Z(N117) );
  GTECH_OR2 C417 ( .A(N115), .B(fp_srca_in[37]), .Z(N116) );
  GTECH_OR2 C418 ( .A(N114), .B(fp_srca_in[38]), .Z(N115) );
  GTECH_OR2 C419 ( .A(N113), .B(fp_srca_in[39]), .Z(N114) );
  GTECH_OR2 C420 ( .A(N112), .B(fp_srca_in[40]), .Z(N113) );
  GTECH_OR2 C421 ( .A(N111), .B(fp_srca_in[41]), .Z(N112) );
  GTECH_OR2 C422 ( .A(N110), .B(fp_srca_in[42]), .Z(N111) );
  GTECH_OR2 C423 ( .A(N109), .B(fp_srca_in[43]), .Z(N110) );
  GTECH_OR2 C424 ( .A(N108), .B(fp_srca_in[44]), .Z(N109) );
  GTECH_OR2 C425 ( .A(N107), .B(fp_srca_in[45]), .Z(N108) );
  GTECH_OR2 C426 ( .A(N106), .B(fp_srca_in[46]), .Z(N107) );
  GTECH_OR2 C427 ( .A(N105), .B(fp_srca_in[47]), .Z(N106) );
  GTECH_OR2 C428 ( .A(N104), .B(fp_srca_in[48]), .Z(N105) );
  GTECH_OR2 C429 ( .A(N103), .B(fp_srca_in[49]), .Z(N104) );
  GTECH_OR2 C430 ( .A(N102), .B(fp_srca_in[50]), .Z(N103) );
  GTECH_OR2 C431 ( .A(N101), .B(fp_srca_in[51]), .Z(N102) );
  GTECH_OR2 C432 ( .A(fp_srca_in[53]), .B(fp_srca_in[52]), .Z(N101) );
  GTECH_NOT I_2 ( .A(N131), .Z(fp_srca_exp_eq_0) );
  GTECH_OR2 C434 ( .A(N127), .B(N130), .Z(N131) );
  GTECH_OR2 C435 ( .A(N126), .B(fp_srca_in[55]), .Z(N127) );
  GTECH_OR2 C436 ( .A(N125), .B(fp_srca_in[56]), .Z(N126) );
  GTECH_OR2 C437 ( .A(N124), .B(fp_srca_in[57]), .Z(N125) );
  GTECH_OR2 C438 ( .A(N123), .B(fp_srca_in[58]), .Z(N124) );
  GTECH_OR2 C439 ( .A(N122), .B(fp_srca_in[59]), .Z(N123) );
  GTECH_OR2 C440 ( .A(N121), .B(fp_srca_in[60]), .Z(N122) );
  GTECH_OR2 C441 ( .A(fp_srca_in[62]), .B(fp_srca_in[61]), .Z(N121) );
  GTECH_AND2 C442 ( .A(fp_op_in[1]), .B(N129), .Z(N130) );
  GTECH_OR2 C443 ( .A(N128), .B(fp_srca_in[52]), .Z(N129) );
  GTECH_OR2 C444 ( .A(fp_srca_in[54]), .B(fp_srca_in[53]), .Z(N128) );
  GTECH_NOT I_3 ( .A(N142), .Z(fp_srca_exp_neq_ffs) );
  GTECH_AND2 C446 ( .A(N138), .B(N141), .Z(N142) );
  GTECH_AND2 C447 ( .A(N137), .B(fp_srca_in[55]), .Z(N138) );
  GTECH_AND2 C448 ( .A(N136), .B(fp_srca_in[56]), .Z(N137) );
  GTECH_AND2 C449 ( .A(N135), .B(fp_srca_in[57]), .Z(N136) );
  GTECH_AND2 C450 ( .A(N134), .B(fp_srca_in[58]), .Z(N135) );
  GTECH_AND2 C451 ( .A(N133), .B(fp_srca_in[59]), .Z(N134) );
  GTECH_AND2 C452 ( .A(N132), .B(fp_srca_in[60]), .Z(N133) );
  GTECH_AND2 C453 ( .A(fp_srca_in[62]), .B(fp_srca_in[61]), .Z(N132) );
  GTECH_OR2 C454 ( .A(fp_op_in[0]), .B(N140), .Z(N141) );
  GTECH_AND2 C455 ( .A(N139), .B(fp_srca_in[52]), .Z(N140) );
  GTECH_AND2 C456 ( .A(fp_srca_in[54]), .B(fp_srca_in[53]), .Z(N139) );
  GTECH_OR2 C457 ( .A(N143), .B(fp_op_in[7]), .Z(fp_src1_in[68]) );
  GTECH_AND2 C458 ( .A(fp_op_in_7_inv), .B(fp_srca_exp_neq_ffs), .Z(N143) );
  GTECH_OR2 C459 ( .A(N144), .B(fp_op_in[7]), .Z(fp_src1_in[67]) );
  GTECH_AND2 C460 ( .A(fp_op_in_7_inv), .B(fp_srca_exp_eq_0), .Z(N144) );
  GTECH_AND2 C461 ( .A(fp_op_in_7_inv), .B(fp_srca_53_0_neq_0), .Z(
        fp_src1_in[66]) );
  GTECH_AND2 C462 ( .A(fp_op_in_7_inv), .B(fp_srca_50_0_neq_0), .Z(
        fp_src1_in[65]) );
  GTECH_AND2 C463 ( .A(fp_op_in_7_inv), .B(fp_srca_53_32_neq_0), .Z(
        fp_src1_in[64]) );
  GTECH_AND2 C464 ( .A(fp_op_in_7_inv), .B(fp_srca_in[63]), .Z(fp_src1_in[63])
         );
  GTECH_AND2 C465 ( .A(fp_op_in_7_inv), .B(fp_srca_in[62]), .Z(fp_src1_in[62])
         );
  GTECH_AND2 C466 ( .A(fp_op_in_7_inv), .B(fp_srca_in[61]), .Z(fp_src1_in[61])
         );
  GTECH_AND2 C467 ( .A(fp_op_in_7_inv), .B(fp_srca_in[60]), .Z(fp_src1_in[60])
         );
  GTECH_AND2 C468 ( .A(fp_op_in_7_inv), .B(fp_srca_in[59]), .Z(fp_src1_in[59])
         );
  GTECH_AND2 C469 ( .A(fp_op_in_7_inv), .B(fp_srca_in[58]), .Z(fp_src1_in[58])
         );
  GTECH_AND2 C470 ( .A(fp_op_in_7_inv), .B(fp_srca_in[57]), .Z(fp_src1_in[57])
         );
  GTECH_AND2 C471 ( .A(fp_op_in_7_inv), .B(fp_srca_in[56]), .Z(fp_src1_in[56])
         );
  GTECH_AND2 C472 ( .A(fp_op_in_7_inv), .B(fp_srca_in[55]), .Z(fp_src1_in[55])
         );
  GTECH_AND2 C473 ( .A(fp_op_in_7_inv), .B(fp_srca_in[54]), .Z(fp_src1_in[54])
         );
  GTECH_AND2 C474 ( .A(fp_op_in_7_inv), .B(fp_srca_in[53]), .Z(fp_src1_in[53])
         );
  GTECH_AND2 C475 ( .A(fp_op_in_7_inv), .B(fp_srca_in[52]), .Z(fp_src1_in[52])
         );
  GTECH_AND2 C476 ( .A(fp_op_in_7_inv), .B(fp_srca_in[51]), .Z(fp_src1_in[51])
         );
  GTECH_AND2 C477 ( .A(fp_op_in_7_inv), .B(fp_srca_in[50]), .Z(fp_src1_in[50])
         );
  GTECH_AND2 C478 ( .A(fp_op_in_7_inv), .B(fp_srca_in[49]), .Z(fp_src1_in[49])
         );
  GTECH_AND2 C479 ( .A(fp_op_in_7_inv), .B(fp_srca_in[48]), .Z(fp_src1_in[48])
         );
  GTECH_AND2 C480 ( .A(fp_op_in_7_inv), .B(fp_srca_in[47]), .Z(fp_src1_in[47])
         );
  GTECH_AND2 C481 ( .A(fp_op_in_7_inv), .B(fp_srca_in[46]), .Z(fp_src1_in[46])
         );
  GTECH_AND2 C482 ( .A(fp_op_in_7_inv), .B(fp_srca_in[45]), .Z(fp_src1_in[45])
         );
  GTECH_AND2 C483 ( .A(fp_op_in_7_inv), .B(fp_srca_in[44]), .Z(fp_src1_in[44])
         );
  GTECH_AND2 C484 ( .A(fp_op_in_7_inv), .B(fp_srca_in[43]), .Z(fp_src1_in[43])
         );
  GTECH_AND2 C485 ( .A(fp_op_in_7_inv), .B(fp_srca_in[42]), .Z(fp_src1_in[42])
         );
  GTECH_AND2 C486 ( .A(fp_op_in_7_inv), .B(fp_srca_in[41]), .Z(fp_src1_in[41])
         );
  GTECH_AND2 C487 ( .A(fp_op_in_7_inv), .B(fp_srca_in[40]), .Z(fp_src1_in[40])
         );
  GTECH_AND2 C488 ( .A(fp_op_in_7_inv), .B(fp_srca_in[39]), .Z(fp_src1_in[39])
         );
  GTECH_AND2 C489 ( .A(fp_op_in_7_inv), .B(fp_srca_in[38]), .Z(fp_src1_in[38])
         );
  GTECH_AND2 C490 ( .A(fp_op_in_7_inv), .B(fp_srca_in[37]), .Z(fp_src1_in[37])
         );
  GTECH_AND2 C491 ( .A(fp_op_in_7_inv), .B(fp_srca_in[36]), .Z(fp_src1_in[36])
         );
  GTECH_AND2 C492 ( .A(fp_op_in_7_inv), .B(fp_srca_in[35]), .Z(fp_src1_in[35])
         );
  GTECH_AND2 C493 ( .A(fp_op_in_7_inv), .B(fp_srca_in[34]), .Z(fp_src1_in[34])
         );
  GTECH_AND2 C494 ( .A(fp_op_in_7_inv), .B(fp_srca_in[33]), .Z(fp_src1_in[33])
         );
  GTECH_AND2 C495 ( .A(fp_op_in_7_inv), .B(fp_srca_in[32]), .Z(fp_src1_in[32])
         );
  GTECH_AND2 C496 ( .A(fp_op_in_7_inv), .B(fp_srca_in[31]), .Z(fp_src1_in[31])
         );
  GTECH_AND2 C497 ( .A(fp_op_in_7_inv), .B(fp_srca_in[30]), .Z(fp_src1_in[30])
         );
  GTECH_AND2 C498 ( .A(fp_op_in_7_inv), .B(fp_srca_in[29]), .Z(fp_src1_in[29])
         );
  GTECH_AND2 C499 ( .A(fp_op_in_7_inv), .B(fp_srca_in[28]), .Z(fp_src1_in[28])
         );
  GTECH_AND2 C500 ( .A(fp_op_in_7_inv), .B(fp_srca_in[27]), .Z(fp_src1_in[27])
         );
  GTECH_AND2 C501 ( .A(fp_op_in_7_inv), .B(fp_srca_in[26]), .Z(fp_src1_in[26])
         );
  GTECH_AND2 C502 ( .A(fp_op_in_7_inv), .B(fp_srca_in[25]), .Z(fp_src1_in[25])
         );
  GTECH_AND2 C503 ( .A(fp_op_in_7_inv), .B(fp_srca_in[24]), .Z(fp_src1_in[24])
         );
  GTECH_AND2 C504 ( .A(fp_op_in_7_inv), .B(fp_srca_in[23]), .Z(fp_src1_in[23])
         );
  GTECH_AND2 C505 ( .A(fp_op_in_7_inv), .B(fp_srca_in[22]), .Z(fp_src1_in[22])
         );
  GTECH_AND2 C506 ( .A(fp_op_in_7_inv), .B(fp_srca_in[21]), .Z(fp_src1_in[21])
         );
  GTECH_AND2 C507 ( .A(fp_op_in_7_inv), .B(fp_srca_in[20]), .Z(fp_src1_in[20])
         );
  GTECH_AND2 C508 ( .A(fp_op_in_7_inv), .B(fp_srca_in[19]), .Z(fp_src1_in[19])
         );
  GTECH_AND2 C509 ( .A(fp_op_in_7_inv), .B(fp_srca_in[18]), .Z(fp_src1_in[18])
         );
  GTECH_AND2 C510 ( .A(fp_op_in_7_inv), .B(fp_srca_in[17]), .Z(fp_src1_in[17])
         );
  GTECH_AND2 C511 ( .A(fp_op_in_7_inv), .B(fp_srca_in[16]), .Z(fp_src1_in[16])
         );
  GTECH_AND2 C512 ( .A(fp_op_in_7_inv), .B(fp_srca_in[15]), .Z(fp_src1_in[15])
         );
  GTECH_AND2 C513 ( .A(fp_op_in_7_inv), .B(fp_srca_in[14]), .Z(fp_src1_in[14])
         );
  GTECH_AND2 C514 ( .A(fp_op_in_7_inv), .B(fp_srca_in[13]), .Z(fp_src1_in[13])
         );
  GTECH_AND2 C515 ( .A(fp_op_in_7_inv), .B(fp_srca_in[12]), .Z(fp_src1_in[12])
         );
  GTECH_AND2 C516 ( .A(fp_op_in_7_inv), .B(fp_srca_in[11]), .Z(fp_src1_in[11])
         );
  GTECH_AND2 C517 ( .A(fp_op_in_7_inv), .B(fp_srca_in[10]), .Z(fp_src1_in[10])
         );
  GTECH_AND2 C518 ( .A(fp_op_in_7_inv), .B(fp_srca_in[9]), .Z(fp_src1_in[9])
         );
  GTECH_AND2 C519 ( .A(fp_op_in_7_inv), .B(fp_srca_in[8]), .Z(fp_src1_in[8])
         );
  GTECH_AND2 C520 ( .A(fp_op_in_7_inv), .B(fp_srca_in[7]), .Z(fp_src1_in[7])
         );
  GTECH_AND2 C521 ( .A(fp_op_in_7_inv), .B(fp_srca_in[6]), .Z(fp_src1_in[6])
         );
  GTECH_AND2 C522 ( .A(fp_op_in_7_inv), .B(fp_srca_in[5]), .Z(fp_src1_in[5])
         );
  GTECH_AND2 C523 ( .A(fp_op_in_7_inv), .B(fp_srca_in[4]), .Z(fp_src1_in[4])
         );
  GTECH_AND2 C524 ( .A(fp_op_in_7_inv), .B(fp_srca_in[3]), .Z(fp_src1_in[3])
         );
  GTECH_AND2 C525 ( .A(fp_op_in_7_inv), .B(fp_srca_in[2]), .Z(fp_src1_in[2])
         );
  GTECH_AND2 C526 ( .A(fp_op_in_7_inv), .B(fp_srca_in[1]), .Z(fp_src1_in[1])
         );
  GTECH_AND2 C527 ( .A(fp_op_in_7_inv), .B(fp_srca_in[0]), .Z(fp_src1_in[0])
         );
  GTECH_OR2 C528 ( .A(N145), .B(N146), .Z(fp_src2_in[68]) );
  GTECH_AND2 C529 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[68]), .Z(N145) );
  GTECH_AND2 C530 ( .A(fp_op_in[7]), .B(fp_srca_exp_neq_ffs), .Z(N146) );
  GTECH_OR2 C531 ( .A(N147), .B(N148), .Z(fp_src2_in[67]) );
  GTECH_AND2 C532 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[67]), .Z(N147) );
  GTECH_AND2 C533 ( .A(fp_op_in[7]), .B(fp_srca_exp_eq_0), .Z(N148) );
  GTECH_OR2 C534 ( .A(N149), .B(N150), .Z(fp_src2_in[66]) );
  GTECH_AND2 C535 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[66]), .Z(N149) );
  GTECH_AND2 C536 ( .A(fp_op_in[7]), .B(fp_srca_53_0_neq_0), .Z(N150) );
  GTECH_OR2 C537 ( .A(N151), .B(N152), .Z(fp_src2_in[65]) );
  GTECH_AND2 C538 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[65]), .Z(N151) );
  GTECH_AND2 C539 ( .A(fp_op_in[7]), .B(fp_srca_50_0_neq_0), .Z(N152) );
  GTECH_OR2 C540 ( .A(N153), .B(N154), .Z(fp_src2_in[64]) );
  GTECH_AND2 C541 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[64]), .Z(N153) );
  GTECH_AND2 C542 ( .A(fp_op_in[7]), .B(fp_srca_53_32_neq_0), .Z(N154) );
  GTECH_OR2 C543 ( .A(N155), .B(N156), .Z(fp_src2_in[63]) );
  GTECH_AND2 C544 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[63]), .Z(N155) );
  GTECH_AND2 C545 ( .A(fp_op_in[7]), .B(fp_srca_in[63]), .Z(N156) );
  GTECH_OR2 C546 ( .A(N157), .B(N158), .Z(fp_src2_in[62]) );
  GTECH_AND2 C547 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[62]), .Z(N157) );
  GTECH_AND2 C548 ( .A(fp_op_in[7]), .B(fp_srca_in[62]), .Z(N158) );
  GTECH_OR2 C549 ( .A(N159), .B(N160), .Z(fp_src2_in[61]) );
  GTECH_AND2 C550 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[61]), .Z(N159) );
  GTECH_AND2 C551 ( .A(fp_op_in[7]), .B(fp_srca_in[61]), .Z(N160) );
  GTECH_OR2 C552 ( .A(N161), .B(N162), .Z(fp_src2_in[60]) );
  GTECH_AND2 C553 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[60]), .Z(N161) );
  GTECH_AND2 C554 ( .A(fp_op_in[7]), .B(fp_srca_in[60]), .Z(N162) );
  GTECH_OR2 C555 ( .A(N163), .B(N164), .Z(fp_src2_in[59]) );
  GTECH_AND2 C556 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[59]), .Z(N163) );
  GTECH_AND2 C557 ( .A(fp_op_in[7]), .B(fp_srca_in[59]), .Z(N164) );
  GTECH_OR2 C558 ( .A(N165), .B(N166), .Z(fp_src2_in[58]) );
  GTECH_AND2 C559 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[58]), .Z(N165) );
  GTECH_AND2 C560 ( .A(fp_op_in[7]), .B(fp_srca_in[58]), .Z(N166) );
  GTECH_OR2 C561 ( .A(N167), .B(N168), .Z(fp_src2_in[57]) );
  GTECH_AND2 C562 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[57]), .Z(N167) );
  GTECH_AND2 C563 ( .A(fp_op_in[7]), .B(fp_srca_in[57]), .Z(N168) );
  GTECH_OR2 C564 ( .A(N169), .B(N170), .Z(fp_src2_in[56]) );
  GTECH_AND2 C565 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[56]), .Z(N169) );
  GTECH_AND2 C566 ( .A(fp_op_in[7]), .B(fp_srca_in[56]), .Z(N170) );
  GTECH_OR2 C567 ( .A(N171), .B(N172), .Z(fp_src2_in[55]) );
  GTECH_AND2 C568 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[55]), .Z(N171) );
  GTECH_AND2 C569 ( .A(fp_op_in[7]), .B(fp_srca_in[55]), .Z(N172) );
  GTECH_OR2 C570 ( .A(N173), .B(N174), .Z(fp_src2_in[54]) );
  GTECH_AND2 C571 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[54]), .Z(N173) );
  GTECH_AND2 C572 ( .A(fp_op_in[7]), .B(fp_srca_in[54]), .Z(N174) );
  GTECH_OR2 C573 ( .A(N175), .B(N176), .Z(fp_src2_in[53]) );
  GTECH_AND2 C574 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[53]), .Z(N175) );
  GTECH_AND2 C575 ( .A(fp_op_in[7]), .B(fp_srca_in[53]), .Z(N176) );
  GTECH_OR2 C576 ( .A(N177), .B(N178), .Z(fp_src2_in[52]) );
  GTECH_AND2 C577 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[52]), .Z(N177) );
  GTECH_AND2 C578 ( .A(fp_op_in[7]), .B(fp_srca_in[52]), .Z(N178) );
  GTECH_OR2 C579 ( .A(N179), .B(N180), .Z(fp_src2_in[51]) );
  GTECH_AND2 C580 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[51]), .Z(N179) );
  GTECH_AND2 C581 ( .A(fp_op_in[7]), .B(fp_srca_in[51]), .Z(N180) );
  GTECH_OR2 C582 ( .A(N181), .B(N182), .Z(fp_src2_in[50]) );
  GTECH_AND2 C583 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[50]), .Z(N181) );
  GTECH_AND2 C584 ( .A(fp_op_in[7]), .B(fp_srca_in[50]), .Z(N182) );
  GTECH_OR2 C585 ( .A(N183), .B(N184), .Z(fp_src2_in[49]) );
  GTECH_AND2 C586 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[49]), .Z(N183) );
  GTECH_AND2 C587 ( .A(fp_op_in[7]), .B(fp_srca_in[49]), .Z(N184) );
  GTECH_OR2 C588 ( .A(N185), .B(N186), .Z(fp_src2_in[48]) );
  GTECH_AND2 C589 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[48]), .Z(N185) );
  GTECH_AND2 C590 ( .A(fp_op_in[7]), .B(fp_srca_in[48]), .Z(N186) );
  GTECH_OR2 C591 ( .A(N187), .B(N188), .Z(fp_src2_in[47]) );
  GTECH_AND2 C592 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[47]), .Z(N187) );
  GTECH_AND2 C593 ( .A(fp_op_in[7]), .B(fp_srca_in[47]), .Z(N188) );
  GTECH_OR2 C594 ( .A(N189), .B(N190), .Z(fp_src2_in[46]) );
  GTECH_AND2 C595 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[46]), .Z(N189) );
  GTECH_AND2 C596 ( .A(fp_op_in[7]), .B(fp_srca_in[46]), .Z(N190) );
  GTECH_OR2 C597 ( .A(N191), .B(N192), .Z(fp_src2_in[45]) );
  GTECH_AND2 C598 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[45]), .Z(N191) );
  GTECH_AND2 C599 ( .A(fp_op_in[7]), .B(fp_srca_in[45]), .Z(N192) );
  GTECH_OR2 C600 ( .A(N193), .B(N194), .Z(fp_src2_in[44]) );
  GTECH_AND2 C601 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[44]), .Z(N193) );
  GTECH_AND2 C602 ( .A(fp_op_in[7]), .B(fp_srca_in[44]), .Z(N194) );
  GTECH_OR2 C603 ( .A(N195), .B(N196), .Z(fp_src2_in[43]) );
  GTECH_AND2 C604 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[43]), .Z(N195) );
  GTECH_AND2 C605 ( .A(fp_op_in[7]), .B(fp_srca_in[43]), .Z(N196) );
  GTECH_OR2 C606 ( .A(N197), .B(N198), .Z(fp_src2_in[42]) );
  GTECH_AND2 C607 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[42]), .Z(N197) );
  GTECH_AND2 C608 ( .A(fp_op_in[7]), .B(fp_srca_in[42]), .Z(N198) );
  GTECH_OR2 C609 ( .A(N199), .B(N200), .Z(fp_src2_in[41]) );
  GTECH_AND2 C610 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[41]), .Z(N199) );
  GTECH_AND2 C611 ( .A(fp_op_in[7]), .B(fp_srca_in[41]), .Z(N200) );
  GTECH_OR2 C612 ( .A(N201), .B(N202), .Z(fp_src2_in[40]) );
  GTECH_AND2 C613 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[40]), .Z(N201) );
  GTECH_AND2 C614 ( .A(fp_op_in[7]), .B(fp_srca_in[40]), .Z(N202) );
  GTECH_OR2 C615 ( .A(N203), .B(N204), .Z(fp_src2_in[39]) );
  GTECH_AND2 C616 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[39]), .Z(N203) );
  GTECH_AND2 C617 ( .A(fp_op_in[7]), .B(fp_srca_in[39]), .Z(N204) );
  GTECH_OR2 C618 ( .A(N205), .B(N206), .Z(fp_src2_in[38]) );
  GTECH_AND2 C619 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[38]), .Z(N205) );
  GTECH_AND2 C620 ( .A(fp_op_in[7]), .B(fp_srca_in[38]), .Z(N206) );
  GTECH_OR2 C621 ( .A(N207), .B(N208), .Z(fp_src2_in[37]) );
  GTECH_AND2 C622 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[37]), .Z(N207) );
  GTECH_AND2 C623 ( .A(fp_op_in[7]), .B(fp_srca_in[37]), .Z(N208) );
  GTECH_OR2 C624 ( .A(N209), .B(N210), .Z(fp_src2_in[36]) );
  GTECH_AND2 C625 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[36]), .Z(N209) );
  GTECH_AND2 C626 ( .A(fp_op_in[7]), .B(fp_srca_in[36]), .Z(N210) );
  GTECH_OR2 C627 ( .A(N211), .B(N212), .Z(fp_src2_in[35]) );
  GTECH_AND2 C628 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[35]), .Z(N211) );
  GTECH_AND2 C629 ( .A(fp_op_in[7]), .B(fp_srca_in[35]), .Z(N212) );
  GTECH_OR2 C630 ( .A(N213), .B(N214), .Z(fp_src2_in[34]) );
  GTECH_AND2 C631 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[34]), .Z(N213) );
  GTECH_AND2 C632 ( .A(fp_op_in[7]), .B(fp_srca_in[34]), .Z(N214) );
  GTECH_OR2 C633 ( .A(N215), .B(N216), .Z(fp_src2_in[33]) );
  GTECH_AND2 C634 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[33]), .Z(N215) );
  GTECH_AND2 C635 ( .A(fp_op_in[7]), .B(fp_srca_in[33]), .Z(N216) );
  GTECH_OR2 C636 ( .A(N217), .B(N218), .Z(fp_src2_in[32]) );
  GTECH_AND2 C637 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[32]), .Z(N217) );
  GTECH_AND2 C638 ( .A(fp_op_in[7]), .B(fp_srca_in[32]), .Z(N218) );
  GTECH_OR2 C639 ( .A(N219), .B(N220), .Z(fp_src2_in[31]) );
  GTECH_AND2 C640 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[31]), .Z(N219) );
  GTECH_AND2 C641 ( .A(fp_op_in[7]), .B(fp_srca_in[31]), .Z(N220) );
  GTECH_OR2 C642 ( .A(N221), .B(N222), .Z(fp_src2_in[30]) );
  GTECH_AND2 C643 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[30]), .Z(N221) );
  GTECH_AND2 C644 ( .A(fp_op_in[7]), .B(fp_srca_in[30]), .Z(N222) );
  GTECH_OR2 C645 ( .A(N223), .B(N224), .Z(fp_src2_in[29]) );
  GTECH_AND2 C646 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[29]), .Z(N223) );
  GTECH_AND2 C647 ( .A(fp_op_in[7]), .B(fp_srca_in[29]), .Z(N224) );
  GTECH_OR2 C648 ( .A(N225), .B(N226), .Z(fp_src2_in[28]) );
  GTECH_AND2 C649 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[28]), .Z(N225) );
  GTECH_AND2 C650 ( .A(fp_op_in[7]), .B(fp_srca_in[28]), .Z(N226) );
  GTECH_OR2 C651 ( .A(N227), .B(N228), .Z(fp_src2_in[27]) );
  GTECH_AND2 C652 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[27]), .Z(N227) );
  GTECH_AND2 C653 ( .A(fp_op_in[7]), .B(fp_srca_in[27]), .Z(N228) );
  GTECH_OR2 C654 ( .A(N229), .B(N230), .Z(fp_src2_in[26]) );
  GTECH_AND2 C655 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[26]), .Z(N229) );
  GTECH_AND2 C656 ( .A(fp_op_in[7]), .B(fp_srca_in[26]), .Z(N230) );
  GTECH_OR2 C657 ( .A(N231), .B(N232), .Z(fp_src2_in[25]) );
  GTECH_AND2 C658 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[25]), .Z(N231) );
  GTECH_AND2 C659 ( .A(fp_op_in[7]), .B(fp_srca_in[25]), .Z(N232) );
  GTECH_OR2 C660 ( .A(N233), .B(N234), .Z(fp_src2_in[24]) );
  GTECH_AND2 C661 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[24]), .Z(N233) );
  GTECH_AND2 C662 ( .A(fp_op_in[7]), .B(fp_srca_in[24]), .Z(N234) );
  GTECH_OR2 C663 ( .A(N235), .B(N236), .Z(fp_src2_in[23]) );
  GTECH_AND2 C664 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[23]), .Z(N235) );
  GTECH_AND2 C665 ( .A(fp_op_in[7]), .B(fp_srca_in[23]), .Z(N236) );
  GTECH_OR2 C666 ( .A(N237), .B(N238), .Z(fp_src2_in[22]) );
  GTECH_AND2 C667 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[22]), .Z(N237) );
  GTECH_AND2 C668 ( .A(fp_op_in[7]), .B(fp_srca_in[22]), .Z(N238) );
  GTECH_OR2 C669 ( .A(N239), .B(N240), .Z(fp_src2_in[21]) );
  GTECH_AND2 C670 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[21]), .Z(N239) );
  GTECH_AND2 C671 ( .A(fp_op_in[7]), .B(fp_srca_in[21]), .Z(N240) );
  GTECH_OR2 C672 ( .A(N241), .B(N242), .Z(fp_src2_in[20]) );
  GTECH_AND2 C673 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[20]), .Z(N241) );
  GTECH_AND2 C674 ( .A(fp_op_in[7]), .B(fp_srca_in[20]), .Z(N242) );
  GTECH_OR2 C675 ( .A(N243), .B(N244), .Z(fp_src2_in[19]) );
  GTECH_AND2 C676 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[19]), .Z(N243) );
  GTECH_AND2 C677 ( .A(fp_op_in[7]), .B(fp_srca_in[19]), .Z(N244) );
  GTECH_OR2 C678 ( .A(N245), .B(N246), .Z(fp_src2_in[18]) );
  GTECH_AND2 C679 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[18]), .Z(N245) );
  GTECH_AND2 C680 ( .A(fp_op_in[7]), .B(fp_srca_in[18]), .Z(N246) );
  GTECH_OR2 C681 ( .A(N247), .B(N248), .Z(fp_src2_in[17]) );
  GTECH_AND2 C682 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[17]), .Z(N247) );
  GTECH_AND2 C683 ( .A(fp_op_in[7]), .B(fp_srca_in[17]), .Z(N248) );
  GTECH_OR2 C684 ( .A(N249), .B(N250), .Z(fp_src2_in[16]) );
  GTECH_AND2 C685 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[16]), .Z(N249) );
  GTECH_AND2 C686 ( .A(fp_op_in[7]), .B(fp_srca_in[16]), .Z(N250) );
  GTECH_OR2 C687 ( .A(N251), .B(N252), .Z(fp_src2_in[15]) );
  GTECH_AND2 C688 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[15]), .Z(N251) );
  GTECH_AND2 C689 ( .A(fp_op_in[7]), .B(fp_srca_in[15]), .Z(N252) );
  GTECH_OR2 C690 ( .A(N253), .B(N254), .Z(fp_src2_in[14]) );
  GTECH_AND2 C691 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[14]), .Z(N253) );
  GTECH_AND2 C692 ( .A(fp_op_in[7]), .B(fp_srca_in[14]), .Z(N254) );
  GTECH_OR2 C693 ( .A(N255), .B(N256), .Z(fp_src2_in[13]) );
  GTECH_AND2 C694 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[13]), .Z(N255) );
  GTECH_AND2 C695 ( .A(fp_op_in[7]), .B(fp_srca_in[13]), .Z(N256) );
  GTECH_OR2 C696 ( .A(N257), .B(N258), .Z(fp_src2_in[12]) );
  GTECH_AND2 C697 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[12]), .Z(N257) );
  GTECH_AND2 C698 ( .A(fp_op_in[7]), .B(fp_srca_in[12]), .Z(N258) );
  GTECH_OR2 C699 ( .A(N259), .B(N260), .Z(fp_src2_in[11]) );
  GTECH_AND2 C700 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[11]), .Z(N259) );
  GTECH_AND2 C701 ( .A(fp_op_in[7]), .B(fp_srca_in[11]), .Z(N260) );
  GTECH_OR2 C702 ( .A(N261), .B(N262), .Z(fp_src2_in[10]) );
  GTECH_AND2 C703 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[10]), .Z(N261) );
  GTECH_AND2 C704 ( .A(fp_op_in[7]), .B(fp_srca_in[10]), .Z(N262) );
  GTECH_OR2 C705 ( .A(N263), .B(N264), .Z(fp_src2_in[9]) );
  GTECH_AND2 C706 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[9]), .Z(N263) );
  GTECH_AND2 C707 ( .A(fp_op_in[7]), .B(fp_srca_in[9]), .Z(N264) );
  GTECH_OR2 C708 ( .A(N265), .B(N266), .Z(fp_src2_in[8]) );
  GTECH_AND2 C709 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[8]), .Z(N265) );
  GTECH_AND2 C710 ( .A(fp_op_in[7]), .B(fp_srca_in[8]), .Z(N266) );
  GTECH_OR2 C711 ( .A(N267), .B(N268), .Z(fp_src2_in[7]) );
  GTECH_AND2 C712 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[7]), .Z(N267) );
  GTECH_AND2 C713 ( .A(fp_op_in[7]), .B(fp_srca_in[7]), .Z(N268) );
  GTECH_OR2 C714 ( .A(N269), .B(N270), .Z(fp_src2_in[6]) );
  GTECH_AND2 C715 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[6]), .Z(N269) );
  GTECH_AND2 C716 ( .A(fp_op_in[7]), .B(fp_srca_in[6]), .Z(N270) );
  GTECH_OR2 C717 ( .A(N271), .B(N272), .Z(fp_src2_in[5]) );
  GTECH_AND2 C718 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[5]), .Z(N271) );
  GTECH_AND2 C719 ( .A(fp_op_in[7]), .B(fp_srca_in[5]), .Z(N272) );
  GTECH_OR2 C720 ( .A(N273), .B(N274), .Z(fp_src2_in[4]) );
  GTECH_AND2 C721 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[4]), .Z(N273) );
  GTECH_AND2 C722 ( .A(fp_op_in[7]), .B(fp_srca_in[4]), .Z(N274) );
  GTECH_OR2 C723 ( .A(N275), .B(N276), .Z(fp_src2_in[3]) );
  GTECH_AND2 C724 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[3]), .Z(N275) );
  GTECH_AND2 C725 ( .A(fp_op_in[7]), .B(fp_srca_in[3]), .Z(N276) );
  GTECH_OR2 C726 ( .A(N277), .B(N278), .Z(fp_src2_in[2]) );
  GTECH_AND2 C727 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[2]), .Z(N277) );
  GTECH_AND2 C728 ( .A(fp_op_in[7]), .B(fp_srca_in[2]), .Z(N278) );
  GTECH_OR2 C729 ( .A(N279), .B(N280), .Z(fp_src2_in[1]) );
  GTECH_AND2 C730 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[1]), .Z(N279) );
  GTECH_AND2 C731 ( .A(fp_op_in[7]), .B(fp_srca_in[1]), .Z(N280) );
  GTECH_OR2 C732 ( .A(N281), .B(N282), .Z(fp_src2_in[0]) );
  GTECH_AND2 C733 ( .A(fp_op_in_7_inv), .B(fp_srcb_in[0]), .Z(N281) );
  GTECH_AND2 C734 ( .A(fp_op_in[7]), .B(fp_srca_in[0]), .Z(N282) );
  GTECH_OR2 C735 ( .A(N283), .B(N287), .Z(inq_id[4]) );
  GTECH_AND2 C736 ( .A(inq_fwrd), .B(fp_id_in[4]), .Z(N283) );
  GTECH_AND2 C737 ( .A(inq_fwrd_inv), .B(N286), .Z(N287) );
  GTECH_OR2 C738 ( .A(N284), .B(N285), .Z(N286) );
  GTECH_AND2 C739 ( .A(inq_bp), .B(inq_din_d1[154]), .Z(N284) );
  GTECH_AND2 C740 ( .A(inq_bp_inv), .B(inq_dout[154]), .Z(N285) );
  GTECH_OR2 C741 ( .A(N288), .B(N292), .Z(inq_id[3]) );
  GTECH_AND2 C742 ( .A(inq_fwrd), .B(fp_id_in[3]), .Z(N288) );
  GTECH_AND2 C743 ( .A(inq_fwrd_inv), .B(N291), .Z(N292) );
  GTECH_OR2 C744 ( .A(N289), .B(N290), .Z(N291) );
  GTECH_AND2 C745 ( .A(inq_bp), .B(inq_din_d1[153]), .Z(N289) );
  GTECH_AND2 C746 ( .A(inq_bp_inv), .B(inq_dout[153]), .Z(N290) );
  GTECH_OR2 C747 ( .A(N293), .B(N297), .Z(inq_id[2]) );
  GTECH_AND2 C748 ( .A(inq_fwrd), .B(fp_id_in[2]), .Z(N293) );
  GTECH_AND2 C749 ( .A(inq_fwrd_inv), .B(N296), .Z(N297) );
  GTECH_OR2 C750 ( .A(N294), .B(N295), .Z(N296) );
  GTECH_AND2 C751 ( .A(inq_bp), .B(inq_din_d1[152]), .Z(N294) );
  GTECH_AND2 C752 ( .A(inq_bp_inv), .B(inq_dout[152]), .Z(N295) );
  GTECH_OR2 C753 ( .A(N298), .B(N302), .Z(inq_id[1]) );
  GTECH_AND2 C754 ( .A(inq_fwrd), .B(fp_id_in[1]), .Z(N298) );
  GTECH_AND2 C755 ( .A(inq_fwrd_inv), .B(N301), .Z(N302) );
  GTECH_OR2 C756 ( .A(N299), .B(N300), .Z(N301) );
  GTECH_AND2 C757 ( .A(inq_bp), .B(inq_din_d1[151]), .Z(N299) );
  GTECH_AND2 C758 ( .A(inq_bp_inv), .B(inq_dout[151]), .Z(N300) );
  GTECH_OR2 C759 ( .A(N303), .B(N307), .Z(inq_id[0]) );
  GTECH_AND2 C760 ( .A(inq_fwrd), .B(fp_id_in[0]), .Z(N303) );
  GTECH_AND2 C761 ( .A(inq_fwrd_inv), .B(N306), .Z(N307) );
  GTECH_OR2 C762 ( .A(N304), .B(N305), .Z(N306) );
  GTECH_AND2 C763 ( .A(inq_bp), .B(inq_din_d1[150]), .Z(N304) );
  GTECH_AND2 C764 ( .A(inq_bp_inv), .B(inq_dout[150]), .Z(N305) );
  GTECH_OR2 C765 ( .A(N308), .B(N312), .Z(inq_rnd_mode[1]) );
  GTECH_AND2 C766 ( .A(inq_fwrd), .B(fp_rnd_mode_in[1]), .Z(N308) );
  GTECH_AND2 C767 ( .A(inq_fwrd_inv), .B(N311), .Z(N312) );
  GTECH_OR2 C768 ( .A(N309), .B(N310), .Z(N311) );
  GTECH_AND2 C769 ( .A(inq_bp), .B(inq_din_d1[149]), .Z(N309) );
  GTECH_AND2 C770 ( .A(inq_bp_inv), .B(inq_dout[149]), .Z(N310) );
  GTECH_OR2 C771 ( .A(N313), .B(N317), .Z(inq_rnd_mode[0]) );
  GTECH_AND2 C772 ( .A(inq_fwrd), .B(fp_rnd_mode_in[0]), .Z(N313) );
  GTECH_AND2 C773 ( .A(inq_fwrd_inv), .B(N316), .Z(N317) );
  GTECH_OR2 C774 ( .A(N314), .B(N315), .Z(N316) );
  GTECH_AND2 C775 ( .A(inq_bp), .B(inq_din_d1[148]), .Z(N314) );
  GTECH_AND2 C776 ( .A(inq_bp_inv), .B(inq_dout[148]), .Z(N315) );
  GTECH_OR2 C777 ( .A(N318), .B(N322), .Z(inq_fcc[1]) );
  GTECH_AND2 C778 ( .A(inq_fwrd), .B(fp_fcc_in[1]), .Z(N318) );
  GTECH_AND2 C779 ( .A(inq_fwrd_inv), .B(N321), .Z(N322) );
  GTECH_OR2 C780 ( .A(N319), .B(N320), .Z(N321) );
  GTECH_AND2 C781 ( .A(inq_bp), .B(inq_din_d1[147]), .Z(N319) );
  GTECH_AND2 C782 ( .A(inq_bp_inv), .B(inq_dout[147]), .Z(N320) );
  GTECH_OR2 C783 ( .A(N323), .B(N327), .Z(inq_fcc[0]) );
  GTECH_AND2 C784 ( .A(inq_fwrd), .B(fp_fcc_in[0]), .Z(N323) );
  GTECH_AND2 C785 ( .A(inq_fwrd_inv), .B(N326), .Z(N327) );
  GTECH_OR2 C786 ( .A(N324), .B(N325), .Z(N326) );
  GTECH_AND2 C787 ( .A(inq_bp), .B(inq_din_d1[146]), .Z(N324) );
  GTECH_AND2 C788 ( .A(inq_bp_inv), .B(inq_dout[146]), .Z(N325) );
  GTECH_OR2 C789 ( .A(N328), .B(N332), .Z(inq_op[7]) );
  GTECH_AND2 C790 ( .A(inq_fwrd), .B(fp_op_in[7]), .Z(N328) );
  GTECH_AND2 C791 ( .A(inq_fwrd_inv), .B(N331), .Z(N332) );
  GTECH_OR2 C792 ( .A(N329), .B(N330), .Z(N331) );
  GTECH_AND2 C793 ( .A(inq_bp), .B(inq_din_d1[145]), .Z(N329) );
  GTECH_AND2 C794 ( .A(inq_bp_inv), .B(inq_dout[145]), .Z(N330) );
  GTECH_OR2 C795 ( .A(N333), .B(N337), .Z(inq_op[6]) );
  GTECH_AND2 C796 ( .A(inq_fwrd), .B(fp_op_in[6]), .Z(N333) );
  GTECH_AND2 C797 ( .A(inq_fwrd_inv), .B(N336), .Z(N337) );
  GTECH_OR2 C798 ( .A(N334), .B(N335), .Z(N336) );
  GTECH_AND2 C799 ( .A(inq_bp), .B(inq_din_d1[144]), .Z(N334) );
  GTECH_AND2 C800 ( .A(inq_bp_inv), .B(inq_dout[144]), .Z(N335) );
  GTECH_OR2 C801 ( .A(N338), .B(N342), .Z(inq_op[5]) );
  GTECH_AND2 C802 ( .A(inq_fwrd), .B(fp_op_in[5]), .Z(N338) );
  GTECH_AND2 C803 ( .A(inq_fwrd_inv), .B(N341), .Z(N342) );
  GTECH_OR2 C804 ( .A(N339), .B(N340), .Z(N341) );
  GTECH_AND2 C805 ( .A(inq_bp), .B(inq_din_d1[143]), .Z(N339) );
  GTECH_AND2 C806 ( .A(inq_bp_inv), .B(inq_dout[143]), .Z(N340) );
  GTECH_OR2 C807 ( .A(N343), .B(N347), .Z(inq_op[4]) );
  GTECH_AND2 C808 ( .A(inq_fwrd), .B(fp_op_in[4]), .Z(N343) );
  GTECH_AND2 C809 ( .A(inq_fwrd_inv), .B(N346), .Z(N347) );
  GTECH_OR2 C810 ( .A(N344), .B(N345), .Z(N346) );
  GTECH_AND2 C811 ( .A(inq_bp), .B(inq_din_d1[142]), .Z(N344) );
  GTECH_AND2 C812 ( .A(inq_bp_inv), .B(inq_dout[142]), .Z(N345) );
  GTECH_OR2 C813 ( .A(N348), .B(N352), .Z(inq_op[3]) );
  GTECH_AND2 C814 ( .A(inq_fwrd), .B(fp_op_in[3]), .Z(N348) );
  GTECH_AND2 C815 ( .A(inq_fwrd_inv), .B(N351), .Z(N352) );
  GTECH_OR2 C816 ( .A(N349), .B(N350), .Z(N351) );
  GTECH_AND2 C817 ( .A(inq_bp), .B(inq_din_d1[141]), .Z(N349) );
  GTECH_AND2 C818 ( .A(inq_bp_inv), .B(inq_dout[141]), .Z(N350) );
  GTECH_OR2 C819 ( .A(N353), .B(N357), .Z(inq_op[2]) );
  GTECH_AND2 C820 ( .A(inq_fwrd), .B(fp_op_in[2]), .Z(N353) );
  GTECH_AND2 C821 ( .A(inq_fwrd_inv), .B(N356), .Z(N357) );
  GTECH_OR2 C822 ( .A(N354), .B(N355), .Z(N356) );
  GTECH_AND2 C823 ( .A(inq_bp), .B(inq_din_d1[140]), .Z(N354) );
  GTECH_AND2 C824 ( .A(inq_bp_inv), .B(inq_dout[140]), .Z(N355) );
  GTECH_OR2 C825 ( .A(N358), .B(N362), .Z(inq_op[1]) );
  GTECH_AND2 C826 ( .A(inq_fwrd), .B(fp_op_in[1]), .Z(N358) );
  GTECH_AND2 C827 ( .A(inq_fwrd_inv), .B(N361), .Z(N362) );
  GTECH_OR2 C828 ( .A(N359), .B(N360), .Z(N361) );
  GTECH_AND2 C829 ( .A(inq_bp), .B(inq_din_d1[139]), .Z(N359) );
  GTECH_AND2 C830 ( .A(inq_bp_inv), .B(inq_dout[139]), .Z(N360) );
  GTECH_OR2 C831 ( .A(N363), .B(N367), .Z(inq_op[0]) );
  GTECH_AND2 C832 ( .A(inq_fwrd), .B(fp_op_in[0]), .Z(N363) );
  GTECH_AND2 C833 ( .A(inq_fwrd_inv), .B(N366), .Z(N367) );
  GTECH_OR2 C834 ( .A(N364), .B(N365), .Z(N366) );
  GTECH_AND2 C835 ( .A(inq_bp), .B(inq_din_d1[138]), .Z(N364) );
  GTECH_AND2 C836 ( .A(inq_bp_inv), .B(inq_dout[138]), .Z(N365) );
  GTECH_OR2 C837 ( .A(N368), .B(N372), .Z(inq_in1_exp_neq_ffs) );
  GTECH_AND2 C838 ( .A(inq_fwrd), .B(fp_src1_in[68]), .Z(N368) );
  GTECH_AND2 C839 ( .A(inq_fwrd_inv), .B(N371), .Z(N372) );
  GTECH_OR2 C840 ( .A(N369), .B(N370), .Z(N371) );
  GTECH_AND2 C841 ( .A(inq_bp), .B(inq_din_d1[137]), .Z(N369) );
  GTECH_AND2 C842 ( .A(inq_bp_inv), .B(inq_dout[137]), .Z(N370) );
  GTECH_OR2 C843 ( .A(N373), .B(N377), .Z(inq_in1_exp_eq_0) );
  GTECH_AND2 C844 ( .A(inq_fwrd), .B(fp_src1_in[67]), .Z(N373) );
  GTECH_AND2 C845 ( .A(inq_fwrd_inv), .B(N376), .Z(N377) );
  GTECH_OR2 C846 ( .A(N374), .B(N375), .Z(N376) );
  GTECH_AND2 C847 ( .A(inq_bp), .B(inq_din_d1[136]), .Z(N374) );
  GTECH_AND2 C848 ( .A(inq_bp_inv), .B(inq_dout[136]), .Z(N375) );
  GTECH_OR2 C849 ( .A(N378), .B(N382), .Z(inq_in1_53_0_neq_0) );
  GTECH_AND2 C850 ( .A(inq_fwrd), .B(fp_src1_in[66]), .Z(N378) );
  GTECH_AND2 C851 ( .A(inq_fwrd_inv), .B(N381), .Z(N382) );
  GTECH_OR2 C852 ( .A(N379), .B(N380), .Z(N381) );
  GTECH_AND2 C853 ( .A(inq_bp), .B(inq_din_d1[135]), .Z(N379) );
  GTECH_AND2 C854 ( .A(inq_bp_inv), .B(inq_dout[135]), .Z(N380) );
  GTECH_OR2 C855 ( .A(N383), .B(N387), .Z(inq_in1_50_0_neq_0) );
  GTECH_AND2 C856 ( .A(inq_fwrd), .B(fp_src1_in[65]), .Z(N383) );
  GTECH_AND2 C857 ( .A(inq_fwrd_inv), .B(N386), .Z(N387) );
  GTECH_OR2 C858 ( .A(N384), .B(N385), .Z(N386) );
  GTECH_AND2 C859 ( .A(inq_bp), .B(inq_din_d1[134]), .Z(N384) );
  GTECH_AND2 C860 ( .A(inq_bp_inv), .B(inq_dout[134]), .Z(N385) );
  GTECH_OR2 C861 ( .A(N388), .B(N392), .Z(inq_in1_53_32_neq_0) );
  GTECH_AND2 C862 ( .A(inq_fwrd), .B(fp_src1_in[64]), .Z(N388) );
  GTECH_AND2 C863 ( .A(inq_fwrd_inv), .B(N391), .Z(N392) );
  GTECH_OR2 C864 ( .A(N389), .B(N390), .Z(N391) );
  GTECH_AND2 C865 ( .A(inq_bp), .B(inq_din_d1[133]), .Z(N389) );
  GTECH_AND2 C866 ( .A(inq_bp_inv), .B(inq_dout[133]), .Z(N390) );
  GTECH_OR2 C867 ( .A(N393), .B(N397), .Z(inq_in1[63]) );
  GTECH_AND2 C868 ( .A(inq_fwrd), .B(fp_src1_in[63]), .Z(N393) );
  GTECH_AND2 C869 ( .A(inq_fwrd_inv), .B(N396), .Z(N397) );
  GTECH_OR2 C870 ( .A(N394), .B(N395), .Z(N396) );
  GTECH_AND2 C871 ( .A(inq_bp), .B(inq_din_d1[132]), .Z(N394) );
  GTECH_AND2 C872 ( .A(inq_bp_inv), .B(inq_dout[132]), .Z(N395) );
  GTECH_OR2 C873 ( .A(N398), .B(N402), .Z(inq_in1[62]) );
  GTECH_AND2 C874 ( .A(inq_fwrd), .B(fp_src1_in[62]), .Z(N398) );
  GTECH_AND2 C875 ( .A(inq_fwrd_inv), .B(N401), .Z(N402) );
  GTECH_OR2 C876 ( .A(N399), .B(N400), .Z(N401) );
  GTECH_AND2 C877 ( .A(inq_bp), .B(inq_din_d1[131]), .Z(N399) );
  GTECH_AND2 C878 ( .A(inq_bp_inv), .B(inq_dout[131]), .Z(N400) );
  GTECH_OR2 C879 ( .A(N403), .B(N407), .Z(inq_in1[61]) );
  GTECH_AND2 C880 ( .A(inq_fwrd), .B(fp_src1_in[61]), .Z(N403) );
  GTECH_AND2 C881 ( .A(inq_fwrd_inv), .B(N406), .Z(N407) );
  GTECH_OR2 C882 ( .A(N404), .B(N405), .Z(N406) );
  GTECH_AND2 C883 ( .A(inq_bp), .B(inq_din_d1[130]), .Z(N404) );
  GTECH_AND2 C884 ( .A(inq_bp_inv), .B(inq_dout[130]), .Z(N405) );
  GTECH_OR2 C885 ( .A(N408), .B(N412), .Z(inq_in1[60]) );
  GTECH_AND2 C886 ( .A(inq_fwrd), .B(fp_src1_in[60]), .Z(N408) );
  GTECH_AND2 C887 ( .A(inq_fwrd_inv), .B(N411), .Z(N412) );
  GTECH_OR2 C888 ( .A(N409), .B(N410), .Z(N411) );
  GTECH_AND2 C889 ( .A(inq_bp), .B(inq_din_d1[129]), .Z(N409) );
  GTECH_AND2 C890 ( .A(inq_bp_inv), .B(inq_dout[129]), .Z(N410) );
  GTECH_OR2 C891 ( .A(N413), .B(N417), .Z(inq_in1[59]) );
  GTECH_AND2 C892 ( .A(inq_fwrd), .B(fp_src1_in[59]), .Z(N413) );
  GTECH_AND2 C893 ( .A(inq_fwrd_inv), .B(N416), .Z(N417) );
  GTECH_OR2 C894 ( .A(N414), .B(N415), .Z(N416) );
  GTECH_AND2 C895 ( .A(inq_bp), .B(inq_din_d1[128]), .Z(N414) );
  GTECH_AND2 C896 ( .A(inq_bp_inv), .B(inq_dout[128]), .Z(N415) );
  GTECH_OR2 C897 ( .A(N418), .B(N422), .Z(inq_in1[58]) );
  GTECH_AND2 C898 ( .A(inq_fwrd), .B(fp_src1_in[58]), .Z(N418) );
  GTECH_AND2 C899 ( .A(inq_fwrd_inv), .B(N421), .Z(N422) );
  GTECH_OR2 C900 ( .A(N419), .B(N420), .Z(N421) );
  GTECH_AND2 C901 ( .A(inq_bp), .B(inq_din_d1[127]), .Z(N419) );
  GTECH_AND2 C902 ( .A(inq_bp_inv), .B(inq_dout[127]), .Z(N420) );
  GTECH_OR2 C903 ( .A(N423), .B(N427), .Z(inq_in1[57]) );
  GTECH_AND2 C904 ( .A(inq_fwrd), .B(fp_src1_in[57]), .Z(N423) );
  GTECH_AND2 C905 ( .A(inq_fwrd_inv), .B(N426), .Z(N427) );
  GTECH_OR2 C906 ( .A(N424), .B(N425), .Z(N426) );
  GTECH_AND2 C907 ( .A(inq_bp), .B(inq_din_d1[126]), .Z(N424) );
  GTECH_AND2 C908 ( .A(inq_bp_inv), .B(inq_dout[126]), .Z(N425) );
  GTECH_OR2 C909 ( .A(N428), .B(N432), .Z(inq_in1[56]) );
  GTECH_AND2 C910 ( .A(inq_fwrd), .B(fp_src1_in[56]), .Z(N428) );
  GTECH_AND2 C911 ( .A(inq_fwrd_inv), .B(N431), .Z(N432) );
  GTECH_OR2 C912 ( .A(N429), .B(N430), .Z(N431) );
  GTECH_AND2 C913 ( .A(inq_bp), .B(inq_din_d1[125]), .Z(N429) );
  GTECH_AND2 C914 ( .A(inq_bp_inv), .B(inq_dout[125]), .Z(N430) );
  GTECH_OR2 C915 ( .A(N433), .B(N437), .Z(inq_in1[55]) );
  GTECH_AND2 C916 ( .A(inq_fwrd), .B(fp_src1_in[55]), .Z(N433) );
  GTECH_AND2 C917 ( .A(inq_fwrd_inv), .B(N436), .Z(N437) );
  GTECH_OR2 C918 ( .A(N434), .B(N435), .Z(N436) );
  GTECH_AND2 C919 ( .A(inq_bp), .B(inq_din_d1[124]), .Z(N434) );
  GTECH_AND2 C920 ( .A(inq_bp_inv), .B(inq_dout[124]), .Z(N435) );
  GTECH_OR2 C921 ( .A(N438), .B(N442), .Z(inq_in1[54]) );
  GTECH_AND2 C922 ( .A(inq_fwrd), .B(fp_src1_in[54]), .Z(N438) );
  GTECH_AND2 C923 ( .A(inq_fwrd_inv), .B(N441), .Z(N442) );
  GTECH_OR2 C924 ( .A(N439), .B(N440), .Z(N441) );
  GTECH_AND2 C925 ( .A(inq_bp), .B(inq_din_d1[123]), .Z(N439) );
  GTECH_AND2 C926 ( .A(inq_bp_inv), .B(inq_dout[123]), .Z(N440) );
  GTECH_OR2 C927 ( .A(N443), .B(N447), .Z(inq_in1[53]) );
  GTECH_AND2 C928 ( .A(inq_fwrd), .B(fp_src1_in[53]), .Z(N443) );
  GTECH_AND2 C929 ( .A(inq_fwrd_inv), .B(N446), .Z(N447) );
  GTECH_OR2 C930 ( .A(N444), .B(N445), .Z(N446) );
  GTECH_AND2 C931 ( .A(inq_bp), .B(inq_din_d1[122]), .Z(N444) );
  GTECH_AND2 C932 ( .A(inq_bp_inv), .B(inq_dout[122]), .Z(N445) );
  GTECH_OR2 C933 ( .A(N448), .B(N452), .Z(inq_in1[52]) );
  GTECH_AND2 C934 ( .A(inq_fwrd), .B(fp_src1_in[52]), .Z(N448) );
  GTECH_AND2 C935 ( .A(inq_fwrd_inv), .B(N451), .Z(N452) );
  GTECH_OR2 C936 ( .A(N449), .B(N450), .Z(N451) );
  GTECH_AND2 C937 ( .A(inq_bp), .B(inq_din_d1[121]), .Z(N449) );
  GTECH_AND2 C938 ( .A(inq_bp_inv), .B(inq_dout[121]), .Z(N450) );
  GTECH_OR2 C939 ( .A(N453), .B(N457), .Z(inq_in1[51]) );
  GTECH_AND2 C940 ( .A(inq_fwrd), .B(fp_src1_in[51]), .Z(N453) );
  GTECH_AND2 C941 ( .A(inq_fwrd_inv), .B(N456), .Z(N457) );
  GTECH_OR2 C942 ( .A(N454), .B(N455), .Z(N456) );
  GTECH_AND2 C943 ( .A(inq_bp), .B(inq_din_d1[120]), .Z(N454) );
  GTECH_AND2 C944 ( .A(inq_bp_inv), .B(inq_dout[120]), .Z(N455) );
  GTECH_OR2 C945 ( .A(N458), .B(N462), .Z(inq_in1[50]) );
  GTECH_AND2 C946 ( .A(inq_fwrd), .B(fp_src1_in[50]), .Z(N458) );
  GTECH_AND2 C947 ( .A(inq_fwrd_inv), .B(N461), .Z(N462) );
  GTECH_OR2 C948 ( .A(N459), .B(N460), .Z(N461) );
  GTECH_AND2 C949 ( .A(inq_bp), .B(inq_din_d1[119]), .Z(N459) );
  GTECH_AND2 C950 ( .A(inq_bp_inv), .B(inq_dout[119]), .Z(N460) );
  GTECH_OR2 C951 ( .A(N463), .B(N467), .Z(inq_in1[49]) );
  GTECH_AND2 C952 ( .A(inq_fwrd), .B(fp_src1_in[49]), .Z(N463) );
  GTECH_AND2 C953 ( .A(inq_fwrd_inv), .B(N466), .Z(N467) );
  GTECH_OR2 C954 ( .A(N464), .B(N465), .Z(N466) );
  GTECH_AND2 C955 ( .A(inq_bp), .B(inq_din_d1[118]), .Z(N464) );
  GTECH_AND2 C956 ( .A(inq_bp_inv), .B(inq_dout[118]), .Z(N465) );
  GTECH_OR2 C957 ( .A(N468), .B(N472), .Z(inq_in1[48]) );
  GTECH_AND2 C958 ( .A(inq_fwrd), .B(fp_src1_in[48]), .Z(N468) );
  GTECH_AND2 C959 ( .A(inq_fwrd_inv), .B(N471), .Z(N472) );
  GTECH_OR2 C960 ( .A(N469), .B(N470), .Z(N471) );
  GTECH_AND2 C961 ( .A(inq_bp), .B(inq_din_d1[117]), .Z(N469) );
  GTECH_AND2 C962 ( .A(inq_bp_inv), .B(inq_dout[117]), .Z(N470) );
  GTECH_OR2 C963 ( .A(N473), .B(N477), .Z(inq_in1[47]) );
  GTECH_AND2 C964 ( .A(inq_fwrd), .B(fp_src1_in[47]), .Z(N473) );
  GTECH_AND2 C965 ( .A(inq_fwrd_inv), .B(N476), .Z(N477) );
  GTECH_OR2 C966 ( .A(N474), .B(N475), .Z(N476) );
  GTECH_AND2 C967 ( .A(inq_bp), .B(inq_din_d1[116]), .Z(N474) );
  GTECH_AND2 C968 ( .A(inq_bp_inv), .B(inq_dout[116]), .Z(N475) );
  GTECH_OR2 C969 ( .A(N478), .B(N482), .Z(inq_in1[46]) );
  GTECH_AND2 C970 ( .A(inq_fwrd), .B(fp_src1_in[46]), .Z(N478) );
  GTECH_AND2 C971 ( .A(inq_fwrd_inv), .B(N481), .Z(N482) );
  GTECH_OR2 C972 ( .A(N479), .B(N480), .Z(N481) );
  GTECH_AND2 C973 ( .A(inq_bp), .B(inq_din_d1[115]), .Z(N479) );
  GTECH_AND2 C974 ( .A(inq_bp_inv), .B(inq_dout[115]), .Z(N480) );
  GTECH_OR2 C975 ( .A(N483), .B(N487), .Z(inq_in1[45]) );
  GTECH_AND2 C976 ( .A(inq_fwrd), .B(fp_src1_in[45]), .Z(N483) );
  GTECH_AND2 C977 ( .A(inq_fwrd_inv), .B(N486), .Z(N487) );
  GTECH_OR2 C978 ( .A(N484), .B(N485), .Z(N486) );
  GTECH_AND2 C979 ( .A(inq_bp), .B(inq_din_d1[114]), .Z(N484) );
  GTECH_AND2 C980 ( .A(inq_bp_inv), .B(inq_dout[114]), .Z(N485) );
  GTECH_OR2 C981 ( .A(N488), .B(N492), .Z(inq_in1[44]) );
  GTECH_AND2 C982 ( .A(inq_fwrd), .B(fp_src1_in[44]), .Z(N488) );
  GTECH_AND2 C983 ( .A(inq_fwrd_inv), .B(N491), .Z(N492) );
  GTECH_OR2 C984 ( .A(N489), .B(N490), .Z(N491) );
  GTECH_AND2 C985 ( .A(inq_bp), .B(inq_din_d1[113]), .Z(N489) );
  GTECH_AND2 C986 ( .A(inq_bp_inv), .B(inq_dout[113]), .Z(N490) );
  GTECH_OR2 C987 ( .A(N493), .B(N497), .Z(inq_in1[43]) );
  GTECH_AND2 C988 ( .A(inq_fwrd), .B(fp_src1_in[43]), .Z(N493) );
  GTECH_AND2 C989 ( .A(inq_fwrd_inv), .B(N496), .Z(N497) );
  GTECH_OR2 C990 ( .A(N494), .B(N495), .Z(N496) );
  GTECH_AND2 C991 ( .A(inq_bp), .B(inq_din_d1[112]), .Z(N494) );
  GTECH_AND2 C992 ( .A(inq_bp_inv), .B(inq_dout[112]), .Z(N495) );
  GTECH_OR2 C993 ( .A(N498), .B(N502), .Z(inq_in1[42]) );
  GTECH_AND2 C994 ( .A(inq_fwrd), .B(fp_src1_in[42]), .Z(N498) );
  GTECH_AND2 C995 ( .A(inq_fwrd_inv), .B(N501), .Z(N502) );
  GTECH_OR2 C996 ( .A(N499), .B(N500), .Z(N501) );
  GTECH_AND2 C997 ( .A(inq_bp), .B(inq_din_d1[111]), .Z(N499) );
  GTECH_AND2 C998 ( .A(inq_bp_inv), .B(inq_dout[111]), .Z(N500) );
  GTECH_OR2 C999 ( .A(N503), .B(N507), .Z(inq_in1[41]) );
  GTECH_AND2 C1000 ( .A(inq_fwrd), .B(fp_src1_in[41]), .Z(N503) );
  GTECH_AND2 C1001 ( .A(inq_fwrd_inv), .B(N506), .Z(N507) );
  GTECH_OR2 C1002 ( .A(N504), .B(N505), .Z(N506) );
  GTECH_AND2 C1003 ( .A(inq_bp), .B(inq_din_d1[110]), .Z(N504) );
  GTECH_AND2 C1004 ( .A(inq_bp_inv), .B(inq_dout[110]), .Z(N505) );
  GTECH_OR2 C1005 ( .A(N508), .B(N512), .Z(inq_in1[40]) );
  GTECH_AND2 C1006 ( .A(inq_fwrd), .B(fp_src1_in[40]), .Z(N508) );
  GTECH_AND2 C1007 ( .A(inq_fwrd_inv), .B(N511), .Z(N512) );
  GTECH_OR2 C1008 ( .A(N509), .B(N510), .Z(N511) );
  GTECH_AND2 C1009 ( .A(inq_bp), .B(inq_din_d1[109]), .Z(N509) );
  GTECH_AND2 C1010 ( .A(inq_bp_inv), .B(inq_dout[109]), .Z(N510) );
  GTECH_OR2 C1011 ( .A(N513), .B(N517), .Z(inq_in1[39]) );
  GTECH_AND2 C1012 ( .A(inq_fwrd), .B(fp_src1_in[39]), .Z(N513) );
  GTECH_AND2 C1013 ( .A(inq_fwrd_inv), .B(N516), .Z(N517) );
  GTECH_OR2 C1014 ( .A(N514), .B(N515), .Z(N516) );
  GTECH_AND2 C1015 ( .A(inq_bp), .B(inq_din_d1[108]), .Z(N514) );
  GTECH_AND2 C1016 ( .A(inq_bp_inv), .B(inq_dout[108]), .Z(N515) );
  GTECH_OR2 C1017 ( .A(N518), .B(N522), .Z(inq_in1[38]) );
  GTECH_AND2 C1018 ( .A(inq_fwrd), .B(fp_src1_in[38]), .Z(N518) );
  GTECH_AND2 C1019 ( .A(inq_fwrd_inv), .B(N521), .Z(N522) );
  GTECH_OR2 C1020 ( .A(N519), .B(N520), .Z(N521) );
  GTECH_AND2 C1021 ( .A(inq_bp), .B(inq_din_d1[107]), .Z(N519) );
  GTECH_AND2 C1022 ( .A(inq_bp_inv), .B(inq_dout[107]), .Z(N520) );
  GTECH_OR2 C1023 ( .A(N523), .B(N527), .Z(inq_in1[37]) );
  GTECH_AND2 C1024 ( .A(inq_fwrd), .B(fp_src1_in[37]), .Z(N523) );
  GTECH_AND2 C1025 ( .A(inq_fwrd_inv), .B(N526), .Z(N527) );
  GTECH_OR2 C1026 ( .A(N524), .B(N525), .Z(N526) );
  GTECH_AND2 C1027 ( .A(inq_bp), .B(inq_din_d1[106]), .Z(N524) );
  GTECH_AND2 C1028 ( .A(inq_bp_inv), .B(inq_dout[106]), .Z(N525) );
  GTECH_OR2 C1029 ( .A(N528), .B(N532), .Z(inq_in1[36]) );
  GTECH_AND2 C1030 ( .A(inq_fwrd), .B(fp_src1_in[36]), .Z(N528) );
  GTECH_AND2 C1031 ( .A(inq_fwrd_inv), .B(N531), .Z(N532) );
  GTECH_OR2 C1032 ( .A(N529), .B(N530), .Z(N531) );
  GTECH_AND2 C1033 ( .A(inq_bp), .B(inq_din_d1[105]), .Z(N529) );
  GTECH_AND2 C1034 ( .A(inq_bp_inv), .B(inq_dout[105]), .Z(N530) );
  GTECH_OR2 C1035 ( .A(N533), .B(N537), .Z(inq_in1[35]) );
  GTECH_AND2 C1036 ( .A(inq_fwrd), .B(fp_src1_in[35]), .Z(N533) );
  GTECH_AND2 C1037 ( .A(inq_fwrd_inv), .B(N536), .Z(N537) );
  GTECH_OR2 C1038 ( .A(N534), .B(N535), .Z(N536) );
  GTECH_AND2 C1039 ( .A(inq_bp), .B(inq_din_d1[104]), .Z(N534) );
  GTECH_AND2 C1040 ( .A(inq_bp_inv), .B(inq_dout[104]), .Z(N535) );
  GTECH_OR2 C1041 ( .A(N538), .B(N542), .Z(inq_in1[34]) );
  GTECH_AND2 C1042 ( .A(inq_fwrd), .B(fp_src1_in[34]), .Z(N538) );
  GTECH_AND2 C1043 ( .A(inq_fwrd_inv), .B(N541), .Z(N542) );
  GTECH_OR2 C1044 ( .A(N539), .B(N540), .Z(N541) );
  GTECH_AND2 C1045 ( .A(inq_bp), .B(inq_din_d1[103]), .Z(N539) );
  GTECH_AND2 C1046 ( .A(inq_bp_inv), .B(inq_dout[103]), .Z(N540) );
  GTECH_OR2 C1047 ( .A(N543), .B(N547), .Z(inq_in1[33]) );
  GTECH_AND2 C1048 ( .A(inq_fwrd), .B(fp_src1_in[33]), .Z(N543) );
  GTECH_AND2 C1049 ( .A(inq_fwrd_inv), .B(N546), .Z(N547) );
  GTECH_OR2 C1050 ( .A(N544), .B(N545), .Z(N546) );
  GTECH_AND2 C1051 ( .A(inq_bp), .B(inq_din_d1[102]), .Z(N544) );
  GTECH_AND2 C1052 ( .A(inq_bp_inv), .B(inq_dout[102]), .Z(N545) );
  GTECH_OR2 C1053 ( .A(N548), .B(N552), .Z(inq_in1[32]) );
  GTECH_AND2 C1054 ( .A(inq_fwrd), .B(fp_src1_in[32]), .Z(N548) );
  GTECH_AND2 C1055 ( .A(inq_fwrd_inv), .B(N551), .Z(N552) );
  GTECH_OR2 C1056 ( .A(N549), .B(N550), .Z(N551) );
  GTECH_AND2 C1057 ( .A(inq_bp), .B(inq_din_d1[101]), .Z(N549) );
  GTECH_AND2 C1058 ( .A(inq_bp_inv), .B(inq_dout[101]), .Z(N550) );
  GTECH_OR2 C1059 ( .A(N553), .B(N557), .Z(inq_in1[31]) );
  GTECH_AND2 C1060 ( .A(inq_fwrd), .B(fp_src1_in[31]), .Z(N553) );
  GTECH_AND2 C1061 ( .A(inq_fwrd_inv), .B(N556), .Z(N557) );
  GTECH_OR2 C1062 ( .A(N554), .B(N555), .Z(N556) );
  GTECH_AND2 C1063 ( .A(inq_bp), .B(inq_din_d1[100]), .Z(N554) );
  GTECH_AND2 C1064 ( .A(inq_bp_inv), .B(inq_dout[100]), .Z(N555) );
  GTECH_OR2 C1065 ( .A(N558), .B(N562), .Z(inq_in1[30]) );
  GTECH_AND2 C1066 ( .A(inq_fwrd), .B(fp_src1_in[30]), .Z(N558) );
  GTECH_AND2 C1067 ( .A(inq_fwrd_inv), .B(N561), .Z(N562) );
  GTECH_OR2 C1068 ( .A(N559), .B(N560), .Z(N561) );
  GTECH_AND2 C1069 ( .A(inq_bp), .B(inq_din_d1[99]), .Z(N559) );
  GTECH_AND2 C1070 ( .A(inq_bp_inv), .B(inq_dout[99]), .Z(N560) );
  GTECH_OR2 C1071 ( .A(N563), .B(N567), .Z(inq_in1[29]) );
  GTECH_AND2 C1072 ( .A(inq_fwrd), .B(fp_src1_in[29]), .Z(N563) );
  GTECH_AND2 C1073 ( .A(inq_fwrd_inv), .B(N566), .Z(N567) );
  GTECH_OR2 C1074 ( .A(N564), .B(N565), .Z(N566) );
  GTECH_AND2 C1075 ( .A(inq_bp), .B(inq_din_d1[98]), .Z(N564) );
  GTECH_AND2 C1076 ( .A(inq_bp_inv), .B(inq_dout[98]), .Z(N565) );
  GTECH_OR2 C1077 ( .A(N568), .B(N572), .Z(inq_in1[28]) );
  GTECH_AND2 C1078 ( .A(inq_fwrd), .B(fp_src1_in[28]), .Z(N568) );
  GTECH_AND2 C1079 ( .A(inq_fwrd_inv), .B(N571), .Z(N572) );
  GTECH_OR2 C1080 ( .A(N569), .B(N570), .Z(N571) );
  GTECH_AND2 C1081 ( .A(inq_bp), .B(inq_din_d1[97]), .Z(N569) );
  GTECH_AND2 C1082 ( .A(inq_bp_inv), .B(inq_dout[97]), .Z(N570) );
  GTECH_OR2 C1083 ( .A(N573), .B(N577), .Z(inq_in1[27]) );
  GTECH_AND2 C1084 ( .A(inq_fwrd), .B(fp_src1_in[27]), .Z(N573) );
  GTECH_AND2 C1085 ( .A(inq_fwrd_inv), .B(N576), .Z(N577) );
  GTECH_OR2 C1086 ( .A(N574), .B(N575), .Z(N576) );
  GTECH_AND2 C1087 ( .A(inq_bp), .B(inq_din_d1[96]), .Z(N574) );
  GTECH_AND2 C1088 ( .A(inq_bp_inv), .B(inq_dout[96]), .Z(N575) );
  GTECH_OR2 C1089 ( .A(N578), .B(N582), .Z(inq_in1[26]) );
  GTECH_AND2 C1090 ( .A(inq_fwrd), .B(fp_src1_in[26]), .Z(N578) );
  GTECH_AND2 C1091 ( .A(inq_fwrd_inv), .B(N581), .Z(N582) );
  GTECH_OR2 C1092 ( .A(N579), .B(N580), .Z(N581) );
  GTECH_AND2 C1093 ( .A(inq_bp), .B(inq_din_d1[95]), .Z(N579) );
  GTECH_AND2 C1094 ( .A(inq_bp_inv), .B(inq_dout[95]), .Z(N580) );
  GTECH_OR2 C1095 ( .A(N583), .B(N587), .Z(inq_in1[25]) );
  GTECH_AND2 C1096 ( .A(inq_fwrd), .B(fp_src1_in[25]), .Z(N583) );
  GTECH_AND2 C1097 ( .A(inq_fwrd_inv), .B(N586), .Z(N587) );
  GTECH_OR2 C1098 ( .A(N584), .B(N585), .Z(N586) );
  GTECH_AND2 C1099 ( .A(inq_bp), .B(inq_din_d1[94]), .Z(N584) );
  GTECH_AND2 C1100 ( .A(inq_bp_inv), .B(inq_dout[94]), .Z(N585) );
  GTECH_OR2 C1101 ( .A(N588), .B(N592), .Z(inq_in1[24]) );
  GTECH_AND2 C1102 ( .A(inq_fwrd), .B(fp_src1_in[24]), .Z(N588) );
  GTECH_AND2 C1103 ( .A(inq_fwrd_inv), .B(N591), .Z(N592) );
  GTECH_OR2 C1104 ( .A(N589), .B(N590), .Z(N591) );
  GTECH_AND2 C1105 ( .A(inq_bp), .B(inq_din_d1[93]), .Z(N589) );
  GTECH_AND2 C1106 ( .A(inq_bp_inv), .B(inq_dout[93]), .Z(N590) );
  GTECH_OR2 C1107 ( .A(N593), .B(N597), .Z(inq_in1[23]) );
  GTECH_AND2 C1108 ( .A(inq_fwrd), .B(fp_src1_in[23]), .Z(N593) );
  GTECH_AND2 C1109 ( .A(inq_fwrd_inv), .B(N596), .Z(N597) );
  GTECH_OR2 C1110 ( .A(N594), .B(N595), .Z(N596) );
  GTECH_AND2 C1111 ( .A(inq_bp), .B(inq_din_d1[92]), .Z(N594) );
  GTECH_AND2 C1112 ( .A(inq_bp_inv), .B(inq_dout[92]), .Z(N595) );
  GTECH_OR2 C1113 ( .A(N598), .B(N602), .Z(inq_in1[22]) );
  GTECH_AND2 C1114 ( .A(inq_fwrd), .B(fp_src1_in[22]), .Z(N598) );
  GTECH_AND2 C1115 ( .A(inq_fwrd_inv), .B(N601), .Z(N602) );
  GTECH_OR2 C1116 ( .A(N599), .B(N600), .Z(N601) );
  GTECH_AND2 C1117 ( .A(inq_bp), .B(inq_din_d1[91]), .Z(N599) );
  GTECH_AND2 C1118 ( .A(inq_bp_inv), .B(inq_dout[91]), .Z(N600) );
  GTECH_OR2 C1119 ( .A(N603), .B(N607), .Z(inq_in1[21]) );
  GTECH_AND2 C1120 ( .A(inq_fwrd), .B(fp_src1_in[21]), .Z(N603) );
  GTECH_AND2 C1121 ( .A(inq_fwrd_inv), .B(N606), .Z(N607) );
  GTECH_OR2 C1122 ( .A(N604), .B(N605), .Z(N606) );
  GTECH_AND2 C1123 ( .A(inq_bp), .B(inq_din_d1[90]), .Z(N604) );
  GTECH_AND2 C1124 ( .A(inq_bp_inv), .B(inq_dout[90]), .Z(N605) );
  GTECH_OR2 C1125 ( .A(N608), .B(N612), .Z(inq_in1[20]) );
  GTECH_AND2 C1126 ( .A(inq_fwrd), .B(fp_src1_in[20]), .Z(N608) );
  GTECH_AND2 C1127 ( .A(inq_fwrd_inv), .B(N611), .Z(N612) );
  GTECH_OR2 C1128 ( .A(N609), .B(N610), .Z(N611) );
  GTECH_AND2 C1129 ( .A(inq_bp), .B(inq_din_d1[89]), .Z(N609) );
  GTECH_AND2 C1130 ( .A(inq_bp_inv), .B(inq_dout[89]), .Z(N610) );
  GTECH_OR2 C1131 ( .A(N613), .B(N617), .Z(inq_in1[19]) );
  GTECH_AND2 C1132 ( .A(inq_fwrd), .B(fp_src1_in[19]), .Z(N613) );
  GTECH_AND2 C1133 ( .A(inq_fwrd_inv), .B(N616), .Z(N617) );
  GTECH_OR2 C1134 ( .A(N614), .B(N615), .Z(N616) );
  GTECH_AND2 C1135 ( .A(inq_bp), .B(inq_din_d1[88]), .Z(N614) );
  GTECH_AND2 C1136 ( .A(inq_bp_inv), .B(inq_dout[88]), .Z(N615) );
  GTECH_OR2 C1137 ( .A(N618), .B(N622), .Z(inq_in1[18]) );
  GTECH_AND2 C1138 ( .A(inq_fwrd), .B(fp_src1_in[18]), .Z(N618) );
  GTECH_AND2 C1139 ( .A(inq_fwrd_inv), .B(N621), .Z(N622) );
  GTECH_OR2 C1140 ( .A(N619), .B(N620), .Z(N621) );
  GTECH_AND2 C1141 ( .A(inq_bp), .B(inq_din_d1[87]), .Z(N619) );
  GTECH_AND2 C1142 ( .A(inq_bp_inv), .B(inq_dout[87]), .Z(N620) );
  GTECH_OR2 C1143 ( .A(N623), .B(N627), .Z(inq_in1[17]) );
  GTECH_AND2 C1144 ( .A(inq_fwrd), .B(fp_src1_in[17]), .Z(N623) );
  GTECH_AND2 C1145 ( .A(inq_fwrd_inv), .B(N626), .Z(N627) );
  GTECH_OR2 C1146 ( .A(N624), .B(N625), .Z(N626) );
  GTECH_AND2 C1147 ( .A(inq_bp), .B(inq_din_d1[86]), .Z(N624) );
  GTECH_AND2 C1148 ( .A(inq_bp_inv), .B(inq_dout[86]), .Z(N625) );
  GTECH_OR2 C1149 ( .A(N628), .B(N632), .Z(inq_in1[16]) );
  GTECH_AND2 C1150 ( .A(inq_fwrd), .B(fp_src1_in[16]), .Z(N628) );
  GTECH_AND2 C1151 ( .A(inq_fwrd_inv), .B(N631), .Z(N632) );
  GTECH_OR2 C1152 ( .A(N629), .B(N630), .Z(N631) );
  GTECH_AND2 C1153 ( .A(inq_bp), .B(inq_din_d1[85]), .Z(N629) );
  GTECH_AND2 C1154 ( .A(inq_bp_inv), .B(inq_dout[85]), .Z(N630) );
  GTECH_OR2 C1155 ( .A(N633), .B(N637), .Z(inq_in1[15]) );
  GTECH_AND2 C1156 ( .A(inq_fwrd), .B(fp_src1_in[15]), .Z(N633) );
  GTECH_AND2 C1157 ( .A(inq_fwrd_inv), .B(N636), .Z(N637) );
  GTECH_OR2 C1158 ( .A(N634), .B(N635), .Z(N636) );
  GTECH_AND2 C1159 ( .A(inq_bp), .B(inq_din_d1[84]), .Z(N634) );
  GTECH_AND2 C1160 ( .A(inq_bp_inv), .B(inq_dout[84]), .Z(N635) );
  GTECH_OR2 C1161 ( .A(N638), .B(N642), .Z(inq_in1[14]) );
  GTECH_AND2 C1162 ( .A(inq_fwrd), .B(fp_src1_in[14]), .Z(N638) );
  GTECH_AND2 C1163 ( .A(inq_fwrd_inv), .B(N641), .Z(N642) );
  GTECH_OR2 C1164 ( .A(N639), .B(N640), .Z(N641) );
  GTECH_AND2 C1165 ( .A(inq_bp), .B(inq_din_d1[83]), .Z(N639) );
  GTECH_AND2 C1166 ( .A(inq_bp_inv), .B(inq_dout[83]), .Z(N640) );
  GTECH_OR2 C1167 ( .A(N643), .B(N647), .Z(inq_in1[13]) );
  GTECH_AND2 C1168 ( .A(inq_fwrd), .B(fp_src1_in[13]), .Z(N643) );
  GTECH_AND2 C1169 ( .A(inq_fwrd_inv), .B(N646), .Z(N647) );
  GTECH_OR2 C1170 ( .A(N644), .B(N645), .Z(N646) );
  GTECH_AND2 C1171 ( .A(inq_bp), .B(inq_din_d1[82]), .Z(N644) );
  GTECH_AND2 C1172 ( .A(inq_bp_inv), .B(inq_dout[82]), .Z(N645) );
  GTECH_OR2 C1173 ( .A(N648), .B(N652), .Z(inq_in1[12]) );
  GTECH_AND2 C1174 ( .A(inq_fwrd), .B(fp_src1_in[12]), .Z(N648) );
  GTECH_AND2 C1175 ( .A(inq_fwrd_inv), .B(N651), .Z(N652) );
  GTECH_OR2 C1176 ( .A(N649), .B(N650), .Z(N651) );
  GTECH_AND2 C1177 ( .A(inq_bp), .B(inq_din_d1[81]), .Z(N649) );
  GTECH_AND2 C1178 ( .A(inq_bp_inv), .B(inq_dout[81]), .Z(N650) );
  GTECH_OR2 C1179 ( .A(N653), .B(N657), .Z(inq_in1[11]) );
  GTECH_AND2 C1180 ( .A(inq_fwrd), .B(fp_src1_in[11]), .Z(N653) );
  GTECH_AND2 C1181 ( .A(inq_fwrd_inv), .B(N656), .Z(N657) );
  GTECH_OR2 C1182 ( .A(N654), .B(N655), .Z(N656) );
  GTECH_AND2 C1183 ( .A(inq_bp), .B(inq_din_d1[80]), .Z(N654) );
  GTECH_AND2 C1184 ( .A(inq_bp_inv), .B(inq_dout[80]), .Z(N655) );
  GTECH_OR2 C1185 ( .A(N658), .B(N662), .Z(inq_in1[10]) );
  GTECH_AND2 C1186 ( .A(inq_fwrd), .B(fp_src1_in[10]), .Z(N658) );
  GTECH_AND2 C1187 ( .A(inq_fwrd_inv), .B(N661), .Z(N662) );
  GTECH_OR2 C1188 ( .A(N659), .B(N660), .Z(N661) );
  GTECH_AND2 C1189 ( .A(inq_bp), .B(inq_din_d1[79]), .Z(N659) );
  GTECH_AND2 C1190 ( .A(inq_bp_inv), .B(inq_dout[79]), .Z(N660) );
  GTECH_OR2 C1191 ( .A(N663), .B(N667), .Z(inq_in1[9]) );
  GTECH_AND2 C1192 ( .A(inq_fwrd), .B(fp_src1_in[9]), .Z(N663) );
  GTECH_AND2 C1193 ( .A(inq_fwrd_inv), .B(N666), .Z(N667) );
  GTECH_OR2 C1194 ( .A(N664), .B(N665), .Z(N666) );
  GTECH_AND2 C1195 ( .A(inq_bp), .B(inq_din_d1[78]), .Z(N664) );
  GTECH_AND2 C1196 ( .A(inq_bp_inv), .B(inq_dout[78]), .Z(N665) );
  GTECH_OR2 C1197 ( .A(N668), .B(N672), .Z(inq_in1[8]) );
  GTECH_AND2 C1198 ( .A(inq_fwrd), .B(fp_src1_in[8]), .Z(N668) );
  GTECH_AND2 C1199 ( .A(inq_fwrd_inv), .B(N671), .Z(N672) );
  GTECH_OR2 C1200 ( .A(N669), .B(N670), .Z(N671) );
  GTECH_AND2 C1201 ( .A(inq_bp), .B(inq_din_d1[77]), .Z(N669) );
  GTECH_AND2 C1202 ( .A(inq_bp_inv), .B(inq_dout[77]), .Z(N670) );
  GTECH_OR2 C1203 ( .A(N673), .B(N677), .Z(inq_in1[7]) );
  GTECH_AND2 C1204 ( .A(inq_fwrd), .B(fp_src1_in[7]), .Z(N673) );
  GTECH_AND2 C1205 ( .A(inq_fwrd_inv), .B(N676), .Z(N677) );
  GTECH_OR2 C1206 ( .A(N674), .B(N675), .Z(N676) );
  GTECH_AND2 C1207 ( .A(inq_bp), .B(inq_din_d1[76]), .Z(N674) );
  GTECH_AND2 C1208 ( .A(inq_bp_inv), .B(inq_dout[76]), .Z(N675) );
  GTECH_OR2 C1209 ( .A(N678), .B(N682), .Z(inq_in1[6]) );
  GTECH_AND2 C1210 ( .A(inq_fwrd), .B(fp_src1_in[6]), .Z(N678) );
  GTECH_AND2 C1211 ( .A(inq_fwrd_inv), .B(N681), .Z(N682) );
  GTECH_OR2 C1212 ( .A(N679), .B(N680), .Z(N681) );
  GTECH_AND2 C1213 ( .A(inq_bp), .B(inq_din_d1[75]), .Z(N679) );
  GTECH_AND2 C1214 ( .A(inq_bp_inv), .B(inq_dout[75]), .Z(N680) );
  GTECH_OR2 C1215 ( .A(N683), .B(N687), .Z(inq_in1[5]) );
  GTECH_AND2 C1216 ( .A(inq_fwrd), .B(fp_src1_in[5]), .Z(N683) );
  GTECH_AND2 C1217 ( .A(inq_fwrd_inv), .B(N686), .Z(N687) );
  GTECH_OR2 C1218 ( .A(N684), .B(N685), .Z(N686) );
  GTECH_AND2 C1219 ( .A(inq_bp), .B(inq_din_d1[74]), .Z(N684) );
  GTECH_AND2 C1220 ( .A(inq_bp_inv), .B(inq_dout[74]), .Z(N685) );
  GTECH_OR2 C1221 ( .A(N688), .B(N692), .Z(inq_in1[4]) );
  GTECH_AND2 C1222 ( .A(inq_fwrd), .B(fp_src1_in[4]), .Z(N688) );
  GTECH_AND2 C1223 ( .A(inq_fwrd_inv), .B(N691), .Z(N692) );
  GTECH_OR2 C1224 ( .A(N689), .B(N690), .Z(N691) );
  GTECH_AND2 C1225 ( .A(inq_bp), .B(inq_din_d1[73]), .Z(N689) );
  GTECH_AND2 C1226 ( .A(inq_bp_inv), .B(inq_dout[73]), .Z(N690) );
  GTECH_OR2 C1227 ( .A(N693), .B(N697), .Z(inq_in1[3]) );
  GTECH_AND2 C1228 ( .A(inq_fwrd), .B(fp_src1_in[3]), .Z(N693) );
  GTECH_AND2 C1229 ( .A(inq_fwrd_inv), .B(N696), .Z(N697) );
  GTECH_OR2 C1230 ( .A(N694), .B(N695), .Z(N696) );
  GTECH_AND2 C1231 ( .A(inq_bp), .B(inq_din_d1[72]), .Z(N694) );
  GTECH_AND2 C1232 ( .A(inq_bp_inv), .B(inq_dout[72]), .Z(N695) );
  GTECH_OR2 C1233 ( .A(N698), .B(N702), .Z(inq_in1[2]) );
  GTECH_AND2 C1234 ( .A(inq_fwrd), .B(fp_src1_in[2]), .Z(N698) );
  GTECH_AND2 C1235 ( .A(inq_fwrd_inv), .B(N701), .Z(N702) );
  GTECH_OR2 C1236 ( .A(N699), .B(N700), .Z(N701) );
  GTECH_AND2 C1237 ( .A(inq_bp), .B(inq_din_d1[71]), .Z(N699) );
  GTECH_AND2 C1238 ( .A(inq_bp_inv), .B(inq_dout[71]), .Z(N700) );
  GTECH_OR2 C1239 ( .A(N703), .B(N707), .Z(inq_in1[1]) );
  GTECH_AND2 C1240 ( .A(inq_fwrd), .B(fp_src1_in[1]), .Z(N703) );
  GTECH_AND2 C1241 ( .A(inq_fwrd_inv), .B(N706), .Z(N707) );
  GTECH_OR2 C1242 ( .A(N704), .B(N705), .Z(N706) );
  GTECH_AND2 C1243 ( .A(inq_bp), .B(inq_din_d1[70]), .Z(N704) );
  GTECH_AND2 C1244 ( .A(inq_bp_inv), .B(inq_dout[70]), .Z(N705) );
  GTECH_OR2 C1245 ( .A(N708), .B(N712), .Z(inq_in1[0]) );
  GTECH_AND2 C1246 ( .A(inq_fwrd), .B(fp_src1_in[0]), .Z(N708) );
  GTECH_AND2 C1247 ( .A(inq_fwrd_inv), .B(N711), .Z(N712) );
  GTECH_OR2 C1248 ( .A(N709), .B(N710), .Z(N711) );
  GTECH_AND2 C1249 ( .A(inq_bp), .B(inq_din_d1[69]), .Z(N709) );
  GTECH_AND2 C1250 ( .A(inq_bp_inv), .B(inq_dout[69]), .Z(N710) );
  GTECH_OR2 C1251 ( .A(N713), .B(N717), .Z(inq_in2_exp_neq_ffs) );
  GTECH_AND2 C1252 ( .A(inq_fwrd), .B(fp_src2_in[68]), .Z(N713) );
  GTECH_AND2 C1253 ( .A(inq_fwrd_inv), .B(N716), .Z(N717) );
  GTECH_OR2 C1254 ( .A(N714), .B(N715), .Z(N716) );
  GTECH_AND2 C1255 ( .A(inq_bp), .B(inq_din_d1[68]), .Z(N714) );
  GTECH_AND2 C1256 ( .A(inq_bp_inv), .B(inq_dout[68]), .Z(N715) );
  GTECH_OR2 C1257 ( .A(N718), .B(N722), .Z(inq_in2_exp_eq_0) );
  GTECH_AND2 C1258 ( .A(inq_fwrd), .B(fp_src2_in[67]), .Z(N718) );
  GTECH_AND2 C1259 ( .A(inq_fwrd_inv), .B(N721), .Z(N722) );
  GTECH_OR2 C1260 ( .A(N719), .B(N720), .Z(N721) );
  GTECH_AND2 C1261 ( .A(inq_bp), .B(inq_din_d1[67]), .Z(N719) );
  GTECH_AND2 C1262 ( .A(inq_bp_inv), .B(inq_dout[67]), .Z(N720) );
  GTECH_OR2 C1263 ( .A(N723), .B(N727), .Z(inq_in2_53_0_neq_0) );
  GTECH_AND2 C1264 ( .A(inq_fwrd), .B(fp_src2_in[66]), .Z(N723) );
  GTECH_AND2 C1265 ( .A(inq_fwrd_inv), .B(N726), .Z(N727) );
  GTECH_OR2 C1266 ( .A(N724), .B(N725), .Z(N726) );
  GTECH_AND2 C1267 ( .A(inq_bp), .B(inq_din_d1[66]), .Z(N724) );
  GTECH_AND2 C1268 ( .A(inq_bp_inv), .B(inq_dout[66]), .Z(N725) );
  GTECH_OR2 C1269 ( .A(N728), .B(N732), .Z(inq_in2_50_0_neq_0) );
  GTECH_AND2 C1270 ( .A(inq_fwrd), .B(fp_src2_in[65]), .Z(N728) );
  GTECH_AND2 C1271 ( .A(inq_fwrd_inv), .B(N731), .Z(N732) );
  GTECH_OR2 C1272 ( .A(N729), .B(N730), .Z(N731) );
  GTECH_AND2 C1273 ( .A(inq_bp), .B(inq_din_d1[65]), .Z(N729) );
  GTECH_AND2 C1274 ( .A(inq_bp_inv), .B(inq_dout[65]), .Z(N730) );
  GTECH_OR2 C1275 ( .A(N733), .B(N737), .Z(inq_in2_53_32_neq_0) );
  GTECH_AND2 C1276 ( .A(inq_fwrd), .B(fp_src2_in[64]), .Z(N733) );
  GTECH_AND2 C1277 ( .A(inq_fwrd_inv), .B(N736), .Z(N737) );
  GTECH_OR2 C1278 ( .A(N734), .B(N735), .Z(N736) );
  GTECH_AND2 C1279 ( .A(inq_bp), .B(inq_din_d1[64]), .Z(N734) );
  GTECH_AND2 C1280 ( .A(inq_bp_inv), .B(inq_dout[64]), .Z(N735) );
  GTECH_OR2 C1281 ( .A(N738), .B(N742), .Z(inq_in2[63]) );
  GTECH_AND2 C1282 ( .A(inq_fwrd), .B(fp_src2_in[63]), .Z(N738) );
  GTECH_AND2 C1283 ( .A(inq_fwrd_inv), .B(N741), .Z(N742) );
  GTECH_OR2 C1284 ( .A(N739), .B(N740), .Z(N741) );
  GTECH_AND2 C1285 ( .A(inq_bp), .B(inq_din_d1[63]), .Z(N739) );
  GTECH_AND2 C1286 ( .A(inq_bp_inv), .B(inq_dout[63]), .Z(N740) );
  GTECH_OR2 C1287 ( .A(N743), .B(N747), .Z(inq_in2[62]) );
  GTECH_AND2 C1288 ( .A(inq_fwrd), .B(fp_src2_in[62]), .Z(N743) );
  GTECH_AND2 C1289 ( .A(inq_fwrd_inv), .B(N746), .Z(N747) );
  GTECH_OR2 C1290 ( .A(N744), .B(N745), .Z(N746) );
  GTECH_AND2 C1291 ( .A(inq_bp), .B(inq_din_d1[62]), .Z(N744) );
  GTECH_AND2 C1292 ( .A(inq_bp_inv), .B(inq_dout[62]), .Z(N745) );
  GTECH_OR2 C1293 ( .A(N748), .B(N752), .Z(inq_in2[61]) );
  GTECH_AND2 C1294 ( .A(inq_fwrd), .B(fp_src2_in[61]), .Z(N748) );
  GTECH_AND2 C1295 ( .A(inq_fwrd_inv), .B(N751), .Z(N752) );
  GTECH_OR2 C1296 ( .A(N749), .B(N750), .Z(N751) );
  GTECH_AND2 C1297 ( .A(inq_bp), .B(inq_din_d1[61]), .Z(N749) );
  GTECH_AND2 C1298 ( .A(inq_bp_inv), .B(inq_dout[61]), .Z(N750) );
  GTECH_OR2 C1299 ( .A(N753), .B(N757), .Z(inq_in2[60]) );
  GTECH_AND2 C1300 ( .A(inq_fwrd), .B(fp_src2_in[60]), .Z(N753) );
  GTECH_AND2 C1301 ( .A(inq_fwrd_inv), .B(N756), .Z(N757) );
  GTECH_OR2 C1302 ( .A(N754), .B(N755), .Z(N756) );
  GTECH_AND2 C1303 ( .A(inq_bp), .B(inq_din_d1[60]), .Z(N754) );
  GTECH_AND2 C1304 ( .A(inq_bp_inv), .B(inq_dout[60]), .Z(N755) );
  GTECH_OR2 C1305 ( .A(N758), .B(N762), .Z(inq_in2[59]) );
  GTECH_AND2 C1306 ( .A(inq_fwrd), .B(fp_src2_in[59]), .Z(N758) );
  GTECH_AND2 C1307 ( .A(inq_fwrd_inv), .B(N761), .Z(N762) );
  GTECH_OR2 C1308 ( .A(N759), .B(N760), .Z(N761) );
  GTECH_AND2 C1309 ( .A(inq_bp), .B(inq_din_d1[59]), .Z(N759) );
  GTECH_AND2 C1310 ( .A(inq_bp_inv), .B(inq_dout[59]), .Z(N760) );
  GTECH_OR2 C1311 ( .A(N763), .B(N767), .Z(inq_in2[58]) );
  GTECH_AND2 C1312 ( .A(inq_fwrd), .B(fp_src2_in[58]), .Z(N763) );
  GTECH_AND2 C1313 ( .A(inq_fwrd_inv), .B(N766), .Z(N767) );
  GTECH_OR2 C1314 ( .A(N764), .B(N765), .Z(N766) );
  GTECH_AND2 C1315 ( .A(inq_bp), .B(inq_din_d1[58]), .Z(N764) );
  GTECH_AND2 C1316 ( .A(inq_bp_inv), .B(inq_dout[58]), .Z(N765) );
  GTECH_OR2 C1317 ( .A(N768), .B(N772), .Z(inq_in2[57]) );
  GTECH_AND2 C1318 ( .A(inq_fwrd), .B(fp_src2_in[57]), .Z(N768) );
  GTECH_AND2 C1319 ( .A(inq_fwrd_inv), .B(N771), .Z(N772) );
  GTECH_OR2 C1320 ( .A(N769), .B(N770), .Z(N771) );
  GTECH_AND2 C1321 ( .A(inq_bp), .B(inq_din_d1[57]), .Z(N769) );
  GTECH_AND2 C1322 ( .A(inq_bp_inv), .B(inq_dout[57]), .Z(N770) );
  GTECH_OR2 C1323 ( .A(N773), .B(N777), .Z(inq_in2[56]) );
  GTECH_AND2 C1324 ( .A(inq_fwrd), .B(fp_src2_in[56]), .Z(N773) );
  GTECH_AND2 C1325 ( .A(inq_fwrd_inv), .B(N776), .Z(N777) );
  GTECH_OR2 C1326 ( .A(N774), .B(N775), .Z(N776) );
  GTECH_AND2 C1327 ( .A(inq_bp), .B(inq_din_d1[56]), .Z(N774) );
  GTECH_AND2 C1328 ( .A(inq_bp_inv), .B(inq_dout[56]), .Z(N775) );
  GTECH_OR2 C1329 ( .A(N778), .B(N782), .Z(inq_in2[55]) );
  GTECH_AND2 C1330 ( .A(inq_fwrd), .B(fp_src2_in[55]), .Z(N778) );
  GTECH_AND2 C1331 ( .A(inq_fwrd_inv), .B(N781), .Z(N782) );
  GTECH_OR2 C1332 ( .A(N779), .B(N780), .Z(N781) );
  GTECH_AND2 C1333 ( .A(inq_bp), .B(inq_din_d1[55]), .Z(N779) );
  GTECH_AND2 C1334 ( .A(inq_bp_inv), .B(inq_dout[55]), .Z(N780) );
  GTECH_OR2 C1335 ( .A(N783), .B(N787), .Z(inq_in2[54]) );
  GTECH_AND2 C1336 ( .A(inq_fwrd), .B(fp_src2_in[54]), .Z(N783) );
  GTECH_AND2 C1337 ( .A(inq_fwrd_inv), .B(N786), .Z(N787) );
  GTECH_OR2 C1338 ( .A(N784), .B(N785), .Z(N786) );
  GTECH_AND2 C1339 ( .A(inq_bp), .B(inq_din_d1[54]), .Z(N784) );
  GTECH_AND2 C1340 ( .A(inq_bp_inv), .B(inq_dout[54]), .Z(N785) );
  GTECH_OR2 C1341 ( .A(N788), .B(N792), .Z(inq_in2[53]) );
  GTECH_AND2 C1342 ( .A(inq_fwrd), .B(fp_src2_in[53]), .Z(N788) );
  GTECH_AND2 C1343 ( .A(inq_fwrd_inv), .B(N791), .Z(N792) );
  GTECH_OR2 C1344 ( .A(N789), .B(N790), .Z(N791) );
  GTECH_AND2 C1345 ( .A(inq_bp), .B(inq_din_d1[53]), .Z(N789) );
  GTECH_AND2 C1346 ( .A(inq_bp_inv), .B(inq_dout[53]), .Z(N790) );
  GTECH_OR2 C1347 ( .A(N793), .B(N797), .Z(inq_in2[52]) );
  GTECH_AND2 C1348 ( .A(inq_fwrd), .B(fp_src2_in[52]), .Z(N793) );
  GTECH_AND2 C1349 ( .A(inq_fwrd_inv), .B(N796), .Z(N797) );
  GTECH_OR2 C1350 ( .A(N794), .B(N795), .Z(N796) );
  GTECH_AND2 C1351 ( .A(inq_bp), .B(inq_din_d1[52]), .Z(N794) );
  GTECH_AND2 C1352 ( .A(inq_bp_inv), .B(inq_dout[52]), .Z(N795) );
  GTECH_OR2 C1353 ( .A(N798), .B(N802), .Z(inq_in2[51]) );
  GTECH_AND2 C1354 ( .A(inq_fwrd), .B(fp_src2_in[51]), .Z(N798) );
  GTECH_AND2 C1355 ( .A(inq_fwrd_inv), .B(N801), .Z(N802) );
  GTECH_OR2 C1356 ( .A(N799), .B(N800), .Z(N801) );
  GTECH_AND2 C1357 ( .A(inq_bp), .B(inq_din_d1[51]), .Z(N799) );
  GTECH_AND2 C1358 ( .A(inq_bp_inv), .B(inq_dout[51]), .Z(N800) );
  GTECH_OR2 C1359 ( .A(N803), .B(N807), .Z(inq_in2[50]) );
  GTECH_AND2 C1360 ( .A(inq_fwrd), .B(fp_src2_in[50]), .Z(N803) );
  GTECH_AND2 C1361 ( .A(inq_fwrd_inv), .B(N806), .Z(N807) );
  GTECH_OR2 C1362 ( .A(N804), .B(N805), .Z(N806) );
  GTECH_AND2 C1363 ( .A(inq_bp), .B(inq_din_d1[50]), .Z(N804) );
  GTECH_AND2 C1364 ( .A(inq_bp_inv), .B(inq_dout[50]), .Z(N805) );
  GTECH_OR2 C1365 ( .A(N808), .B(N812), .Z(inq_in2[49]) );
  GTECH_AND2 C1366 ( .A(inq_fwrd), .B(fp_src2_in[49]), .Z(N808) );
  GTECH_AND2 C1367 ( .A(inq_fwrd_inv), .B(N811), .Z(N812) );
  GTECH_OR2 C1368 ( .A(N809), .B(N810), .Z(N811) );
  GTECH_AND2 C1369 ( .A(inq_bp), .B(inq_din_d1[49]), .Z(N809) );
  GTECH_AND2 C1370 ( .A(inq_bp_inv), .B(inq_dout[49]), .Z(N810) );
  GTECH_OR2 C1371 ( .A(N813), .B(N817), .Z(inq_in2[48]) );
  GTECH_AND2 C1372 ( .A(inq_fwrd), .B(fp_src2_in[48]), .Z(N813) );
  GTECH_AND2 C1373 ( .A(inq_fwrd_inv), .B(N816), .Z(N817) );
  GTECH_OR2 C1374 ( .A(N814), .B(N815), .Z(N816) );
  GTECH_AND2 C1375 ( .A(inq_bp), .B(inq_din_d1[48]), .Z(N814) );
  GTECH_AND2 C1376 ( .A(inq_bp_inv), .B(inq_dout[48]), .Z(N815) );
  GTECH_OR2 C1377 ( .A(N818), .B(N822), .Z(inq_in2[47]) );
  GTECH_AND2 C1378 ( .A(inq_fwrd), .B(fp_src2_in[47]), .Z(N818) );
  GTECH_AND2 C1379 ( .A(inq_fwrd_inv), .B(N821), .Z(N822) );
  GTECH_OR2 C1380 ( .A(N819), .B(N820), .Z(N821) );
  GTECH_AND2 C1381 ( .A(inq_bp), .B(inq_din_d1[47]), .Z(N819) );
  GTECH_AND2 C1382 ( .A(inq_bp_inv), .B(inq_dout[47]), .Z(N820) );
  GTECH_OR2 C1383 ( .A(N823), .B(N827), .Z(inq_in2[46]) );
  GTECH_AND2 C1384 ( .A(inq_fwrd), .B(fp_src2_in[46]), .Z(N823) );
  GTECH_AND2 C1385 ( .A(inq_fwrd_inv), .B(N826), .Z(N827) );
  GTECH_OR2 C1386 ( .A(N824), .B(N825), .Z(N826) );
  GTECH_AND2 C1387 ( .A(inq_bp), .B(inq_din_d1[46]), .Z(N824) );
  GTECH_AND2 C1388 ( .A(inq_bp_inv), .B(inq_dout[46]), .Z(N825) );
  GTECH_OR2 C1389 ( .A(N828), .B(N832), .Z(inq_in2[45]) );
  GTECH_AND2 C1390 ( .A(inq_fwrd), .B(fp_src2_in[45]), .Z(N828) );
  GTECH_AND2 C1391 ( .A(inq_fwrd_inv), .B(N831), .Z(N832) );
  GTECH_OR2 C1392 ( .A(N829), .B(N830), .Z(N831) );
  GTECH_AND2 C1393 ( .A(inq_bp), .B(inq_din_d1[45]), .Z(N829) );
  GTECH_AND2 C1394 ( .A(inq_bp_inv), .B(inq_dout[45]), .Z(N830) );
  GTECH_OR2 C1395 ( .A(N833), .B(N837), .Z(inq_in2[44]) );
  GTECH_AND2 C1396 ( .A(inq_fwrd), .B(fp_src2_in[44]), .Z(N833) );
  GTECH_AND2 C1397 ( .A(inq_fwrd_inv), .B(N836), .Z(N837) );
  GTECH_OR2 C1398 ( .A(N834), .B(N835), .Z(N836) );
  GTECH_AND2 C1399 ( .A(inq_bp), .B(inq_din_d1[44]), .Z(N834) );
  GTECH_AND2 C1400 ( .A(inq_bp_inv), .B(inq_dout[44]), .Z(N835) );
  GTECH_OR2 C1401 ( .A(N838), .B(N842), .Z(inq_in2[43]) );
  GTECH_AND2 C1402 ( .A(inq_fwrd), .B(fp_src2_in[43]), .Z(N838) );
  GTECH_AND2 C1403 ( .A(inq_fwrd_inv), .B(N841), .Z(N842) );
  GTECH_OR2 C1404 ( .A(N839), .B(N840), .Z(N841) );
  GTECH_AND2 C1405 ( .A(inq_bp), .B(inq_din_d1[43]), .Z(N839) );
  GTECH_AND2 C1406 ( .A(inq_bp_inv), .B(inq_dout[43]), .Z(N840) );
  GTECH_OR2 C1407 ( .A(N843), .B(N847), .Z(inq_in2[42]) );
  GTECH_AND2 C1408 ( .A(inq_fwrd), .B(fp_src2_in[42]), .Z(N843) );
  GTECH_AND2 C1409 ( .A(inq_fwrd_inv), .B(N846), .Z(N847) );
  GTECH_OR2 C1410 ( .A(N844), .B(N845), .Z(N846) );
  GTECH_AND2 C1411 ( .A(inq_bp), .B(inq_din_d1[42]), .Z(N844) );
  GTECH_AND2 C1412 ( .A(inq_bp_inv), .B(inq_dout[42]), .Z(N845) );
  GTECH_OR2 C1413 ( .A(N848), .B(N852), .Z(inq_in2[41]) );
  GTECH_AND2 C1414 ( .A(inq_fwrd), .B(fp_src2_in[41]), .Z(N848) );
  GTECH_AND2 C1415 ( .A(inq_fwrd_inv), .B(N851), .Z(N852) );
  GTECH_OR2 C1416 ( .A(N849), .B(N850), .Z(N851) );
  GTECH_AND2 C1417 ( .A(inq_bp), .B(inq_din_d1[41]), .Z(N849) );
  GTECH_AND2 C1418 ( .A(inq_bp_inv), .B(inq_dout[41]), .Z(N850) );
  GTECH_OR2 C1419 ( .A(N853), .B(N857), .Z(inq_in2[40]) );
  GTECH_AND2 C1420 ( .A(inq_fwrd), .B(fp_src2_in[40]), .Z(N853) );
  GTECH_AND2 C1421 ( .A(inq_fwrd_inv), .B(N856), .Z(N857) );
  GTECH_OR2 C1422 ( .A(N854), .B(N855), .Z(N856) );
  GTECH_AND2 C1423 ( .A(inq_bp), .B(inq_din_d1[40]), .Z(N854) );
  GTECH_AND2 C1424 ( .A(inq_bp_inv), .B(inq_dout[40]), .Z(N855) );
  GTECH_OR2 C1425 ( .A(N858), .B(N862), .Z(inq_in2[39]) );
  GTECH_AND2 C1426 ( .A(inq_fwrd), .B(fp_src2_in[39]), .Z(N858) );
  GTECH_AND2 C1427 ( .A(inq_fwrd_inv), .B(N861), .Z(N862) );
  GTECH_OR2 C1428 ( .A(N859), .B(N860), .Z(N861) );
  GTECH_AND2 C1429 ( .A(inq_bp), .B(inq_din_d1[39]), .Z(N859) );
  GTECH_AND2 C1430 ( .A(inq_bp_inv), .B(inq_dout[39]), .Z(N860) );
  GTECH_OR2 C1431 ( .A(N863), .B(N867), .Z(inq_in2[38]) );
  GTECH_AND2 C1432 ( .A(inq_fwrd), .B(fp_src2_in[38]), .Z(N863) );
  GTECH_AND2 C1433 ( .A(inq_fwrd_inv), .B(N866), .Z(N867) );
  GTECH_OR2 C1434 ( .A(N864), .B(N865), .Z(N866) );
  GTECH_AND2 C1435 ( .A(inq_bp), .B(inq_din_d1[38]), .Z(N864) );
  GTECH_AND2 C1436 ( .A(inq_bp_inv), .B(inq_dout[38]), .Z(N865) );
  GTECH_OR2 C1437 ( .A(N868), .B(N872), .Z(inq_in2[37]) );
  GTECH_AND2 C1438 ( .A(inq_fwrd), .B(fp_src2_in[37]), .Z(N868) );
  GTECH_AND2 C1439 ( .A(inq_fwrd_inv), .B(N871), .Z(N872) );
  GTECH_OR2 C1440 ( .A(N869), .B(N870), .Z(N871) );
  GTECH_AND2 C1441 ( .A(inq_bp), .B(inq_din_d1[37]), .Z(N869) );
  GTECH_AND2 C1442 ( .A(inq_bp_inv), .B(inq_dout[37]), .Z(N870) );
  GTECH_OR2 C1443 ( .A(N873), .B(N877), .Z(inq_in2[36]) );
  GTECH_AND2 C1444 ( .A(inq_fwrd), .B(fp_src2_in[36]), .Z(N873) );
  GTECH_AND2 C1445 ( .A(inq_fwrd_inv), .B(N876), .Z(N877) );
  GTECH_OR2 C1446 ( .A(N874), .B(N875), .Z(N876) );
  GTECH_AND2 C1447 ( .A(inq_bp), .B(inq_din_d1[36]), .Z(N874) );
  GTECH_AND2 C1448 ( .A(inq_bp_inv), .B(inq_dout[36]), .Z(N875) );
  GTECH_OR2 C1449 ( .A(N878), .B(N882), .Z(inq_in2[35]) );
  GTECH_AND2 C1450 ( .A(inq_fwrd), .B(fp_src2_in[35]), .Z(N878) );
  GTECH_AND2 C1451 ( .A(inq_fwrd_inv), .B(N881), .Z(N882) );
  GTECH_OR2 C1452 ( .A(N879), .B(N880), .Z(N881) );
  GTECH_AND2 C1453 ( .A(inq_bp), .B(inq_din_d1[35]), .Z(N879) );
  GTECH_AND2 C1454 ( .A(inq_bp_inv), .B(inq_dout[35]), .Z(N880) );
  GTECH_OR2 C1455 ( .A(N883), .B(N887), .Z(inq_in2[34]) );
  GTECH_AND2 C1456 ( .A(inq_fwrd), .B(fp_src2_in[34]), .Z(N883) );
  GTECH_AND2 C1457 ( .A(inq_fwrd_inv), .B(N886), .Z(N887) );
  GTECH_OR2 C1458 ( .A(N884), .B(N885), .Z(N886) );
  GTECH_AND2 C1459 ( .A(inq_bp), .B(inq_din_d1[34]), .Z(N884) );
  GTECH_AND2 C1460 ( .A(inq_bp_inv), .B(inq_dout[34]), .Z(N885) );
  GTECH_OR2 C1461 ( .A(N888), .B(N892), .Z(inq_in2[33]) );
  GTECH_AND2 C1462 ( .A(inq_fwrd), .B(fp_src2_in[33]), .Z(N888) );
  GTECH_AND2 C1463 ( .A(inq_fwrd_inv), .B(N891), .Z(N892) );
  GTECH_OR2 C1464 ( .A(N889), .B(N890), .Z(N891) );
  GTECH_AND2 C1465 ( .A(inq_bp), .B(inq_din_d1[33]), .Z(N889) );
  GTECH_AND2 C1466 ( .A(inq_bp_inv), .B(inq_dout[33]), .Z(N890) );
  GTECH_OR2 C1467 ( .A(N893), .B(N897), .Z(inq_in2[32]) );
  GTECH_AND2 C1468 ( .A(inq_fwrd), .B(fp_src2_in[32]), .Z(N893) );
  GTECH_AND2 C1469 ( .A(inq_fwrd_inv), .B(N896), .Z(N897) );
  GTECH_OR2 C1470 ( .A(N894), .B(N895), .Z(N896) );
  GTECH_AND2 C1471 ( .A(inq_bp), .B(inq_din_d1[32]), .Z(N894) );
  GTECH_AND2 C1472 ( .A(inq_bp_inv), .B(inq_dout[32]), .Z(N895) );
  GTECH_OR2 C1473 ( .A(N898), .B(N902), .Z(inq_in2[31]) );
  GTECH_AND2 C1474 ( .A(inq_fwrd), .B(fp_src2_in[31]), .Z(N898) );
  GTECH_AND2 C1475 ( .A(inq_fwrd_inv), .B(N901), .Z(N902) );
  GTECH_OR2 C1476 ( .A(N899), .B(N900), .Z(N901) );
  GTECH_AND2 C1477 ( .A(inq_bp), .B(inq_din_d1[31]), .Z(N899) );
  GTECH_AND2 C1478 ( .A(inq_bp_inv), .B(inq_dout[31]), .Z(N900) );
  GTECH_OR2 C1479 ( .A(N903), .B(N907), .Z(inq_in2[30]) );
  GTECH_AND2 C1480 ( .A(inq_fwrd), .B(fp_src2_in[30]), .Z(N903) );
  GTECH_AND2 C1481 ( .A(inq_fwrd_inv), .B(N906), .Z(N907) );
  GTECH_OR2 C1482 ( .A(N904), .B(N905), .Z(N906) );
  GTECH_AND2 C1483 ( .A(inq_bp), .B(inq_din_d1[30]), .Z(N904) );
  GTECH_AND2 C1484 ( .A(inq_bp_inv), .B(inq_dout[30]), .Z(N905) );
  GTECH_OR2 C1485 ( .A(N908), .B(N912), .Z(inq_in2[29]) );
  GTECH_AND2 C1486 ( .A(inq_fwrd), .B(fp_src2_in[29]), .Z(N908) );
  GTECH_AND2 C1487 ( .A(inq_fwrd_inv), .B(N911), .Z(N912) );
  GTECH_OR2 C1488 ( .A(N909), .B(N910), .Z(N911) );
  GTECH_AND2 C1489 ( .A(inq_bp), .B(inq_din_d1[29]), .Z(N909) );
  GTECH_AND2 C1490 ( .A(inq_bp_inv), .B(inq_dout[29]), .Z(N910) );
  GTECH_OR2 C1491 ( .A(N913), .B(N917), .Z(inq_in2[28]) );
  GTECH_AND2 C1492 ( .A(inq_fwrd), .B(fp_src2_in[28]), .Z(N913) );
  GTECH_AND2 C1493 ( .A(inq_fwrd_inv), .B(N916), .Z(N917) );
  GTECH_OR2 C1494 ( .A(N914), .B(N915), .Z(N916) );
  GTECH_AND2 C1495 ( .A(inq_bp), .B(inq_din_d1[28]), .Z(N914) );
  GTECH_AND2 C1496 ( .A(inq_bp_inv), .B(inq_dout[28]), .Z(N915) );
  GTECH_OR2 C1497 ( .A(N918), .B(N922), .Z(inq_in2[27]) );
  GTECH_AND2 C1498 ( .A(inq_fwrd), .B(fp_src2_in[27]), .Z(N918) );
  GTECH_AND2 C1499 ( .A(inq_fwrd_inv), .B(N921), .Z(N922) );
  GTECH_OR2 C1500 ( .A(N919), .B(N920), .Z(N921) );
  GTECH_AND2 C1501 ( .A(inq_bp), .B(inq_din_d1[27]), .Z(N919) );
  GTECH_AND2 C1502 ( .A(inq_bp_inv), .B(inq_dout[27]), .Z(N920) );
  GTECH_OR2 C1503 ( .A(N923), .B(N927), .Z(inq_in2[26]) );
  GTECH_AND2 C1504 ( .A(inq_fwrd), .B(fp_src2_in[26]), .Z(N923) );
  GTECH_AND2 C1505 ( .A(inq_fwrd_inv), .B(N926), .Z(N927) );
  GTECH_OR2 C1506 ( .A(N924), .B(N925), .Z(N926) );
  GTECH_AND2 C1507 ( .A(inq_bp), .B(inq_din_d1[26]), .Z(N924) );
  GTECH_AND2 C1508 ( .A(inq_bp_inv), .B(inq_dout[26]), .Z(N925) );
  GTECH_OR2 C1509 ( .A(N928), .B(N932), .Z(inq_in2[25]) );
  GTECH_AND2 C1510 ( .A(inq_fwrd), .B(fp_src2_in[25]), .Z(N928) );
  GTECH_AND2 C1511 ( .A(inq_fwrd_inv), .B(N931), .Z(N932) );
  GTECH_OR2 C1512 ( .A(N929), .B(N930), .Z(N931) );
  GTECH_AND2 C1513 ( .A(inq_bp), .B(inq_din_d1[25]), .Z(N929) );
  GTECH_AND2 C1514 ( .A(inq_bp_inv), .B(inq_dout[25]), .Z(N930) );
  GTECH_OR2 C1515 ( .A(N933), .B(N937), .Z(inq_in2[24]) );
  GTECH_AND2 C1516 ( .A(inq_fwrd), .B(fp_src2_in[24]), .Z(N933) );
  GTECH_AND2 C1517 ( .A(inq_fwrd_inv), .B(N936), .Z(N937) );
  GTECH_OR2 C1518 ( .A(N934), .B(N935), .Z(N936) );
  GTECH_AND2 C1519 ( .A(inq_bp), .B(inq_din_d1[24]), .Z(N934) );
  GTECH_AND2 C1520 ( .A(inq_bp_inv), .B(inq_dout[24]), .Z(N935) );
  GTECH_OR2 C1521 ( .A(N938), .B(N942), .Z(inq_in2[23]) );
  GTECH_AND2 C1522 ( .A(inq_fwrd), .B(fp_src2_in[23]), .Z(N938) );
  GTECH_AND2 C1523 ( .A(inq_fwrd_inv), .B(N941), .Z(N942) );
  GTECH_OR2 C1524 ( .A(N939), .B(N940), .Z(N941) );
  GTECH_AND2 C1525 ( .A(inq_bp), .B(inq_din_d1[23]), .Z(N939) );
  GTECH_AND2 C1526 ( .A(inq_bp_inv), .B(inq_dout[23]), .Z(N940) );
  GTECH_OR2 C1527 ( .A(N943), .B(N947), .Z(inq_in2[22]) );
  GTECH_AND2 C1528 ( .A(inq_fwrd), .B(fp_src2_in[22]), .Z(N943) );
  GTECH_AND2 C1529 ( .A(inq_fwrd_inv), .B(N946), .Z(N947) );
  GTECH_OR2 C1530 ( .A(N944), .B(N945), .Z(N946) );
  GTECH_AND2 C1531 ( .A(inq_bp), .B(inq_din_d1[22]), .Z(N944) );
  GTECH_AND2 C1532 ( .A(inq_bp_inv), .B(inq_dout[22]), .Z(N945) );
  GTECH_OR2 C1533 ( .A(N948), .B(N952), .Z(inq_in2[21]) );
  GTECH_AND2 C1534 ( .A(inq_fwrd), .B(fp_src2_in[21]), .Z(N948) );
  GTECH_AND2 C1535 ( .A(inq_fwrd_inv), .B(N951), .Z(N952) );
  GTECH_OR2 C1536 ( .A(N949), .B(N950), .Z(N951) );
  GTECH_AND2 C1537 ( .A(inq_bp), .B(inq_din_d1[21]), .Z(N949) );
  GTECH_AND2 C1538 ( .A(inq_bp_inv), .B(inq_dout[21]), .Z(N950) );
  GTECH_OR2 C1539 ( .A(N953), .B(N957), .Z(inq_in2[20]) );
  GTECH_AND2 C1540 ( .A(inq_fwrd), .B(fp_src2_in[20]), .Z(N953) );
  GTECH_AND2 C1541 ( .A(inq_fwrd_inv), .B(N956), .Z(N957) );
  GTECH_OR2 C1542 ( .A(N954), .B(N955), .Z(N956) );
  GTECH_AND2 C1543 ( .A(inq_bp), .B(inq_din_d1[20]), .Z(N954) );
  GTECH_AND2 C1544 ( .A(inq_bp_inv), .B(inq_dout[20]), .Z(N955) );
  GTECH_OR2 C1545 ( .A(N958), .B(N962), .Z(inq_in2[19]) );
  GTECH_AND2 C1546 ( .A(inq_fwrd), .B(fp_src2_in[19]), .Z(N958) );
  GTECH_AND2 C1547 ( .A(inq_fwrd_inv), .B(N961), .Z(N962) );
  GTECH_OR2 C1548 ( .A(N959), .B(N960), .Z(N961) );
  GTECH_AND2 C1549 ( .A(inq_bp), .B(inq_din_d1[19]), .Z(N959) );
  GTECH_AND2 C1550 ( .A(inq_bp_inv), .B(inq_dout[19]), .Z(N960) );
  GTECH_OR2 C1551 ( .A(N963), .B(N967), .Z(inq_in2[18]) );
  GTECH_AND2 C1552 ( .A(inq_fwrd), .B(fp_src2_in[18]), .Z(N963) );
  GTECH_AND2 C1553 ( .A(inq_fwrd_inv), .B(N966), .Z(N967) );
  GTECH_OR2 C1554 ( .A(N964), .B(N965), .Z(N966) );
  GTECH_AND2 C1555 ( .A(inq_bp), .B(inq_din_d1[18]), .Z(N964) );
  GTECH_AND2 C1556 ( .A(inq_bp_inv), .B(inq_dout[18]), .Z(N965) );
  GTECH_OR2 C1557 ( .A(N968), .B(N972), .Z(inq_in2[17]) );
  GTECH_AND2 C1558 ( .A(inq_fwrd), .B(fp_src2_in[17]), .Z(N968) );
  GTECH_AND2 C1559 ( .A(inq_fwrd_inv), .B(N971), .Z(N972) );
  GTECH_OR2 C1560 ( .A(N969), .B(N970), .Z(N971) );
  GTECH_AND2 C1561 ( .A(inq_bp), .B(inq_din_d1[17]), .Z(N969) );
  GTECH_AND2 C1562 ( .A(inq_bp_inv), .B(inq_dout[17]), .Z(N970) );
  GTECH_OR2 C1563 ( .A(N973), .B(N977), .Z(inq_in2[16]) );
  GTECH_AND2 C1564 ( .A(inq_fwrd), .B(fp_src2_in[16]), .Z(N973) );
  GTECH_AND2 C1565 ( .A(inq_fwrd_inv), .B(N976), .Z(N977) );
  GTECH_OR2 C1566 ( .A(N974), .B(N975), .Z(N976) );
  GTECH_AND2 C1567 ( .A(inq_bp), .B(inq_din_d1[16]), .Z(N974) );
  GTECH_AND2 C1568 ( .A(inq_bp_inv), .B(inq_dout[16]), .Z(N975) );
  GTECH_OR2 C1569 ( .A(N978), .B(N982), .Z(inq_in2[15]) );
  GTECH_AND2 C1570 ( .A(inq_fwrd), .B(fp_src2_in[15]), .Z(N978) );
  GTECH_AND2 C1571 ( .A(inq_fwrd_inv), .B(N981), .Z(N982) );
  GTECH_OR2 C1572 ( .A(N979), .B(N980), .Z(N981) );
  GTECH_AND2 C1573 ( .A(inq_bp), .B(inq_din_d1[15]), .Z(N979) );
  GTECH_AND2 C1574 ( .A(inq_bp_inv), .B(inq_dout[15]), .Z(N980) );
  GTECH_OR2 C1575 ( .A(N983), .B(N987), .Z(inq_in2[14]) );
  GTECH_AND2 C1576 ( .A(inq_fwrd), .B(fp_src2_in[14]), .Z(N983) );
  GTECH_AND2 C1577 ( .A(inq_fwrd_inv), .B(N986), .Z(N987) );
  GTECH_OR2 C1578 ( .A(N984), .B(N985), .Z(N986) );
  GTECH_AND2 C1579 ( .A(inq_bp), .B(inq_din_d1[14]), .Z(N984) );
  GTECH_AND2 C1580 ( .A(inq_bp_inv), .B(inq_dout[14]), .Z(N985) );
  GTECH_OR2 C1581 ( .A(N988), .B(N992), .Z(inq_in2[13]) );
  GTECH_AND2 C1582 ( .A(inq_fwrd), .B(fp_src2_in[13]), .Z(N988) );
  GTECH_AND2 C1583 ( .A(inq_fwrd_inv), .B(N991), .Z(N992) );
  GTECH_OR2 C1584 ( .A(N989), .B(N990), .Z(N991) );
  GTECH_AND2 C1585 ( .A(inq_bp), .B(inq_din_d1[13]), .Z(N989) );
  GTECH_AND2 C1586 ( .A(inq_bp_inv), .B(inq_dout[13]), .Z(N990) );
  GTECH_OR2 C1587 ( .A(N993), .B(N997), .Z(inq_in2[12]) );
  GTECH_AND2 C1588 ( .A(inq_fwrd), .B(fp_src2_in[12]), .Z(N993) );
  GTECH_AND2 C1589 ( .A(inq_fwrd_inv), .B(N996), .Z(N997) );
  GTECH_OR2 C1590 ( .A(N994), .B(N995), .Z(N996) );
  GTECH_AND2 C1591 ( .A(inq_bp), .B(inq_din_d1[12]), .Z(N994) );
  GTECH_AND2 C1592 ( .A(inq_bp_inv), .B(inq_dout[12]), .Z(N995) );
  GTECH_OR2 C1593 ( .A(N998), .B(N1002), .Z(inq_in2[11]) );
  GTECH_AND2 C1594 ( .A(inq_fwrd), .B(fp_src2_in[11]), .Z(N998) );
  GTECH_AND2 C1595 ( .A(inq_fwrd_inv), .B(N1001), .Z(N1002) );
  GTECH_OR2 C1596 ( .A(N999), .B(N1000), .Z(N1001) );
  GTECH_AND2 C1597 ( .A(inq_bp), .B(inq_din_d1[11]), .Z(N999) );
  GTECH_AND2 C1598 ( .A(inq_bp_inv), .B(inq_dout[11]), .Z(N1000) );
  GTECH_OR2 C1599 ( .A(N1003), .B(N1007), .Z(inq_in2[10]) );
  GTECH_AND2 C1600 ( .A(inq_fwrd), .B(fp_src2_in[10]), .Z(N1003) );
  GTECH_AND2 C1601 ( .A(inq_fwrd_inv), .B(N1006), .Z(N1007) );
  GTECH_OR2 C1602 ( .A(N1004), .B(N1005), .Z(N1006) );
  GTECH_AND2 C1603 ( .A(inq_bp), .B(inq_din_d1[10]), .Z(N1004) );
  GTECH_AND2 C1604 ( .A(inq_bp_inv), .B(inq_dout[10]), .Z(N1005) );
  GTECH_OR2 C1605 ( .A(N1008), .B(N1012), .Z(inq_in2[9]) );
  GTECH_AND2 C1606 ( .A(inq_fwrd), .B(fp_src2_in[9]), .Z(N1008) );
  GTECH_AND2 C1607 ( .A(inq_fwrd_inv), .B(N1011), .Z(N1012) );
  GTECH_OR2 C1608 ( .A(N1009), .B(N1010), .Z(N1011) );
  GTECH_AND2 C1609 ( .A(inq_bp), .B(inq_din_d1[9]), .Z(N1009) );
  GTECH_AND2 C1610 ( .A(inq_bp_inv), .B(inq_dout[9]), .Z(N1010) );
  GTECH_OR2 C1611 ( .A(N1013), .B(N1017), .Z(inq_in2[8]) );
  GTECH_AND2 C1612 ( .A(inq_fwrd), .B(fp_src2_in[8]), .Z(N1013) );
  GTECH_AND2 C1613 ( .A(inq_fwrd_inv), .B(N1016), .Z(N1017) );
  GTECH_OR2 C1614 ( .A(N1014), .B(N1015), .Z(N1016) );
  GTECH_AND2 C1615 ( .A(inq_bp), .B(inq_din_d1[8]), .Z(N1014) );
  GTECH_AND2 C1616 ( .A(inq_bp_inv), .B(inq_dout[8]), .Z(N1015) );
  GTECH_OR2 C1617 ( .A(N1018), .B(N1022), .Z(inq_in2[7]) );
  GTECH_AND2 C1618 ( .A(inq_fwrd), .B(fp_src2_in[7]), .Z(N1018) );
  GTECH_AND2 C1619 ( .A(inq_fwrd_inv), .B(N1021), .Z(N1022) );
  GTECH_OR2 C1620 ( .A(N1019), .B(N1020), .Z(N1021) );
  GTECH_AND2 C1621 ( .A(inq_bp), .B(inq_din_d1[7]), .Z(N1019) );
  GTECH_AND2 C1622 ( .A(inq_bp_inv), .B(inq_dout[7]), .Z(N1020) );
  GTECH_OR2 C1623 ( .A(N1023), .B(N1027), .Z(inq_in2[6]) );
  GTECH_AND2 C1624 ( .A(inq_fwrd), .B(fp_src2_in[6]), .Z(N1023) );
  GTECH_AND2 C1625 ( .A(inq_fwrd_inv), .B(N1026), .Z(N1027) );
  GTECH_OR2 C1626 ( .A(N1024), .B(N1025), .Z(N1026) );
  GTECH_AND2 C1627 ( .A(inq_bp), .B(inq_din_d1[6]), .Z(N1024) );
  GTECH_AND2 C1628 ( .A(inq_bp_inv), .B(inq_dout[6]), .Z(N1025) );
  GTECH_OR2 C1629 ( .A(N1028), .B(N1032), .Z(inq_in2[5]) );
  GTECH_AND2 C1630 ( .A(inq_fwrd), .B(fp_src2_in[5]), .Z(N1028) );
  GTECH_AND2 C1631 ( .A(inq_fwrd_inv), .B(N1031), .Z(N1032) );
  GTECH_OR2 C1632 ( .A(N1029), .B(N1030), .Z(N1031) );
  GTECH_AND2 C1633 ( .A(inq_bp), .B(inq_din_d1[5]), .Z(N1029) );
  GTECH_AND2 C1634 ( .A(inq_bp_inv), .B(inq_dout[5]), .Z(N1030) );
  GTECH_OR2 C1635 ( .A(N1033), .B(N1037), .Z(inq_in2[4]) );
  GTECH_AND2 C1636 ( .A(inq_fwrd), .B(fp_src2_in[4]), .Z(N1033) );
  GTECH_AND2 C1637 ( .A(inq_fwrd_inv), .B(N1036), .Z(N1037) );
  GTECH_OR2 C1638 ( .A(N1034), .B(N1035), .Z(N1036) );
  GTECH_AND2 C1639 ( .A(inq_bp), .B(inq_din_d1[4]), .Z(N1034) );
  GTECH_AND2 C1640 ( .A(inq_bp_inv), .B(inq_dout[4]), .Z(N1035) );
  GTECH_OR2 C1641 ( .A(N1038), .B(N1042), .Z(inq_in2[3]) );
  GTECH_AND2 C1642 ( .A(inq_fwrd), .B(fp_src2_in[3]), .Z(N1038) );
  GTECH_AND2 C1643 ( .A(inq_fwrd_inv), .B(N1041), .Z(N1042) );
  GTECH_OR2 C1644 ( .A(N1039), .B(N1040), .Z(N1041) );
  GTECH_AND2 C1645 ( .A(inq_bp), .B(inq_din_d1[3]), .Z(N1039) );
  GTECH_AND2 C1646 ( .A(inq_bp_inv), .B(inq_dout[3]), .Z(N1040) );
  GTECH_OR2 C1647 ( .A(N1043), .B(N1047), .Z(inq_in2[2]) );
  GTECH_AND2 C1648 ( .A(inq_fwrd), .B(fp_src2_in[2]), .Z(N1043) );
  GTECH_AND2 C1649 ( .A(inq_fwrd_inv), .B(N1046), .Z(N1047) );
  GTECH_OR2 C1650 ( .A(N1044), .B(N1045), .Z(N1046) );
  GTECH_AND2 C1651 ( .A(inq_bp), .B(inq_din_d1[2]), .Z(N1044) );
  GTECH_AND2 C1652 ( .A(inq_bp_inv), .B(inq_dout[2]), .Z(N1045) );
  GTECH_OR2 C1653 ( .A(N1048), .B(N1052), .Z(inq_in2[1]) );
  GTECH_AND2 C1654 ( .A(inq_fwrd), .B(fp_src2_in[1]), .Z(N1048) );
  GTECH_AND2 C1655 ( .A(inq_fwrd_inv), .B(N1051), .Z(N1052) );
  GTECH_OR2 C1656 ( .A(N1049), .B(N1050), .Z(N1051) );
  GTECH_AND2 C1657 ( .A(inq_bp), .B(inq_din_d1[1]), .Z(N1049) );
  GTECH_AND2 C1658 ( .A(inq_bp_inv), .B(inq_dout[1]), .Z(N1050) );
  GTECH_OR2 C1659 ( .A(N1053), .B(N1057), .Z(inq_in2[0]) );
  GTECH_AND2 C1660 ( .A(inq_fwrd), .B(fp_src2_in[0]), .Z(N1053) );
  GTECH_AND2 C1661 ( .A(inq_fwrd_inv), .B(N1056), .Z(N1057) );
  GTECH_OR2 C1662 ( .A(N1054), .B(N1055), .Z(N1056) );
  GTECH_AND2 C1663 ( .A(inq_bp), .B(inq_din_d1[0]), .Z(N1054) );
  GTECH_AND2 C1664 ( .A(inq_bp_inv), .B(inq_dout[0]), .Z(N1055) );
endmodule


module fpu_in ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, a1stg_step, 
        m1stg_step, d1stg_step, add_pipe_active, mul_pipe_active, 
        div_pipe_active, inq_dout, sehold, arst_l, grst_l, rclk, fadd_clken_l, 
        fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div, inq_id, 
        inq_rnd_mode, inq_fcc, inq_op, inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, 
        inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1, 
        inq_in2_exp_neq_ffs, inq_in2_exp_eq_0, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2, fp_id_in, 
        fp_rnd_mode_in, fp_fcc_in, fp_op_in, fp_src1_in, fp_src2_in, 
        inq_rdaddr, inq_wraddr, inq_read_en, inq_we, se, si, so );
  input [123:0] pcx_fpio_data_px2;
  input [154:0] inq_dout;
  output [4:0] inq_id;
  output [1:0] inq_rnd_mode;
  output [1:0] inq_fcc;
  output [7:0] inq_op;
  output [63:0] inq_in1;
  output [63:0] inq_in2;
  output [4:0] fp_id_in;
  output [1:0] fp_rnd_mode_in;
  output [1:0] fp_fcc_in;
  output [7:0] fp_op_in;
  output [68:0] fp_src1_in;
  output [68:0] fp_src2_in;
  output [3:0] inq_rdaddr;
  output [3:0] inq_wraddr;
  input pcx_fpio_data_rdy_px2, a1stg_step, m1stg_step, d1stg_step,
         add_pipe_active, mul_pipe_active, div_pipe_active, sehold, arst_l,
         grst_l, rclk, se, si;
  output fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div,
         inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, inq_in1_53_0_neq_0,
         inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in2_exp_neq_ffs,
         inq_in2_exp_eq_0, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_read_en, inq_we, so;
  wire   pcx_fpio_data_px2_123, pcx_fpio_data_px2_122, pcx_fpio_data_px2_121,
         pcx_fpio_data_px2_120, pcx_fpio_data_px2_119, pcx_fpio_data_px2_118,
         pcx_fpio_data_px2_116, pcx_fpio_data_px2_115, pcx_fpio_data_px2_114,
         pcx_fpio_data_px2_113, pcx_fpio_data_px2_112, pcx_fpio_data_px2_79,
         pcx_fpio_data_px2_78, pcx_fpio_data_px2_77, pcx_fpio_data_px2_76,
         pcx_fpio_data_px2_75, pcx_fpio_data_px2_74, pcx_fpio_data_px2_73,
         pcx_fpio_data_px2_72, fp_op_in_7in, fp_data_rdy, inq_bp, inq_bp_inv,
         inq_fwrd, inq_fwrd_inv, scan_out_fpu_in_ctl;
  assign pcx_fpio_data_px2_123 = pcx_fpio_data_px2[123];
  assign pcx_fpio_data_px2_122 = pcx_fpio_data_px2[122];
  assign pcx_fpio_data_px2_121 = pcx_fpio_data_px2[121];
  assign pcx_fpio_data_px2_120 = pcx_fpio_data_px2[120];
  assign pcx_fpio_data_px2_119 = pcx_fpio_data_px2[119];
  assign pcx_fpio_data_px2_118 = pcx_fpio_data_px2[118];
  assign pcx_fpio_data_px2_116 = pcx_fpio_data_px2[116];
  assign pcx_fpio_data_px2_115 = pcx_fpio_data_px2[115];
  assign pcx_fpio_data_px2_114 = pcx_fpio_data_px2[114];
  assign pcx_fpio_data_px2_113 = pcx_fpio_data_px2[113];
  assign pcx_fpio_data_px2_112 = pcx_fpio_data_px2[112];
  assign pcx_fpio_data_px2_79 = pcx_fpio_data_px2[79];
  assign pcx_fpio_data_px2_78 = pcx_fpio_data_px2[78];
  assign pcx_fpio_data_px2_77 = pcx_fpio_data_px2[77];
  assign pcx_fpio_data_px2_76 = pcx_fpio_data_px2[76];
  assign pcx_fpio_data_px2_75 = pcx_fpio_data_px2[75];
  assign pcx_fpio_data_px2_74 = pcx_fpio_data_px2[74];
  assign pcx_fpio_data_px2_73 = pcx_fpio_data_px2[73];
  assign pcx_fpio_data_px2_72 = pcx_fpio_data_px2[72];

  fpu_in_ctl fpu_in_ctl ( .pcx_fpio_data_rdy_px2(pcx_fpio_data_rdy_px2), 
        .pcx_fpio_data_px2({pcx_fpio_data_px2_123, pcx_fpio_data_px2_122, 
        pcx_fpio_data_px2_121, pcx_fpio_data_px2_120, pcx_fpio_data_px2_119, 
        pcx_fpio_data_px2_118}), .fp_op_in(fp_op_in[3:2]), .fp_op_in_7in(
        fp_op_in_7in), .a1stg_step(a1stg_step), .m1stg_step(m1stg_step), 
        .d1stg_step(d1stg_step), .add_pipe_active(add_pipe_active), 
        .mul_pipe_active(mul_pipe_active), .div_pipe_active(div_pipe_active), 
        .sehold(sehold), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), 
        .fp_data_rdy(fp_data_rdy), .fadd_clken_l(fadd_clken_l), .fmul_clken_l(
        fmul_clken_l), .fdiv_clken_l(fdiv_clken_l), .inq_we(inq_we), 
        .inq_wraddr(inq_wraddr), .inq_read_en(inq_read_en), .inq_rdaddr(
        inq_rdaddr), .inq_bp(inq_bp), .inq_bp_inv(inq_bp_inv), .inq_fwrd(
        inq_fwrd), .inq_fwrd_inv(inq_fwrd_inv), .inq_add(inq_add), .inq_mul(
        inq_mul), .inq_div(inq_div), .se(se), .si(si), .so(scan_out_fpu_in_ctl) );
  fpu_in_dp fpu_in_dp ( .fp_data_rdy(fp_data_rdy), .fpio_data_px2_116_112({
        pcx_fpio_data_px2_116, pcx_fpio_data_px2_115, pcx_fpio_data_px2_114, 
        pcx_fpio_data_px2_113, pcx_fpio_data_px2_112}), .fpio_data_px2_79_72({
        pcx_fpio_data_px2_79, pcx_fpio_data_px2_78, pcx_fpio_data_px2_77, 
        pcx_fpio_data_px2_76, pcx_fpio_data_px2_75, pcx_fpio_data_px2_74, 
        pcx_fpio_data_px2_73, pcx_fpio_data_px2_72}), .fpio_data_px2_67_0(
        pcx_fpio_data_px2[67:0]), .inq_fwrd(inq_fwrd), .inq_fwrd_inv(
        inq_fwrd_inv), .inq_bp(inq_bp), .inq_bp_inv(inq_bp_inv), .inq_dout(
        inq_dout), .rclk(rclk), .fp_op_in_7in(fp_op_in_7in), .inq_id(inq_id), 
        .inq_rnd_mode(inq_rnd_mode), .inq_fcc(inq_fcc), .inq_op(inq_op), 
        .inq_in1_exp_neq_ffs(inq_in1_exp_neq_ffs), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(
        inq_in1_53_32_neq_0), .inq_in1(inq_in1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), 
        .inq_in2(inq_in2), .fp_id_in(fp_id_in), .fp_rnd_mode_in(fp_rnd_mode_in), .fp_fcc_in(fp_fcc_in), .fp_op_in(fp_op_in), .fp_src1_in(fp_src1_in), 
        .fp_src2_in(fp_src2_in), .se(se), .si(scan_out_fpu_in_ctl), .so(so) );
endmodule


module bw_r_rf16x160 ( dout, so_w, so_r, din, rd_adr, wr_adr, read_en, wr_en, 
        rst_tri_en, word_wen, byte_wen, rd_clk, wr_clk, se, si_r, si_w, 
        reset_l, sehold );
  output [159:0] dout;
  input [159:0] din;
  input [3:0] rd_adr;
  input [3:0] wr_adr;
  input [3:0] word_wen;
  input [19:0] byte_wen;
  input read_en, wr_en, rst_tri_en, rd_clk, wr_clk, se, si_r, si_w, reset_l,
         sehold;
  output so_w, so_r;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         wr_en_d1, ren_d1, \inq_ary[15][159] , \inq_ary[15][158] ,
         \inq_ary[15][157] , \inq_ary[15][156] , \inq_ary[15][155] ,
         \inq_ary[15][154] , \inq_ary[15][153] , \inq_ary[15][152] ,
         \inq_ary[15][151] , \inq_ary[15][150] , \inq_ary[15][149] ,
         \inq_ary[15][148] , \inq_ary[15][147] , \inq_ary[15][146] ,
         \inq_ary[15][145] , \inq_ary[15][144] , \inq_ary[15][143] ,
         \inq_ary[15][142] , \inq_ary[15][141] , \inq_ary[15][140] ,
         \inq_ary[15][139] , \inq_ary[15][138] , \inq_ary[15][137] ,
         \inq_ary[15][136] , \inq_ary[15][135] , \inq_ary[15][134] ,
         \inq_ary[15][133] , \inq_ary[15][132] , \inq_ary[15][131] ,
         \inq_ary[15][130] , \inq_ary[15][129] , \inq_ary[15][128] ,
         \inq_ary[15][127] , \inq_ary[15][126] , \inq_ary[15][125] ,
         \inq_ary[15][124] , \inq_ary[15][123] , \inq_ary[15][122] ,
         \inq_ary[15][121] , \inq_ary[15][120] , \inq_ary[15][119] ,
         \inq_ary[15][118] , \inq_ary[15][117] , \inq_ary[15][116] ,
         \inq_ary[15][115] , \inq_ary[15][114] , \inq_ary[15][113] ,
         \inq_ary[15][112] , \inq_ary[15][111] , \inq_ary[15][110] ,
         \inq_ary[15][109] , \inq_ary[15][108] , \inq_ary[15][107] ,
         \inq_ary[15][106] , \inq_ary[15][105] , \inq_ary[15][104] ,
         \inq_ary[15][103] , \inq_ary[15][102] , \inq_ary[15][101] ,
         \inq_ary[15][100] , \inq_ary[15][99] , \inq_ary[15][98] ,
         \inq_ary[15][97] , \inq_ary[15][96] , \inq_ary[15][95] ,
         \inq_ary[15][94] , \inq_ary[15][93] , \inq_ary[15][92] ,
         \inq_ary[15][91] , \inq_ary[15][90] , \inq_ary[15][89] ,
         \inq_ary[15][88] , \inq_ary[15][87] , \inq_ary[15][86] ,
         \inq_ary[15][85] , \inq_ary[15][84] , \inq_ary[15][83] ,
         \inq_ary[15][82] , \inq_ary[15][81] , \inq_ary[15][80] ,
         \inq_ary[15][79] , \inq_ary[15][78] , \inq_ary[15][77] ,
         \inq_ary[15][76] , \inq_ary[15][75] , \inq_ary[15][74] ,
         \inq_ary[15][73] , \inq_ary[15][72] , \inq_ary[15][71] ,
         \inq_ary[15][70] , \inq_ary[15][69] , \inq_ary[15][68] ,
         \inq_ary[15][67] , \inq_ary[15][66] , \inq_ary[15][65] ,
         \inq_ary[15][64] , \inq_ary[15][63] , \inq_ary[15][62] ,
         \inq_ary[15][61] , \inq_ary[15][60] , \inq_ary[15][59] ,
         \inq_ary[15][58] , \inq_ary[15][57] , \inq_ary[15][56] ,
         \inq_ary[15][55] , \inq_ary[15][54] , \inq_ary[15][53] ,
         \inq_ary[15][52] , \inq_ary[15][51] , \inq_ary[15][50] ,
         \inq_ary[15][49] , \inq_ary[15][48] , \inq_ary[15][47] ,
         \inq_ary[15][46] , \inq_ary[15][45] , \inq_ary[15][44] ,
         \inq_ary[15][43] , \inq_ary[15][42] , \inq_ary[15][41] ,
         \inq_ary[15][40] , \inq_ary[15][39] , \inq_ary[15][38] ,
         \inq_ary[15][37] , \inq_ary[15][36] , \inq_ary[15][35] ,
         \inq_ary[15][34] , \inq_ary[15][33] , \inq_ary[15][32] ,
         \inq_ary[15][31] , \inq_ary[15][30] , \inq_ary[15][29] ,
         \inq_ary[15][28] , \inq_ary[15][27] , \inq_ary[15][26] ,
         \inq_ary[15][25] , \inq_ary[15][24] , \inq_ary[15][23] ,
         \inq_ary[15][22] , \inq_ary[15][21] , \inq_ary[15][20] ,
         \inq_ary[15][19] , \inq_ary[15][18] , \inq_ary[15][17] ,
         \inq_ary[15][16] , \inq_ary[15][15] , \inq_ary[15][14] ,
         \inq_ary[15][13] , \inq_ary[15][12] , \inq_ary[15][11] ,
         \inq_ary[15][10] , \inq_ary[15][9] , \inq_ary[15][8] ,
         \inq_ary[15][7] , \inq_ary[15][6] , \inq_ary[15][5] ,
         \inq_ary[15][4] , \inq_ary[15][3] , \inq_ary[15][2] ,
         \inq_ary[15][1] , \inq_ary[15][0] , \inq_ary[14][159] ,
         \inq_ary[14][158] , \inq_ary[14][157] , \inq_ary[14][156] ,
         \inq_ary[14][155] , \inq_ary[14][154] , \inq_ary[14][153] ,
         \inq_ary[14][152] , \inq_ary[14][151] , \inq_ary[14][150] ,
         \inq_ary[14][149] , \inq_ary[14][148] , \inq_ary[14][147] ,
         \inq_ary[14][146] , \inq_ary[14][145] , \inq_ary[14][144] ,
         \inq_ary[14][143] , \inq_ary[14][142] , \inq_ary[14][141] ,
         \inq_ary[14][140] , \inq_ary[14][139] , \inq_ary[14][138] ,
         \inq_ary[14][137] , \inq_ary[14][136] , \inq_ary[14][135] ,
         \inq_ary[14][134] , \inq_ary[14][133] , \inq_ary[14][132] ,
         \inq_ary[14][131] , \inq_ary[14][130] , \inq_ary[14][129] ,
         \inq_ary[14][128] , \inq_ary[14][127] , \inq_ary[14][126] ,
         \inq_ary[14][125] , \inq_ary[14][124] , \inq_ary[14][123] ,
         \inq_ary[14][122] , \inq_ary[14][121] , \inq_ary[14][120] ,
         \inq_ary[14][119] , \inq_ary[14][118] , \inq_ary[14][117] ,
         \inq_ary[14][116] , \inq_ary[14][115] , \inq_ary[14][114] ,
         \inq_ary[14][113] , \inq_ary[14][112] , \inq_ary[14][111] ,
         \inq_ary[14][110] , \inq_ary[14][109] , \inq_ary[14][108] ,
         \inq_ary[14][107] , \inq_ary[14][106] , \inq_ary[14][105] ,
         \inq_ary[14][104] , \inq_ary[14][103] , \inq_ary[14][102] ,
         \inq_ary[14][101] , \inq_ary[14][100] , \inq_ary[14][99] ,
         \inq_ary[14][98] , \inq_ary[14][97] , \inq_ary[14][96] ,
         \inq_ary[14][95] , \inq_ary[14][94] , \inq_ary[14][93] ,
         \inq_ary[14][92] , \inq_ary[14][91] , \inq_ary[14][90] ,
         \inq_ary[14][89] , \inq_ary[14][88] , \inq_ary[14][87] ,
         \inq_ary[14][86] , \inq_ary[14][85] , \inq_ary[14][84] ,
         \inq_ary[14][83] , \inq_ary[14][82] , \inq_ary[14][81] ,
         \inq_ary[14][80] , \inq_ary[14][79] , \inq_ary[14][78] ,
         \inq_ary[14][77] , \inq_ary[14][76] , \inq_ary[14][75] ,
         \inq_ary[14][74] , \inq_ary[14][73] , \inq_ary[14][72] ,
         \inq_ary[14][71] , \inq_ary[14][70] , \inq_ary[14][69] ,
         \inq_ary[14][68] , \inq_ary[14][67] , \inq_ary[14][66] ,
         \inq_ary[14][65] , \inq_ary[14][64] , \inq_ary[14][63] ,
         \inq_ary[14][62] , \inq_ary[14][61] , \inq_ary[14][60] ,
         \inq_ary[14][59] , \inq_ary[14][58] , \inq_ary[14][57] ,
         \inq_ary[14][56] , \inq_ary[14][55] , \inq_ary[14][54] ,
         \inq_ary[14][53] , \inq_ary[14][52] , \inq_ary[14][51] ,
         \inq_ary[14][50] , \inq_ary[14][49] , \inq_ary[14][48] ,
         \inq_ary[14][47] , \inq_ary[14][46] , \inq_ary[14][45] ,
         \inq_ary[14][44] , \inq_ary[14][43] , \inq_ary[14][42] ,
         \inq_ary[14][41] , \inq_ary[14][40] , \inq_ary[14][39] ,
         \inq_ary[14][38] , \inq_ary[14][37] , \inq_ary[14][36] ,
         \inq_ary[14][35] , \inq_ary[14][34] , \inq_ary[14][33] ,
         \inq_ary[14][32] , \inq_ary[14][31] , \inq_ary[14][30] ,
         \inq_ary[14][29] , \inq_ary[14][28] , \inq_ary[14][27] ,
         \inq_ary[14][26] , \inq_ary[14][25] , \inq_ary[14][24] ,
         \inq_ary[14][23] , \inq_ary[14][22] , \inq_ary[14][21] ,
         \inq_ary[14][20] , \inq_ary[14][19] , \inq_ary[14][18] ,
         \inq_ary[14][17] , \inq_ary[14][16] , \inq_ary[14][15] ,
         \inq_ary[14][14] , \inq_ary[14][13] , \inq_ary[14][12] ,
         \inq_ary[14][11] , \inq_ary[14][10] , \inq_ary[14][9] ,
         \inq_ary[14][8] , \inq_ary[14][7] , \inq_ary[14][6] ,
         \inq_ary[14][5] , \inq_ary[14][4] , \inq_ary[14][3] ,
         \inq_ary[14][2] , \inq_ary[14][1] , \inq_ary[14][0] ,
         \inq_ary[13][159] , \inq_ary[13][158] , \inq_ary[13][157] ,
         \inq_ary[13][156] , \inq_ary[13][155] , \inq_ary[13][154] ,
         \inq_ary[13][153] , \inq_ary[13][152] , \inq_ary[13][151] ,
         \inq_ary[13][150] , \inq_ary[13][149] , \inq_ary[13][148] ,
         \inq_ary[13][147] , \inq_ary[13][146] , \inq_ary[13][145] ,
         \inq_ary[13][144] , \inq_ary[13][143] , \inq_ary[13][142] ,
         \inq_ary[13][141] , \inq_ary[13][140] , \inq_ary[13][139] ,
         \inq_ary[13][138] , \inq_ary[13][137] , \inq_ary[13][136] ,
         \inq_ary[13][135] , \inq_ary[13][134] , \inq_ary[13][133] ,
         \inq_ary[13][132] , \inq_ary[13][131] , \inq_ary[13][130] ,
         \inq_ary[13][129] , \inq_ary[13][128] , \inq_ary[13][127] ,
         \inq_ary[13][126] , \inq_ary[13][125] , \inq_ary[13][124] ,
         \inq_ary[13][123] , \inq_ary[13][122] , \inq_ary[13][121] ,
         \inq_ary[13][120] , \inq_ary[13][119] , \inq_ary[13][118] ,
         \inq_ary[13][117] , \inq_ary[13][116] , \inq_ary[13][115] ,
         \inq_ary[13][114] , \inq_ary[13][113] , \inq_ary[13][112] ,
         \inq_ary[13][111] , \inq_ary[13][110] , \inq_ary[13][109] ,
         \inq_ary[13][108] , \inq_ary[13][107] , \inq_ary[13][106] ,
         \inq_ary[13][105] , \inq_ary[13][104] , \inq_ary[13][103] ,
         \inq_ary[13][102] , \inq_ary[13][101] , \inq_ary[13][100] ,
         \inq_ary[13][99] , \inq_ary[13][98] , \inq_ary[13][97] ,
         \inq_ary[13][96] , \inq_ary[13][95] , \inq_ary[13][94] ,
         \inq_ary[13][93] , \inq_ary[13][92] , \inq_ary[13][91] ,
         \inq_ary[13][90] , \inq_ary[13][89] , \inq_ary[13][88] ,
         \inq_ary[13][87] , \inq_ary[13][86] , \inq_ary[13][85] ,
         \inq_ary[13][84] , \inq_ary[13][83] , \inq_ary[13][82] ,
         \inq_ary[13][81] , \inq_ary[13][80] , \inq_ary[13][79] ,
         \inq_ary[13][78] , \inq_ary[13][77] , \inq_ary[13][76] ,
         \inq_ary[13][75] , \inq_ary[13][74] , \inq_ary[13][73] ,
         \inq_ary[13][72] , \inq_ary[13][71] , \inq_ary[13][70] ,
         \inq_ary[13][69] , \inq_ary[13][68] , \inq_ary[13][67] ,
         \inq_ary[13][66] , \inq_ary[13][65] , \inq_ary[13][64] ,
         \inq_ary[13][63] , \inq_ary[13][62] , \inq_ary[13][61] ,
         \inq_ary[13][60] , \inq_ary[13][59] , \inq_ary[13][58] ,
         \inq_ary[13][57] , \inq_ary[13][56] , \inq_ary[13][55] ,
         \inq_ary[13][54] , \inq_ary[13][53] , \inq_ary[13][52] ,
         \inq_ary[13][51] , \inq_ary[13][50] , \inq_ary[13][49] ,
         \inq_ary[13][48] , \inq_ary[13][47] , \inq_ary[13][46] ,
         \inq_ary[13][45] , \inq_ary[13][44] , \inq_ary[13][43] ,
         \inq_ary[13][42] , \inq_ary[13][41] , \inq_ary[13][40] ,
         \inq_ary[13][39] , \inq_ary[13][38] , \inq_ary[13][37] ,
         \inq_ary[13][36] , \inq_ary[13][35] , \inq_ary[13][34] ,
         \inq_ary[13][33] , \inq_ary[13][32] , \inq_ary[13][31] ,
         \inq_ary[13][30] , \inq_ary[13][29] , \inq_ary[13][28] ,
         \inq_ary[13][27] , \inq_ary[13][26] , \inq_ary[13][25] ,
         \inq_ary[13][24] , \inq_ary[13][23] , \inq_ary[13][22] ,
         \inq_ary[13][21] , \inq_ary[13][20] , \inq_ary[13][19] ,
         \inq_ary[13][18] , \inq_ary[13][17] , \inq_ary[13][16] ,
         \inq_ary[13][15] , \inq_ary[13][14] , \inq_ary[13][13] ,
         \inq_ary[13][12] , \inq_ary[13][11] , \inq_ary[13][10] ,
         \inq_ary[13][9] , \inq_ary[13][8] , \inq_ary[13][7] ,
         \inq_ary[13][6] , \inq_ary[13][5] , \inq_ary[13][4] ,
         \inq_ary[13][3] , \inq_ary[13][2] , \inq_ary[13][1] ,
         \inq_ary[13][0] , \inq_ary[12][159] , \inq_ary[12][158] ,
         \inq_ary[12][157] , \inq_ary[12][156] , \inq_ary[12][155] ,
         \inq_ary[12][154] , \inq_ary[12][153] , \inq_ary[12][152] ,
         \inq_ary[12][151] , \inq_ary[12][150] , \inq_ary[12][149] ,
         \inq_ary[12][148] , \inq_ary[12][147] , \inq_ary[12][146] ,
         \inq_ary[12][145] , \inq_ary[12][144] , \inq_ary[12][143] ,
         \inq_ary[12][142] , \inq_ary[12][141] , \inq_ary[12][140] ,
         \inq_ary[12][139] , \inq_ary[12][138] , \inq_ary[12][137] ,
         \inq_ary[12][136] , \inq_ary[12][135] , \inq_ary[12][134] ,
         \inq_ary[12][133] , \inq_ary[12][132] , \inq_ary[12][131] ,
         \inq_ary[12][130] , \inq_ary[12][129] , \inq_ary[12][128] ,
         \inq_ary[12][127] , \inq_ary[12][126] , \inq_ary[12][125] ,
         \inq_ary[12][124] , \inq_ary[12][123] , \inq_ary[12][122] ,
         \inq_ary[12][121] , \inq_ary[12][120] , \inq_ary[12][119] ,
         \inq_ary[12][118] , \inq_ary[12][117] , \inq_ary[12][116] ,
         \inq_ary[12][115] , \inq_ary[12][114] , \inq_ary[12][113] ,
         \inq_ary[12][112] , \inq_ary[12][111] , \inq_ary[12][110] ,
         \inq_ary[12][109] , \inq_ary[12][108] , \inq_ary[12][107] ,
         \inq_ary[12][106] , \inq_ary[12][105] , \inq_ary[12][104] ,
         \inq_ary[12][103] , \inq_ary[12][102] , \inq_ary[12][101] ,
         \inq_ary[12][100] , \inq_ary[12][99] , \inq_ary[12][98] ,
         \inq_ary[12][97] , \inq_ary[12][96] , \inq_ary[12][95] ,
         \inq_ary[12][94] , \inq_ary[12][93] , \inq_ary[12][92] ,
         \inq_ary[12][91] , \inq_ary[12][90] , \inq_ary[12][89] ,
         \inq_ary[12][88] , \inq_ary[12][87] , \inq_ary[12][86] ,
         \inq_ary[12][85] , \inq_ary[12][84] , \inq_ary[12][83] ,
         \inq_ary[12][82] , \inq_ary[12][81] , \inq_ary[12][80] ,
         \inq_ary[12][79] , \inq_ary[12][78] , \inq_ary[12][77] ,
         \inq_ary[12][76] , \inq_ary[12][75] , \inq_ary[12][74] ,
         \inq_ary[12][73] , \inq_ary[12][72] , \inq_ary[12][71] ,
         \inq_ary[12][70] , \inq_ary[12][69] , \inq_ary[12][68] ,
         \inq_ary[12][67] , \inq_ary[12][66] , \inq_ary[12][65] ,
         \inq_ary[12][64] , \inq_ary[12][63] , \inq_ary[12][62] ,
         \inq_ary[12][61] , \inq_ary[12][60] , \inq_ary[12][59] ,
         \inq_ary[12][58] , \inq_ary[12][57] , \inq_ary[12][56] ,
         \inq_ary[12][55] , \inq_ary[12][54] , \inq_ary[12][53] ,
         \inq_ary[12][52] , \inq_ary[12][51] , \inq_ary[12][50] ,
         \inq_ary[12][49] , \inq_ary[12][48] , \inq_ary[12][47] ,
         \inq_ary[12][46] , \inq_ary[12][45] , \inq_ary[12][44] ,
         \inq_ary[12][43] , \inq_ary[12][42] , \inq_ary[12][41] ,
         \inq_ary[12][40] , \inq_ary[12][39] , \inq_ary[12][38] ,
         \inq_ary[12][37] , \inq_ary[12][36] , \inq_ary[12][35] ,
         \inq_ary[12][34] , \inq_ary[12][33] , \inq_ary[12][32] ,
         \inq_ary[12][31] , \inq_ary[12][30] , \inq_ary[12][29] ,
         \inq_ary[12][28] , \inq_ary[12][27] , \inq_ary[12][26] ,
         \inq_ary[12][25] , \inq_ary[12][24] , \inq_ary[12][23] ,
         \inq_ary[12][22] , \inq_ary[12][21] , \inq_ary[12][20] ,
         \inq_ary[12][19] , \inq_ary[12][18] , \inq_ary[12][17] ,
         \inq_ary[12][16] , \inq_ary[12][15] , \inq_ary[12][14] ,
         \inq_ary[12][13] , \inq_ary[12][12] , \inq_ary[12][11] ,
         \inq_ary[12][10] , \inq_ary[12][9] , \inq_ary[12][8] ,
         \inq_ary[12][7] , \inq_ary[12][6] , \inq_ary[12][5] ,
         \inq_ary[12][4] , \inq_ary[12][3] , \inq_ary[12][2] ,
         \inq_ary[12][1] , \inq_ary[12][0] , \inq_ary[11][159] ,
         \inq_ary[11][158] , \inq_ary[11][157] , \inq_ary[11][156] ,
         \inq_ary[11][155] , \inq_ary[11][154] , \inq_ary[11][153] ,
         \inq_ary[11][152] , \inq_ary[11][151] , \inq_ary[11][150] ,
         \inq_ary[11][149] , \inq_ary[11][148] , \inq_ary[11][147] ,
         \inq_ary[11][146] , \inq_ary[11][145] , \inq_ary[11][144] ,
         \inq_ary[11][143] , \inq_ary[11][142] , \inq_ary[11][141] ,
         \inq_ary[11][140] , \inq_ary[11][139] , \inq_ary[11][138] ,
         \inq_ary[11][137] , \inq_ary[11][136] , \inq_ary[11][135] ,
         \inq_ary[11][134] , \inq_ary[11][133] , \inq_ary[11][132] ,
         \inq_ary[11][131] , \inq_ary[11][130] , \inq_ary[11][129] ,
         \inq_ary[11][128] , \inq_ary[11][127] , \inq_ary[11][126] ,
         \inq_ary[11][125] , \inq_ary[11][124] , \inq_ary[11][123] ,
         \inq_ary[11][122] , \inq_ary[11][121] , \inq_ary[11][120] ,
         \inq_ary[11][119] , \inq_ary[11][118] , \inq_ary[11][117] ,
         \inq_ary[11][116] , \inq_ary[11][115] , \inq_ary[11][114] ,
         \inq_ary[11][113] , \inq_ary[11][112] , \inq_ary[11][111] ,
         \inq_ary[11][110] , \inq_ary[11][109] , \inq_ary[11][108] ,
         \inq_ary[11][107] , \inq_ary[11][106] , \inq_ary[11][105] ,
         \inq_ary[11][104] , \inq_ary[11][103] , \inq_ary[11][102] ,
         \inq_ary[11][101] , \inq_ary[11][100] , \inq_ary[11][99] ,
         \inq_ary[11][98] , \inq_ary[11][97] , \inq_ary[11][96] ,
         \inq_ary[11][95] , \inq_ary[11][94] , \inq_ary[11][93] ,
         \inq_ary[11][92] , \inq_ary[11][91] , \inq_ary[11][90] ,
         \inq_ary[11][89] , \inq_ary[11][88] , \inq_ary[11][87] ,
         \inq_ary[11][86] , \inq_ary[11][85] , \inq_ary[11][84] ,
         \inq_ary[11][83] , \inq_ary[11][82] , \inq_ary[11][81] ,
         \inq_ary[11][80] , \inq_ary[11][79] , \inq_ary[11][78] ,
         \inq_ary[11][77] , \inq_ary[11][76] , \inq_ary[11][75] ,
         \inq_ary[11][74] , \inq_ary[11][73] , \inq_ary[11][72] ,
         \inq_ary[11][71] , \inq_ary[11][70] , \inq_ary[11][69] ,
         \inq_ary[11][68] , \inq_ary[11][67] , \inq_ary[11][66] ,
         \inq_ary[11][65] , \inq_ary[11][64] , \inq_ary[11][63] ,
         \inq_ary[11][62] , \inq_ary[11][61] , \inq_ary[11][60] ,
         \inq_ary[11][59] , \inq_ary[11][58] , \inq_ary[11][57] ,
         \inq_ary[11][56] , \inq_ary[11][55] , \inq_ary[11][54] ,
         \inq_ary[11][53] , \inq_ary[11][52] , \inq_ary[11][51] ,
         \inq_ary[11][50] , \inq_ary[11][49] , \inq_ary[11][48] ,
         \inq_ary[11][47] , \inq_ary[11][46] , \inq_ary[11][45] ,
         \inq_ary[11][44] , \inq_ary[11][43] , \inq_ary[11][42] ,
         \inq_ary[11][41] , \inq_ary[11][40] , \inq_ary[11][39] ,
         \inq_ary[11][38] , \inq_ary[11][37] , \inq_ary[11][36] ,
         \inq_ary[11][35] , \inq_ary[11][34] , \inq_ary[11][33] ,
         \inq_ary[11][32] , \inq_ary[11][31] , \inq_ary[11][30] ,
         \inq_ary[11][29] , \inq_ary[11][28] , \inq_ary[11][27] ,
         \inq_ary[11][26] , \inq_ary[11][25] , \inq_ary[11][24] ,
         \inq_ary[11][23] , \inq_ary[11][22] , \inq_ary[11][21] ,
         \inq_ary[11][20] , \inq_ary[11][19] , \inq_ary[11][18] ,
         \inq_ary[11][17] , \inq_ary[11][16] , \inq_ary[11][15] ,
         \inq_ary[11][14] , \inq_ary[11][13] , \inq_ary[11][12] ,
         \inq_ary[11][11] , \inq_ary[11][10] , \inq_ary[11][9] ,
         \inq_ary[11][8] , \inq_ary[11][7] , \inq_ary[11][6] ,
         \inq_ary[11][5] , \inq_ary[11][4] , \inq_ary[11][3] ,
         \inq_ary[11][2] , \inq_ary[11][1] , \inq_ary[11][0] ,
         \inq_ary[10][159] , \inq_ary[10][158] , \inq_ary[10][157] ,
         \inq_ary[10][156] , \inq_ary[10][155] , \inq_ary[10][154] ,
         \inq_ary[10][153] , \inq_ary[10][152] , \inq_ary[10][151] ,
         \inq_ary[10][150] , \inq_ary[10][149] , \inq_ary[10][148] ,
         \inq_ary[10][147] , \inq_ary[10][146] , \inq_ary[10][145] ,
         \inq_ary[10][144] , \inq_ary[10][143] , \inq_ary[10][142] ,
         \inq_ary[10][141] , \inq_ary[10][140] , \inq_ary[10][139] ,
         \inq_ary[10][138] , \inq_ary[10][137] , \inq_ary[10][136] ,
         \inq_ary[10][135] , \inq_ary[10][134] , \inq_ary[10][133] ,
         \inq_ary[10][132] , \inq_ary[10][131] , \inq_ary[10][130] ,
         \inq_ary[10][129] , \inq_ary[10][128] , \inq_ary[10][127] ,
         \inq_ary[10][126] , \inq_ary[10][125] , \inq_ary[10][124] ,
         \inq_ary[10][123] , \inq_ary[10][122] , \inq_ary[10][121] ,
         \inq_ary[10][120] , \inq_ary[10][119] , \inq_ary[10][118] ,
         \inq_ary[10][117] , \inq_ary[10][116] , \inq_ary[10][115] ,
         \inq_ary[10][114] , \inq_ary[10][113] , \inq_ary[10][112] ,
         \inq_ary[10][111] , \inq_ary[10][110] , \inq_ary[10][109] ,
         \inq_ary[10][108] , \inq_ary[10][107] , \inq_ary[10][106] ,
         \inq_ary[10][105] , \inq_ary[10][104] , \inq_ary[10][103] ,
         \inq_ary[10][102] , \inq_ary[10][101] , \inq_ary[10][100] ,
         \inq_ary[10][99] , \inq_ary[10][98] , \inq_ary[10][97] ,
         \inq_ary[10][96] , \inq_ary[10][95] , \inq_ary[10][94] ,
         \inq_ary[10][93] , \inq_ary[10][92] , \inq_ary[10][91] ,
         \inq_ary[10][90] , \inq_ary[10][89] , \inq_ary[10][88] ,
         \inq_ary[10][87] , \inq_ary[10][86] , \inq_ary[10][85] ,
         \inq_ary[10][84] , \inq_ary[10][83] , \inq_ary[10][82] ,
         \inq_ary[10][81] , \inq_ary[10][80] , \inq_ary[10][79] ,
         \inq_ary[10][78] , \inq_ary[10][77] , \inq_ary[10][76] ,
         \inq_ary[10][75] , \inq_ary[10][74] , \inq_ary[10][73] ,
         \inq_ary[10][72] , \inq_ary[10][71] , \inq_ary[10][70] ,
         \inq_ary[10][69] , \inq_ary[10][68] , \inq_ary[10][67] ,
         \inq_ary[10][66] , \inq_ary[10][65] , \inq_ary[10][64] ,
         \inq_ary[10][63] , \inq_ary[10][62] , \inq_ary[10][61] ,
         \inq_ary[10][60] , \inq_ary[10][59] , \inq_ary[10][58] ,
         \inq_ary[10][57] , \inq_ary[10][56] , \inq_ary[10][55] ,
         \inq_ary[10][54] , \inq_ary[10][53] , \inq_ary[10][52] ,
         \inq_ary[10][51] , \inq_ary[10][50] , \inq_ary[10][49] ,
         \inq_ary[10][48] , \inq_ary[10][47] , \inq_ary[10][46] ,
         \inq_ary[10][45] , \inq_ary[10][44] , \inq_ary[10][43] ,
         \inq_ary[10][42] , \inq_ary[10][41] , \inq_ary[10][40] ,
         \inq_ary[10][39] , \inq_ary[10][38] , \inq_ary[10][37] ,
         \inq_ary[10][36] , \inq_ary[10][35] , \inq_ary[10][34] ,
         \inq_ary[10][33] , \inq_ary[10][32] , \inq_ary[10][31] ,
         \inq_ary[10][30] , \inq_ary[10][29] , \inq_ary[10][28] ,
         \inq_ary[10][27] , \inq_ary[10][26] , \inq_ary[10][25] ,
         \inq_ary[10][24] , \inq_ary[10][23] , \inq_ary[10][22] ,
         \inq_ary[10][21] , \inq_ary[10][20] , \inq_ary[10][19] ,
         \inq_ary[10][18] , \inq_ary[10][17] , \inq_ary[10][16] ,
         \inq_ary[10][15] , \inq_ary[10][14] , \inq_ary[10][13] ,
         \inq_ary[10][12] , \inq_ary[10][11] , \inq_ary[10][10] ,
         \inq_ary[10][9] , \inq_ary[10][8] , \inq_ary[10][7] ,
         \inq_ary[10][6] , \inq_ary[10][5] , \inq_ary[10][4] ,
         \inq_ary[10][3] , \inq_ary[10][2] , \inq_ary[10][1] ,
         \inq_ary[10][0] , \inq_ary[9][159] , \inq_ary[9][158] ,
         \inq_ary[9][157] , \inq_ary[9][156] , \inq_ary[9][155] ,
         \inq_ary[9][154] , \inq_ary[9][153] , \inq_ary[9][152] ,
         \inq_ary[9][151] , \inq_ary[9][150] , \inq_ary[9][149] ,
         \inq_ary[9][148] , \inq_ary[9][147] , \inq_ary[9][146] ,
         \inq_ary[9][145] , \inq_ary[9][144] , \inq_ary[9][143] ,
         \inq_ary[9][142] , \inq_ary[9][141] , \inq_ary[9][140] ,
         \inq_ary[9][139] , \inq_ary[9][138] , \inq_ary[9][137] ,
         \inq_ary[9][136] , \inq_ary[9][135] , \inq_ary[9][134] ,
         \inq_ary[9][133] , \inq_ary[9][132] , \inq_ary[9][131] ,
         \inq_ary[9][130] , \inq_ary[9][129] , \inq_ary[9][128] ,
         \inq_ary[9][127] , \inq_ary[9][126] , \inq_ary[9][125] ,
         \inq_ary[9][124] , \inq_ary[9][123] , \inq_ary[9][122] ,
         \inq_ary[9][121] , \inq_ary[9][120] , \inq_ary[9][119] ,
         \inq_ary[9][118] , \inq_ary[9][117] , \inq_ary[9][116] ,
         \inq_ary[9][115] , \inq_ary[9][114] , \inq_ary[9][113] ,
         \inq_ary[9][112] , \inq_ary[9][111] , \inq_ary[9][110] ,
         \inq_ary[9][109] , \inq_ary[9][108] , \inq_ary[9][107] ,
         \inq_ary[9][106] , \inq_ary[9][105] , \inq_ary[9][104] ,
         \inq_ary[9][103] , \inq_ary[9][102] , \inq_ary[9][101] ,
         \inq_ary[9][100] , \inq_ary[9][99] , \inq_ary[9][98] ,
         \inq_ary[9][97] , \inq_ary[9][96] , \inq_ary[9][95] ,
         \inq_ary[9][94] , \inq_ary[9][93] , \inq_ary[9][92] ,
         \inq_ary[9][91] , \inq_ary[9][90] , \inq_ary[9][89] ,
         \inq_ary[9][88] , \inq_ary[9][87] , \inq_ary[9][86] ,
         \inq_ary[9][85] , \inq_ary[9][84] , \inq_ary[9][83] ,
         \inq_ary[9][82] , \inq_ary[9][81] , \inq_ary[9][80] ,
         \inq_ary[9][79] , \inq_ary[9][78] , \inq_ary[9][77] ,
         \inq_ary[9][76] , \inq_ary[9][75] , \inq_ary[9][74] ,
         \inq_ary[9][73] , \inq_ary[9][72] , \inq_ary[9][71] ,
         \inq_ary[9][70] , \inq_ary[9][69] , \inq_ary[9][68] ,
         \inq_ary[9][67] , \inq_ary[9][66] , \inq_ary[9][65] ,
         \inq_ary[9][64] , \inq_ary[9][63] , \inq_ary[9][62] ,
         \inq_ary[9][61] , \inq_ary[9][60] , \inq_ary[9][59] ,
         \inq_ary[9][58] , \inq_ary[9][57] , \inq_ary[9][56] ,
         \inq_ary[9][55] , \inq_ary[9][54] , \inq_ary[9][53] ,
         \inq_ary[9][52] , \inq_ary[9][51] , \inq_ary[9][50] ,
         \inq_ary[9][49] , \inq_ary[9][48] , \inq_ary[9][47] ,
         \inq_ary[9][46] , \inq_ary[9][45] , \inq_ary[9][44] ,
         \inq_ary[9][43] , \inq_ary[9][42] , \inq_ary[9][41] ,
         \inq_ary[9][40] , \inq_ary[9][39] , \inq_ary[9][38] ,
         \inq_ary[9][37] , \inq_ary[9][36] , \inq_ary[9][35] ,
         \inq_ary[9][34] , \inq_ary[9][33] , \inq_ary[9][32] ,
         \inq_ary[9][31] , \inq_ary[9][30] , \inq_ary[9][29] ,
         \inq_ary[9][28] , \inq_ary[9][27] , \inq_ary[9][26] ,
         \inq_ary[9][25] , \inq_ary[9][24] , \inq_ary[9][23] ,
         \inq_ary[9][22] , \inq_ary[9][21] , \inq_ary[9][20] ,
         \inq_ary[9][19] , \inq_ary[9][18] , \inq_ary[9][17] ,
         \inq_ary[9][16] , \inq_ary[9][15] , \inq_ary[9][14] ,
         \inq_ary[9][13] , \inq_ary[9][12] , \inq_ary[9][11] ,
         \inq_ary[9][10] , \inq_ary[9][9] , \inq_ary[9][8] , \inq_ary[9][7] ,
         \inq_ary[9][6] , \inq_ary[9][5] , \inq_ary[9][4] , \inq_ary[9][3] ,
         \inq_ary[9][2] , \inq_ary[9][1] , \inq_ary[9][0] , \inq_ary[8][159] ,
         \inq_ary[8][158] , \inq_ary[8][157] , \inq_ary[8][156] ,
         \inq_ary[8][155] , \inq_ary[8][154] , \inq_ary[8][153] ,
         \inq_ary[8][152] , \inq_ary[8][151] , \inq_ary[8][150] ,
         \inq_ary[8][149] , \inq_ary[8][148] , \inq_ary[8][147] ,
         \inq_ary[8][146] , \inq_ary[8][145] , \inq_ary[8][144] ,
         \inq_ary[8][143] , \inq_ary[8][142] , \inq_ary[8][141] ,
         \inq_ary[8][140] , \inq_ary[8][139] , \inq_ary[8][138] ,
         \inq_ary[8][137] , \inq_ary[8][136] , \inq_ary[8][135] ,
         \inq_ary[8][134] , \inq_ary[8][133] , \inq_ary[8][132] ,
         \inq_ary[8][131] , \inq_ary[8][130] , \inq_ary[8][129] ,
         \inq_ary[8][128] , \inq_ary[8][127] , \inq_ary[8][126] ,
         \inq_ary[8][125] , \inq_ary[8][124] , \inq_ary[8][123] ,
         \inq_ary[8][122] , \inq_ary[8][121] , \inq_ary[8][120] ,
         \inq_ary[8][119] , \inq_ary[8][118] , \inq_ary[8][117] ,
         \inq_ary[8][116] , \inq_ary[8][115] , \inq_ary[8][114] ,
         \inq_ary[8][113] , \inq_ary[8][112] , \inq_ary[8][111] ,
         \inq_ary[8][110] , \inq_ary[8][109] , \inq_ary[8][108] ,
         \inq_ary[8][107] , \inq_ary[8][106] , \inq_ary[8][105] ,
         \inq_ary[8][104] , \inq_ary[8][103] , \inq_ary[8][102] ,
         \inq_ary[8][101] , \inq_ary[8][100] , \inq_ary[8][99] ,
         \inq_ary[8][98] , \inq_ary[8][97] , \inq_ary[8][96] ,
         \inq_ary[8][95] , \inq_ary[8][94] , \inq_ary[8][93] ,
         \inq_ary[8][92] , \inq_ary[8][91] , \inq_ary[8][90] ,
         \inq_ary[8][89] , \inq_ary[8][88] , \inq_ary[8][87] ,
         \inq_ary[8][86] , \inq_ary[8][85] , \inq_ary[8][84] ,
         \inq_ary[8][83] , \inq_ary[8][82] , \inq_ary[8][81] ,
         \inq_ary[8][80] , \inq_ary[8][79] , \inq_ary[8][78] ,
         \inq_ary[8][77] , \inq_ary[8][76] , \inq_ary[8][75] ,
         \inq_ary[8][74] , \inq_ary[8][73] , \inq_ary[8][72] ,
         \inq_ary[8][71] , \inq_ary[8][70] , \inq_ary[8][69] ,
         \inq_ary[8][68] , \inq_ary[8][67] , \inq_ary[8][66] ,
         \inq_ary[8][65] , \inq_ary[8][64] , \inq_ary[8][63] ,
         \inq_ary[8][62] , \inq_ary[8][61] , \inq_ary[8][60] ,
         \inq_ary[8][59] , \inq_ary[8][58] , \inq_ary[8][57] ,
         \inq_ary[8][56] , \inq_ary[8][55] , \inq_ary[8][54] ,
         \inq_ary[8][53] , \inq_ary[8][52] , \inq_ary[8][51] ,
         \inq_ary[8][50] , \inq_ary[8][49] , \inq_ary[8][48] ,
         \inq_ary[8][47] , \inq_ary[8][46] , \inq_ary[8][45] ,
         \inq_ary[8][44] , \inq_ary[8][43] , \inq_ary[8][42] ,
         \inq_ary[8][41] , \inq_ary[8][40] , \inq_ary[8][39] ,
         \inq_ary[8][38] , \inq_ary[8][37] , \inq_ary[8][36] ,
         \inq_ary[8][35] , \inq_ary[8][34] , \inq_ary[8][33] ,
         \inq_ary[8][32] , \inq_ary[8][31] , \inq_ary[8][30] ,
         \inq_ary[8][29] , \inq_ary[8][28] , \inq_ary[8][27] ,
         \inq_ary[8][26] , \inq_ary[8][25] , \inq_ary[8][24] ,
         \inq_ary[8][23] , \inq_ary[8][22] , \inq_ary[8][21] ,
         \inq_ary[8][20] , \inq_ary[8][19] , \inq_ary[8][18] ,
         \inq_ary[8][17] , \inq_ary[8][16] , \inq_ary[8][15] ,
         \inq_ary[8][14] , \inq_ary[8][13] , \inq_ary[8][12] ,
         \inq_ary[8][11] , \inq_ary[8][10] , \inq_ary[8][9] , \inq_ary[8][8] ,
         \inq_ary[8][7] , \inq_ary[8][6] , \inq_ary[8][5] , \inq_ary[8][4] ,
         \inq_ary[8][3] , \inq_ary[8][2] , \inq_ary[8][1] , \inq_ary[8][0] ,
         \inq_ary[7][159] , \inq_ary[7][158] , \inq_ary[7][157] ,
         \inq_ary[7][156] , \inq_ary[7][155] , \inq_ary[7][154] ,
         \inq_ary[7][153] , \inq_ary[7][152] , \inq_ary[7][151] ,
         \inq_ary[7][150] , \inq_ary[7][149] , \inq_ary[7][148] ,
         \inq_ary[7][147] , \inq_ary[7][146] , \inq_ary[7][145] ,
         \inq_ary[7][144] , \inq_ary[7][143] , \inq_ary[7][142] ,
         \inq_ary[7][141] , \inq_ary[7][140] , \inq_ary[7][139] ,
         \inq_ary[7][138] , \inq_ary[7][137] , \inq_ary[7][136] ,
         \inq_ary[7][135] , \inq_ary[7][134] , \inq_ary[7][133] ,
         \inq_ary[7][132] , \inq_ary[7][131] , \inq_ary[7][130] ,
         \inq_ary[7][129] , \inq_ary[7][128] , \inq_ary[7][127] ,
         \inq_ary[7][126] , \inq_ary[7][125] , \inq_ary[7][124] ,
         \inq_ary[7][123] , \inq_ary[7][122] , \inq_ary[7][121] ,
         \inq_ary[7][120] , \inq_ary[7][119] , \inq_ary[7][118] ,
         \inq_ary[7][117] , \inq_ary[7][116] , \inq_ary[7][115] ,
         \inq_ary[7][114] , \inq_ary[7][113] , \inq_ary[7][112] ,
         \inq_ary[7][111] , \inq_ary[7][110] , \inq_ary[7][109] ,
         \inq_ary[7][108] , \inq_ary[7][107] , \inq_ary[7][106] ,
         \inq_ary[7][105] , \inq_ary[7][104] , \inq_ary[7][103] ,
         \inq_ary[7][102] , \inq_ary[7][101] , \inq_ary[7][100] ,
         \inq_ary[7][99] , \inq_ary[7][98] , \inq_ary[7][97] ,
         \inq_ary[7][96] , \inq_ary[7][95] , \inq_ary[7][94] ,
         \inq_ary[7][93] , \inq_ary[7][92] , \inq_ary[7][91] ,
         \inq_ary[7][90] , \inq_ary[7][89] , \inq_ary[7][88] ,
         \inq_ary[7][87] , \inq_ary[7][86] , \inq_ary[7][85] ,
         \inq_ary[7][84] , \inq_ary[7][83] , \inq_ary[7][82] ,
         \inq_ary[7][81] , \inq_ary[7][80] , \inq_ary[7][79] ,
         \inq_ary[7][78] , \inq_ary[7][77] , \inq_ary[7][76] ,
         \inq_ary[7][75] , \inq_ary[7][74] , \inq_ary[7][73] ,
         \inq_ary[7][72] , \inq_ary[7][71] , \inq_ary[7][70] ,
         \inq_ary[7][69] , \inq_ary[7][68] , \inq_ary[7][67] ,
         \inq_ary[7][66] , \inq_ary[7][65] , \inq_ary[7][64] ,
         \inq_ary[7][63] , \inq_ary[7][62] , \inq_ary[7][61] ,
         \inq_ary[7][60] , \inq_ary[7][59] , \inq_ary[7][58] ,
         \inq_ary[7][57] , \inq_ary[7][56] , \inq_ary[7][55] ,
         \inq_ary[7][54] , \inq_ary[7][53] , \inq_ary[7][52] ,
         \inq_ary[7][51] , \inq_ary[7][50] , \inq_ary[7][49] ,
         \inq_ary[7][48] , \inq_ary[7][47] , \inq_ary[7][46] ,
         \inq_ary[7][45] , \inq_ary[7][44] , \inq_ary[7][43] ,
         \inq_ary[7][42] , \inq_ary[7][41] , \inq_ary[7][40] ,
         \inq_ary[7][39] , \inq_ary[7][38] , \inq_ary[7][37] ,
         \inq_ary[7][36] , \inq_ary[7][35] , \inq_ary[7][34] ,
         \inq_ary[7][33] , \inq_ary[7][32] , \inq_ary[7][31] ,
         \inq_ary[7][30] , \inq_ary[7][29] , \inq_ary[7][28] ,
         \inq_ary[7][27] , \inq_ary[7][26] , \inq_ary[7][25] ,
         \inq_ary[7][24] , \inq_ary[7][23] , \inq_ary[7][22] ,
         \inq_ary[7][21] , \inq_ary[7][20] , \inq_ary[7][19] ,
         \inq_ary[7][18] , \inq_ary[7][17] , \inq_ary[7][16] ,
         \inq_ary[7][15] , \inq_ary[7][14] , \inq_ary[7][13] ,
         \inq_ary[7][12] , \inq_ary[7][11] , \inq_ary[7][10] , \inq_ary[7][9] ,
         \inq_ary[7][8] , \inq_ary[7][7] , \inq_ary[7][6] , \inq_ary[7][5] ,
         \inq_ary[7][4] , \inq_ary[7][3] , \inq_ary[7][2] , \inq_ary[7][1] ,
         \inq_ary[7][0] , \inq_ary[6][159] , \inq_ary[6][158] ,
         \inq_ary[6][157] , \inq_ary[6][156] , \inq_ary[6][155] ,
         \inq_ary[6][154] , \inq_ary[6][153] , \inq_ary[6][152] ,
         \inq_ary[6][151] , \inq_ary[6][150] , \inq_ary[6][149] ,
         \inq_ary[6][148] , \inq_ary[6][147] , \inq_ary[6][146] ,
         \inq_ary[6][145] , \inq_ary[6][144] , \inq_ary[6][143] ,
         \inq_ary[6][142] , \inq_ary[6][141] , \inq_ary[6][140] ,
         \inq_ary[6][139] , \inq_ary[6][138] , \inq_ary[6][137] ,
         \inq_ary[6][136] , \inq_ary[6][135] , \inq_ary[6][134] ,
         \inq_ary[6][133] , \inq_ary[6][132] , \inq_ary[6][131] ,
         \inq_ary[6][130] , \inq_ary[6][129] , \inq_ary[6][128] ,
         \inq_ary[6][127] , \inq_ary[6][126] , \inq_ary[6][125] ,
         \inq_ary[6][124] , \inq_ary[6][123] , \inq_ary[6][122] ,
         \inq_ary[6][121] , \inq_ary[6][120] , \inq_ary[6][119] ,
         \inq_ary[6][118] , \inq_ary[6][117] , \inq_ary[6][116] ,
         \inq_ary[6][115] , \inq_ary[6][114] , \inq_ary[6][113] ,
         \inq_ary[6][112] , \inq_ary[6][111] , \inq_ary[6][110] ,
         \inq_ary[6][109] , \inq_ary[6][108] , \inq_ary[6][107] ,
         \inq_ary[6][106] , \inq_ary[6][105] , \inq_ary[6][104] ,
         \inq_ary[6][103] , \inq_ary[6][102] , \inq_ary[6][101] ,
         \inq_ary[6][100] , \inq_ary[6][99] , \inq_ary[6][98] ,
         \inq_ary[6][97] , \inq_ary[6][96] , \inq_ary[6][95] ,
         \inq_ary[6][94] , \inq_ary[6][93] , \inq_ary[6][92] ,
         \inq_ary[6][91] , \inq_ary[6][90] , \inq_ary[6][89] ,
         \inq_ary[6][88] , \inq_ary[6][87] , \inq_ary[6][86] ,
         \inq_ary[6][85] , \inq_ary[6][84] , \inq_ary[6][83] ,
         \inq_ary[6][82] , \inq_ary[6][81] , \inq_ary[6][80] ,
         \inq_ary[6][79] , \inq_ary[6][78] , \inq_ary[6][77] ,
         \inq_ary[6][76] , \inq_ary[6][75] , \inq_ary[6][74] ,
         \inq_ary[6][73] , \inq_ary[6][72] , \inq_ary[6][71] ,
         \inq_ary[6][70] , \inq_ary[6][69] , \inq_ary[6][68] ,
         \inq_ary[6][67] , \inq_ary[6][66] , \inq_ary[6][65] ,
         \inq_ary[6][64] , \inq_ary[6][63] , \inq_ary[6][62] ,
         \inq_ary[6][61] , \inq_ary[6][60] , \inq_ary[6][59] ,
         \inq_ary[6][58] , \inq_ary[6][57] , \inq_ary[6][56] ,
         \inq_ary[6][55] , \inq_ary[6][54] , \inq_ary[6][53] ,
         \inq_ary[6][52] , \inq_ary[6][51] , \inq_ary[6][50] ,
         \inq_ary[6][49] , \inq_ary[6][48] , \inq_ary[6][47] ,
         \inq_ary[6][46] , \inq_ary[6][45] , \inq_ary[6][44] ,
         \inq_ary[6][43] , \inq_ary[6][42] , \inq_ary[6][41] ,
         \inq_ary[6][40] , \inq_ary[6][39] , \inq_ary[6][38] ,
         \inq_ary[6][37] , \inq_ary[6][36] , \inq_ary[6][35] ,
         \inq_ary[6][34] , \inq_ary[6][33] , \inq_ary[6][32] ,
         \inq_ary[6][31] , \inq_ary[6][30] , \inq_ary[6][29] ,
         \inq_ary[6][28] , \inq_ary[6][27] , \inq_ary[6][26] ,
         \inq_ary[6][25] , \inq_ary[6][24] , \inq_ary[6][23] ,
         \inq_ary[6][22] , \inq_ary[6][21] , \inq_ary[6][20] ,
         \inq_ary[6][19] , \inq_ary[6][18] , \inq_ary[6][17] ,
         \inq_ary[6][16] , \inq_ary[6][15] , \inq_ary[6][14] ,
         \inq_ary[6][13] , \inq_ary[6][12] , \inq_ary[6][11] ,
         \inq_ary[6][10] , \inq_ary[6][9] , \inq_ary[6][8] , \inq_ary[6][7] ,
         \inq_ary[6][6] , \inq_ary[6][5] , \inq_ary[6][4] , \inq_ary[6][3] ,
         \inq_ary[6][2] , \inq_ary[6][1] , \inq_ary[6][0] , \inq_ary[5][159] ,
         \inq_ary[5][158] , \inq_ary[5][157] , \inq_ary[5][156] ,
         \inq_ary[5][155] , \inq_ary[5][154] , \inq_ary[5][153] ,
         \inq_ary[5][152] , \inq_ary[5][151] , \inq_ary[5][150] ,
         \inq_ary[5][149] , \inq_ary[5][148] , \inq_ary[5][147] ,
         \inq_ary[5][146] , \inq_ary[5][145] , \inq_ary[5][144] ,
         \inq_ary[5][143] , \inq_ary[5][142] , \inq_ary[5][141] ,
         \inq_ary[5][140] , \inq_ary[5][139] , \inq_ary[5][138] ,
         \inq_ary[5][137] , \inq_ary[5][136] , \inq_ary[5][135] ,
         \inq_ary[5][134] , \inq_ary[5][133] , \inq_ary[5][132] ,
         \inq_ary[5][131] , \inq_ary[5][130] , \inq_ary[5][129] ,
         \inq_ary[5][128] , \inq_ary[5][127] , \inq_ary[5][126] ,
         \inq_ary[5][125] , \inq_ary[5][124] , \inq_ary[5][123] ,
         \inq_ary[5][122] , \inq_ary[5][121] , \inq_ary[5][120] ,
         \inq_ary[5][119] , \inq_ary[5][118] , \inq_ary[5][117] ,
         \inq_ary[5][116] , \inq_ary[5][115] , \inq_ary[5][114] ,
         \inq_ary[5][113] , \inq_ary[5][112] , \inq_ary[5][111] ,
         \inq_ary[5][110] , \inq_ary[5][109] , \inq_ary[5][108] ,
         \inq_ary[5][107] , \inq_ary[5][106] , \inq_ary[5][105] ,
         \inq_ary[5][104] , \inq_ary[5][103] , \inq_ary[5][102] ,
         \inq_ary[5][101] , \inq_ary[5][100] , \inq_ary[5][99] ,
         \inq_ary[5][98] , \inq_ary[5][97] , \inq_ary[5][96] ,
         \inq_ary[5][95] , \inq_ary[5][94] , \inq_ary[5][93] ,
         \inq_ary[5][92] , \inq_ary[5][91] , \inq_ary[5][90] ,
         \inq_ary[5][89] , \inq_ary[5][88] , \inq_ary[5][87] ,
         \inq_ary[5][86] , \inq_ary[5][85] , \inq_ary[5][84] ,
         \inq_ary[5][83] , \inq_ary[5][82] , \inq_ary[5][81] ,
         \inq_ary[5][80] , \inq_ary[5][79] , \inq_ary[5][78] ,
         \inq_ary[5][77] , \inq_ary[5][76] , \inq_ary[5][75] ,
         \inq_ary[5][74] , \inq_ary[5][73] , \inq_ary[5][72] ,
         \inq_ary[5][71] , \inq_ary[5][70] , \inq_ary[5][69] ,
         \inq_ary[5][68] , \inq_ary[5][67] , \inq_ary[5][66] ,
         \inq_ary[5][65] , \inq_ary[5][64] , \inq_ary[5][63] ,
         \inq_ary[5][62] , \inq_ary[5][61] , \inq_ary[5][60] ,
         \inq_ary[5][59] , \inq_ary[5][58] , \inq_ary[5][57] ,
         \inq_ary[5][56] , \inq_ary[5][55] , \inq_ary[5][54] ,
         \inq_ary[5][53] , \inq_ary[5][52] , \inq_ary[5][51] ,
         \inq_ary[5][50] , \inq_ary[5][49] , \inq_ary[5][48] ,
         \inq_ary[5][47] , \inq_ary[5][46] , \inq_ary[5][45] ,
         \inq_ary[5][44] , \inq_ary[5][43] , \inq_ary[5][42] ,
         \inq_ary[5][41] , \inq_ary[5][40] , \inq_ary[5][39] ,
         \inq_ary[5][38] , \inq_ary[5][37] , \inq_ary[5][36] ,
         \inq_ary[5][35] , \inq_ary[5][34] , \inq_ary[5][33] ,
         \inq_ary[5][32] , \inq_ary[5][31] , \inq_ary[5][30] ,
         \inq_ary[5][29] , \inq_ary[5][28] , \inq_ary[5][27] ,
         \inq_ary[5][26] , \inq_ary[5][25] , \inq_ary[5][24] ,
         \inq_ary[5][23] , \inq_ary[5][22] , \inq_ary[5][21] ,
         \inq_ary[5][20] , \inq_ary[5][19] , \inq_ary[5][18] ,
         \inq_ary[5][17] , \inq_ary[5][16] , \inq_ary[5][15] ,
         \inq_ary[5][14] , \inq_ary[5][13] , \inq_ary[5][12] ,
         \inq_ary[5][11] , \inq_ary[5][10] , \inq_ary[5][9] , \inq_ary[5][8] ,
         \inq_ary[5][7] , \inq_ary[5][6] , \inq_ary[5][5] , \inq_ary[5][4] ,
         \inq_ary[5][3] , \inq_ary[5][2] , \inq_ary[5][1] , \inq_ary[5][0] ,
         \inq_ary[4][159] , \inq_ary[4][158] , \inq_ary[4][157] ,
         \inq_ary[4][156] , \inq_ary[4][155] , \inq_ary[4][154] ,
         \inq_ary[4][153] , \inq_ary[4][152] , \inq_ary[4][151] ,
         \inq_ary[4][150] , \inq_ary[4][149] , \inq_ary[4][148] ,
         \inq_ary[4][147] , \inq_ary[4][146] , \inq_ary[4][145] ,
         \inq_ary[4][144] , \inq_ary[4][143] , \inq_ary[4][142] ,
         \inq_ary[4][141] , \inq_ary[4][140] , \inq_ary[4][139] ,
         \inq_ary[4][138] , \inq_ary[4][137] , \inq_ary[4][136] ,
         \inq_ary[4][135] , \inq_ary[4][134] , \inq_ary[4][133] ,
         \inq_ary[4][132] , \inq_ary[4][131] , \inq_ary[4][130] ,
         \inq_ary[4][129] , \inq_ary[4][128] , \inq_ary[4][127] ,
         \inq_ary[4][126] , \inq_ary[4][125] , \inq_ary[4][124] ,
         \inq_ary[4][123] , \inq_ary[4][122] , \inq_ary[4][121] ,
         \inq_ary[4][120] , \inq_ary[4][119] , \inq_ary[4][118] ,
         \inq_ary[4][117] , \inq_ary[4][116] , \inq_ary[4][115] ,
         \inq_ary[4][114] , \inq_ary[4][113] , \inq_ary[4][112] ,
         \inq_ary[4][111] , \inq_ary[4][110] , \inq_ary[4][109] ,
         \inq_ary[4][108] , \inq_ary[4][107] , \inq_ary[4][106] ,
         \inq_ary[4][105] , \inq_ary[4][104] , \inq_ary[4][103] ,
         \inq_ary[4][102] , \inq_ary[4][101] , \inq_ary[4][100] ,
         \inq_ary[4][99] , \inq_ary[4][98] , \inq_ary[4][97] ,
         \inq_ary[4][96] , \inq_ary[4][95] , \inq_ary[4][94] ,
         \inq_ary[4][93] , \inq_ary[4][92] , \inq_ary[4][91] ,
         \inq_ary[4][90] , \inq_ary[4][89] , \inq_ary[4][88] ,
         \inq_ary[4][87] , \inq_ary[4][86] , \inq_ary[4][85] ,
         \inq_ary[4][84] , \inq_ary[4][83] , \inq_ary[4][82] ,
         \inq_ary[4][81] , \inq_ary[4][80] , \inq_ary[4][79] ,
         \inq_ary[4][78] , \inq_ary[4][77] , \inq_ary[4][76] ,
         \inq_ary[4][75] , \inq_ary[4][74] , \inq_ary[4][73] ,
         \inq_ary[4][72] , \inq_ary[4][71] , \inq_ary[4][70] ,
         \inq_ary[4][69] , \inq_ary[4][68] , \inq_ary[4][67] ,
         \inq_ary[4][66] , \inq_ary[4][65] , \inq_ary[4][64] ,
         \inq_ary[4][63] , \inq_ary[4][62] , \inq_ary[4][61] ,
         \inq_ary[4][60] , \inq_ary[4][59] , \inq_ary[4][58] ,
         \inq_ary[4][57] , \inq_ary[4][56] , \inq_ary[4][55] ,
         \inq_ary[4][54] , \inq_ary[4][53] , \inq_ary[4][52] ,
         \inq_ary[4][51] , \inq_ary[4][50] , \inq_ary[4][49] ,
         \inq_ary[4][48] , \inq_ary[4][47] , \inq_ary[4][46] ,
         \inq_ary[4][45] , \inq_ary[4][44] , \inq_ary[4][43] ,
         \inq_ary[4][42] , \inq_ary[4][41] , \inq_ary[4][40] ,
         \inq_ary[4][39] , \inq_ary[4][38] , \inq_ary[4][37] ,
         \inq_ary[4][36] , \inq_ary[4][35] , \inq_ary[4][34] ,
         \inq_ary[4][33] , \inq_ary[4][32] , \inq_ary[4][31] ,
         \inq_ary[4][30] , \inq_ary[4][29] , \inq_ary[4][28] ,
         \inq_ary[4][27] , \inq_ary[4][26] , \inq_ary[4][25] ,
         \inq_ary[4][24] , \inq_ary[4][23] , \inq_ary[4][22] ,
         \inq_ary[4][21] , \inq_ary[4][20] , \inq_ary[4][19] ,
         \inq_ary[4][18] , \inq_ary[4][17] , \inq_ary[4][16] ,
         \inq_ary[4][15] , \inq_ary[4][14] , \inq_ary[4][13] ,
         \inq_ary[4][12] , \inq_ary[4][11] , \inq_ary[4][10] , \inq_ary[4][9] ,
         \inq_ary[4][8] , \inq_ary[4][7] , \inq_ary[4][6] , \inq_ary[4][5] ,
         \inq_ary[4][4] , \inq_ary[4][3] , \inq_ary[4][2] , \inq_ary[4][1] ,
         \inq_ary[4][0] , \inq_ary[3][159] , \inq_ary[3][158] ,
         \inq_ary[3][157] , \inq_ary[3][156] , \inq_ary[3][155] ,
         \inq_ary[3][154] , \inq_ary[3][153] , \inq_ary[3][152] ,
         \inq_ary[3][151] , \inq_ary[3][150] , \inq_ary[3][149] ,
         \inq_ary[3][148] , \inq_ary[3][147] , \inq_ary[3][146] ,
         \inq_ary[3][145] , \inq_ary[3][144] , \inq_ary[3][143] ,
         \inq_ary[3][142] , \inq_ary[3][141] , \inq_ary[3][140] ,
         \inq_ary[3][139] , \inq_ary[3][138] , \inq_ary[3][137] ,
         \inq_ary[3][136] , \inq_ary[3][135] , \inq_ary[3][134] ,
         \inq_ary[3][133] , \inq_ary[3][132] , \inq_ary[3][131] ,
         \inq_ary[3][130] , \inq_ary[3][129] , \inq_ary[3][128] ,
         \inq_ary[3][127] , \inq_ary[3][126] , \inq_ary[3][125] ,
         \inq_ary[3][124] , \inq_ary[3][123] , \inq_ary[3][122] ,
         \inq_ary[3][121] , \inq_ary[3][120] , \inq_ary[3][119] ,
         \inq_ary[3][118] , \inq_ary[3][117] , \inq_ary[3][116] ,
         \inq_ary[3][115] , \inq_ary[3][114] , \inq_ary[3][113] ,
         \inq_ary[3][112] , \inq_ary[3][111] , \inq_ary[3][110] ,
         \inq_ary[3][109] , \inq_ary[3][108] , \inq_ary[3][107] ,
         \inq_ary[3][106] , \inq_ary[3][105] , \inq_ary[3][104] ,
         \inq_ary[3][103] , \inq_ary[3][102] , \inq_ary[3][101] ,
         \inq_ary[3][100] , \inq_ary[3][99] , \inq_ary[3][98] ,
         \inq_ary[3][97] , \inq_ary[3][96] , \inq_ary[3][95] ,
         \inq_ary[3][94] , \inq_ary[3][93] , \inq_ary[3][92] ,
         \inq_ary[3][91] , \inq_ary[3][90] , \inq_ary[3][89] ,
         \inq_ary[3][88] , \inq_ary[3][87] , \inq_ary[3][86] ,
         \inq_ary[3][85] , \inq_ary[3][84] , \inq_ary[3][83] ,
         \inq_ary[3][82] , \inq_ary[3][81] , \inq_ary[3][80] ,
         \inq_ary[3][79] , \inq_ary[3][78] , \inq_ary[3][77] ,
         \inq_ary[3][76] , \inq_ary[3][75] , \inq_ary[3][74] ,
         \inq_ary[3][73] , \inq_ary[3][72] , \inq_ary[3][71] ,
         \inq_ary[3][70] , \inq_ary[3][69] , \inq_ary[3][68] ,
         \inq_ary[3][67] , \inq_ary[3][66] , \inq_ary[3][65] ,
         \inq_ary[3][64] , \inq_ary[3][63] , \inq_ary[3][62] ,
         \inq_ary[3][61] , \inq_ary[3][60] , \inq_ary[3][59] ,
         \inq_ary[3][58] , \inq_ary[3][57] , \inq_ary[3][56] ,
         \inq_ary[3][55] , \inq_ary[3][54] , \inq_ary[3][53] ,
         \inq_ary[3][52] , \inq_ary[3][51] , \inq_ary[3][50] ,
         \inq_ary[3][49] , \inq_ary[3][48] , \inq_ary[3][47] ,
         \inq_ary[3][46] , \inq_ary[3][45] , \inq_ary[3][44] ,
         \inq_ary[3][43] , \inq_ary[3][42] , \inq_ary[3][41] ,
         \inq_ary[3][40] , \inq_ary[3][39] , \inq_ary[3][38] ,
         \inq_ary[3][37] , \inq_ary[3][36] , \inq_ary[3][35] ,
         \inq_ary[3][34] , \inq_ary[3][33] , \inq_ary[3][32] ,
         \inq_ary[3][31] , \inq_ary[3][30] , \inq_ary[3][29] ,
         \inq_ary[3][28] , \inq_ary[3][27] , \inq_ary[3][26] ,
         \inq_ary[3][25] , \inq_ary[3][24] , \inq_ary[3][23] ,
         \inq_ary[3][22] , \inq_ary[3][21] , \inq_ary[3][20] ,
         \inq_ary[3][19] , \inq_ary[3][18] , \inq_ary[3][17] ,
         \inq_ary[3][16] , \inq_ary[3][15] , \inq_ary[3][14] ,
         \inq_ary[3][13] , \inq_ary[3][12] , \inq_ary[3][11] ,
         \inq_ary[3][10] , \inq_ary[3][9] , \inq_ary[3][8] , \inq_ary[3][7] ,
         \inq_ary[3][6] , \inq_ary[3][5] , \inq_ary[3][4] , \inq_ary[3][3] ,
         \inq_ary[3][2] , \inq_ary[3][1] , \inq_ary[3][0] , \inq_ary[2][159] ,
         \inq_ary[2][158] , \inq_ary[2][157] , \inq_ary[2][156] ,
         \inq_ary[2][155] , \inq_ary[2][154] , \inq_ary[2][153] ,
         \inq_ary[2][152] , \inq_ary[2][151] , \inq_ary[2][150] ,
         \inq_ary[2][149] , \inq_ary[2][148] , \inq_ary[2][147] ,
         \inq_ary[2][146] , \inq_ary[2][145] , \inq_ary[2][144] ,
         \inq_ary[2][143] , \inq_ary[2][142] , \inq_ary[2][141] ,
         \inq_ary[2][140] , \inq_ary[2][139] , \inq_ary[2][138] ,
         \inq_ary[2][137] , \inq_ary[2][136] , \inq_ary[2][135] ,
         \inq_ary[2][134] , \inq_ary[2][133] , \inq_ary[2][132] ,
         \inq_ary[2][131] , \inq_ary[2][130] , \inq_ary[2][129] ,
         \inq_ary[2][128] , \inq_ary[2][127] , \inq_ary[2][126] ,
         \inq_ary[2][125] , \inq_ary[2][124] , \inq_ary[2][123] ,
         \inq_ary[2][122] , \inq_ary[2][121] , \inq_ary[2][120] ,
         \inq_ary[2][119] , \inq_ary[2][118] , \inq_ary[2][117] ,
         \inq_ary[2][116] , \inq_ary[2][115] , \inq_ary[2][114] ,
         \inq_ary[2][113] , \inq_ary[2][112] , \inq_ary[2][111] ,
         \inq_ary[2][110] , \inq_ary[2][109] , \inq_ary[2][108] ,
         \inq_ary[2][107] , \inq_ary[2][106] , \inq_ary[2][105] ,
         \inq_ary[2][104] , \inq_ary[2][103] , \inq_ary[2][102] ,
         \inq_ary[2][101] , \inq_ary[2][100] , \inq_ary[2][99] ,
         \inq_ary[2][98] , \inq_ary[2][97] , \inq_ary[2][96] ,
         \inq_ary[2][95] , \inq_ary[2][94] , \inq_ary[2][93] ,
         \inq_ary[2][92] , \inq_ary[2][91] , \inq_ary[2][90] ,
         \inq_ary[2][89] , \inq_ary[2][88] , \inq_ary[2][87] ,
         \inq_ary[2][86] , \inq_ary[2][85] , \inq_ary[2][84] ,
         \inq_ary[2][83] , \inq_ary[2][82] , \inq_ary[2][81] ,
         \inq_ary[2][80] , \inq_ary[2][79] , \inq_ary[2][78] ,
         \inq_ary[2][77] , \inq_ary[2][76] , \inq_ary[2][75] ,
         \inq_ary[2][74] , \inq_ary[2][73] , \inq_ary[2][72] ,
         \inq_ary[2][71] , \inq_ary[2][70] , \inq_ary[2][69] ,
         \inq_ary[2][68] , \inq_ary[2][67] , \inq_ary[2][66] ,
         \inq_ary[2][65] , \inq_ary[2][64] , \inq_ary[2][63] ,
         \inq_ary[2][62] , \inq_ary[2][61] , \inq_ary[2][60] ,
         \inq_ary[2][59] , \inq_ary[2][58] , \inq_ary[2][57] ,
         \inq_ary[2][56] , \inq_ary[2][55] , \inq_ary[2][54] ,
         \inq_ary[2][53] , \inq_ary[2][52] , \inq_ary[2][51] ,
         \inq_ary[2][50] , \inq_ary[2][49] , \inq_ary[2][48] ,
         \inq_ary[2][47] , \inq_ary[2][46] , \inq_ary[2][45] ,
         \inq_ary[2][44] , \inq_ary[2][43] , \inq_ary[2][42] ,
         \inq_ary[2][41] , \inq_ary[2][40] , \inq_ary[2][39] ,
         \inq_ary[2][38] , \inq_ary[2][37] , \inq_ary[2][36] ,
         \inq_ary[2][35] , \inq_ary[2][34] , \inq_ary[2][33] ,
         \inq_ary[2][32] , \inq_ary[2][31] , \inq_ary[2][30] ,
         \inq_ary[2][29] , \inq_ary[2][28] , \inq_ary[2][27] ,
         \inq_ary[2][26] , \inq_ary[2][25] , \inq_ary[2][24] ,
         \inq_ary[2][23] , \inq_ary[2][22] , \inq_ary[2][21] ,
         \inq_ary[2][20] , \inq_ary[2][19] , \inq_ary[2][18] ,
         \inq_ary[2][17] , \inq_ary[2][16] , \inq_ary[2][15] ,
         \inq_ary[2][14] , \inq_ary[2][13] , \inq_ary[2][12] ,
         \inq_ary[2][11] , \inq_ary[2][10] , \inq_ary[2][9] , \inq_ary[2][8] ,
         \inq_ary[2][7] , \inq_ary[2][6] , \inq_ary[2][5] , \inq_ary[2][4] ,
         \inq_ary[2][3] , \inq_ary[2][2] , \inq_ary[2][1] , \inq_ary[2][0] ,
         \inq_ary[1][159] , \inq_ary[1][158] , \inq_ary[1][157] ,
         \inq_ary[1][156] , \inq_ary[1][155] , \inq_ary[1][154] ,
         \inq_ary[1][153] , \inq_ary[1][152] , \inq_ary[1][151] ,
         \inq_ary[1][150] , \inq_ary[1][149] , \inq_ary[1][148] ,
         \inq_ary[1][147] , \inq_ary[1][146] , \inq_ary[1][145] ,
         \inq_ary[1][144] , \inq_ary[1][143] , \inq_ary[1][142] ,
         \inq_ary[1][141] , \inq_ary[1][140] , \inq_ary[1][139] ,
         \inq_ary[1][138] , \inq_ary[1][137] , \inq_ary[1][136] ,
         \inq_ary[1][135] , \inq_ary[1][134] , \inq_ary[1][133] ,
         \inq_ary[1][132] , \inq_ary[1][131] , \inq_ary[1][130] ,
         \inq_ary[1][129] , \inq_ary[1][128] , \inq_ary[1][127] ,
         \inq_ary[1][126] , \inq_ary[1][125] , \inq_ary[1][124] ,
         \inq_ary[1][123] , \inq_ary[1][122] , \inq_ary[1][121] ,
         \inq_ary[1][120] , \inq_ary[1][119] , \inq_ary[1][118] ,
         \inq_ary[1][117] , \inq_ary[1][116] , \inq_ary[1][115] ,
         \inq_ary[1][114] , \inq_ary[1][113] , \inq_ary[1][112] ,
         \inq_ary[1][111] , \inq_ary[1][110] , \inq_ary[1][109] ,
         \inq_ary[1][108] , \inq_ary[1][107] , \inq_ary[1][106] ,
         \inq_ary[1][105] , \inq_ary[1][104] , \inq_ary[1][103] ,
         \inq_ary[1][102] , \inq_ary[1][101] , \inq_ary[1][100] ,
         \inq_ary[1][99] , \inq_ary[1][98] , \inq_ary[1][97] ,
         \inq_ary[1][96] , \inq_ary[1][95] , \inq_ary[1][94] ,
         \inq_ary[1][93] , \inq_ary[1][92] , \inq_ary[1][91] ,
         \inq_ary[1][90] , \inq_ary[1][89] , \inq_ary[1][88] ,
         \inq_ary[1][87] , \inq_ary[1][86] , \inq_ary[1][85] ,
         \inq_ary[1][84] , \inq_ary[1][83] , \inq_ary[1][82] ,
         \inq_ary[1][81] , \inq_ary[1][80] , \inq_ary[1][79] ,
         \inq_ary[1][78] , \inq_ary[1][77] , \inq_ary[1][76] ,
         \inq_ary[1][75] , \inq_ary[1][74] , \inq_ary[1][73] ,
         \inq_ary[1][72] , \inq_ary[1][71] , \inq_ary[1][70] ,
         \inq_ary[1][69] , \inq_ary[1][68] , \inq_ary[1][67] ,
         \inq_ary[1][66] , \inq_ary[1][65] , \inq_ary[1][64] ,
         \inq_ary[1][63] , \inq_ary[1][62] , \inq_ary[1][61] ,
         \inq_ary[1][60] , \inq_ary[1][59] , \inq_ary[1][58] ,
         \inq_ary[1][57] , \inq_ary[1][56] , \inq_ary[1][55] ,
         \inq_ary[1][54] , \inq_ary[1][53] , \inq_ary[1][52] ,
         \inq_ary[1][51] , \inq_ary[1][50] , \inq_ary[1][49] ,
         \inq_ary[1][48] , \inq_ary[1][47] , \inq_ary[1][46] ,
         \inq_ary[1][45] , \inq_ary[1][44] , \inq_ary[1][43] ,
         \inq_ary[1][42] , \inq_ary[1][41] , \inq_ary[1][40] ,
         \inq_ary[1][39] , \inq_ary[1][38] , \inq_ary[1][37] ,
         \inq_ary[1][36] , \inq_ary[1][35] , \inq_ary[1][34] ,
         \inq_ary[1][33] , \inq_ary[1][32] , \inq_ary[1][31] ,
         \inq_ary[1][30] , \inq_ary[1][29] , \inq_ary[1][28] ,
         \inq_ary[1][27] , \inq_ary[1][26] , \inq_ary[1][25] ,
         \inq_ary[1][24] , \inq_ary[1][23] , \inq_ary[1][22] ,
         \inq_ary[1][21] , \inq_ary[1][20] , \inq_ary[1][19] ,
         \inq_ary[1][18] , \inq_ary[1][17] , \inq_ary[1][16] ,
         \inq_ary[1][15] , \inq_ary[1][14] , \inq_ary[1][13] ,
         \inq_ary[1][12] , \inq_ary[1][11] , \inq_ary[1][10] , \inq_ary[1][9] ,
         \inq_ary[1][8] , \inq_ary[1][7] , \inq_ary[1][6] , \inq_ary[1][5] ,
         \inq_ary[1][4] , \inq_ary[1][3] , \inq_ary[1][2] , \inq_ary[1][1] ,
         \inq_ary[1][0] , \inq_ary[0][159] , \inq_ary[0][158] ,
         \inq_ary[0][157] , \inq_ary[0][156] , \inq_ary[0][155] ,
         \inq_ary[0][154] , \inq_ary[0][153] , \inq_ary[0][152] ,
         \inq_ary[0][151] , \inq_ary[0][150] , \inq_ary[0][149] ,
         \inq_ary[0][148] , \inq_ary[0][147] , \inq_ary[0][146] ,
         \inq_ary[0][145] , \inq_ary[0][144] , \inq_ary[0][143] ,
         \inq_ary[0][142] , \inq_ary[0][141] , \inq_ary[0][140] ,
         \inq_ary[0][139] , \inq_ary[0][138] , \inq_ary[0][137] ,
         \inq_ary[0][136] , \inq_ary[0][135] , \inq_ary[0][134] ,
         \inq_ary[0][133] , \inq_ary[0][132] , \inq_ary[0][131] ,
         \inq_ary[0][130] , \inq_ary[0][129] , \inq_ary[0][128] ,
         \inq_ary[0][127] , \inq_ary[0][126] , \inq_ary[0][125] ,
         \inq_ary[0][124] , \inq_ary[0][123] , \inq_ary[0][122] ,
         \inq_ary[0][121] , \inq_ary[0][120] , \inq_ary[0][119] ,
         \inq_ary[0][118] , \inq_ary[0][117] , \inq_ary[0][116] ,
         \inq_ary[0][115] , \inq_ary[0][114] , \inq_ary[0][113] ,
         \inq_ary[0][112] , \inq_ary[0][111] , \inq_ary[0][110] ,
         \inq_ary[0][109] , \inq_ary[0][108] , \inq_ary[0][107] ,
         \inq_ary[0][106] , \inq_ary[0][105] , \inq_ary[0][104] ,
         \inq_ary[0][103] , \inq_ary[0][102] , \inq_ary[0][101] ,
         \inq_ary[0][100] , \inq_ary[0][99] , \inq_ary[0][98] ,
         \inq_ary[0][97] , \inq_ary[0][96] , \inq_ary[0][95] ,
         \inq_ary[0][94] , \inq_ary[0][93] , \inq_ary[0][92] ,
         \inq_ary[0][91] , \inq_ary[0][90] , \inq_ary[0][89] ,
         \inq_ary[0][88] , \inq_ary[0][87] , \inq_ary[0][86] ,
         \inq_ary[0][85] , \inq_ary[0][84] , \inq_ary[0][83] ,
         \inq_ary[0][82] , \inq_ary[0][81] , \inq_ary[0][80] ,
         \inq_ary[0][79] , \inq_ary[0][78] , \inq_ary[0][77] ,
         \inq_ary[0][76] , \inq_ary[0][75] , \inq_ary[0][74] ,
         \inq_ary[0][73] , \inq_ary[0][72] , \inq_ary[0][71] ,
         \inq_ary[0][70] , \inq_ary[0][69] , \inq_ary[0][68] ,
         \inq_ary[0][67] , \inq_ary[0][66] , \inq_ary[0][65] ,
         \inq_ary[0][64] , \inq_ary[0][63] , \inq_ary[0][62] ,
         \inq_ary[0][61] , \inq_ary[0][60] , \inq_ary[0][59] ,
         \inq_ary[0][58] , \inq_ary[0][57] , \inq_ary[0][56] ,
         \inq_ary[0][55] , \inq_ary[0][54] , \inq_ary[0][53] ,
         \inq_ary[0][52] , \inq_ary[0][51] , \inq_ary[0][50] ,
         \inq_ary[0][49] , \inq_ary[0][48] , \inq_ary[0][47] ,
         \inq_ary[0][46] , \inq_ary[0][45] , \inq_ary[0][44] ,
         \inq_ary[0][43] , \inq_ary[0][42] , \inq_ary[0][41] ,
         \inq_ary[0][40] , \inq_ary[0][39] , \inq_ary[0][38] ,
         \inq_ary[0][37] , \inq_ary[0][36] , \inq_ary[0][35] ,
         \inq_ary[0][34] , \inq_ary[0][33] , \inq_ary[0][32] ,
         \inq_ary[0][31] , \inq_ary[0][30] , \inq_ary[0][29] ,
         \inq_ary[0][28] , \inq_ary[0][27] , \inq_ary[0][26] ,
         \inq_ary[0][25] , \inq_ary[0][24] , \inq_ary[0][23] ,
         \inq_ary[0][22] , \inq_ary[0][21] , \inq_ary[0][20] ,
         \inq_ary[0][19] , \inq_ary[0][18] , \inq_ary[0][17] ,
         \inq_ary[0][16] , \inq_ary[0][15] , \inq_ary[0][14] ,
         \inq_ary[0][13] , \inq_ary[0][12] , \inq_ary[0][11] ,
         \inq_ary[0][10] , \inq_ary[0][9] , \inq_ary[0][8] , \inq_ary[0][7] ,
         \inq_ary[0][6] , \inq_ary[0][5] , \inq_ary[0][4] , \inq_ary[0][3] ,
         \inq_ary[0][2] , \inq_ary[0][1] , \inq_ary[0][0] , N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, net16761, net16762;
  wire   [159:0] wrdata_d1;
  wire   [3:0] word_wen_d1;
  wire   [19:0] byte_wen_d1;
  wire   [3:0] wrptr_d1;
  wire   [3:0] rdptr_d1;

  \**SEQGEN**  \byte_wen_d1_reg[19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[19]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[19]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[18]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[18]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[17]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[17]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[16]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[16]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[15]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[15]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[14]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[14]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[13]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[13]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[12]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[12]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[11]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[11]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[10]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[10]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[9]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[9]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[8]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[8]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[7]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[7]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[6]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[6]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[5]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[5]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[4]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[4]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[3]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[2]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[1]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \byte_wen_d1_reg[0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(byte_wen[0]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(byte_wen_d1[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrptr_d1_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        wr_adr[3]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrptr_d1[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrptr_d1_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        wr_adr[2]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrptr_d1[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrptr_d1_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        wr_adr[1]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrptr_d1[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrptr_d1_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        wr_adr[0]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrptr_d1[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \word_wen_d1_reg[3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(word_wen[3]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(word_wen_d1[3]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \word_wen_d1_reg[2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(word_wen[2]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(word_wen_d1[2]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \word_wen_d1_reg[1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(word_wen[1]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(word_wen_d1[1]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \word_wen_d1_reg[0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(word_wen[0]), .clocked_on(wr_clk), .data_in(1'b0), 
        .enable(1'b0), .Q(word_wen_d1[0]), .synch_clear(1'b0), .synch_preset(
        1'b0), .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[159]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[159]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[158]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[158]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[157]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[157]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[156]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[156]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[155]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[155]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[154]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[154]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[153]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[153]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[152]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[152]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[151]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[151]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[150]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[150]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[149]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[149]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[148]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[148]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[147]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[147]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[146]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[146]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[145]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[145]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[144]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[144]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[143]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[143]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[142]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[142]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[141]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[141]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[140]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[140]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[139]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[139]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[138]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[138]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[137]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[137]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[136]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[136]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[135]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[135]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[134]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[134]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[133]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[133]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[132]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[132]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[131]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[131]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[130]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[130]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[129]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[129]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[128]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[128]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[127]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[127]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[126]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[126]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[125]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[125]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[124]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[124]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[123]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[123]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[122]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[122]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[121]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[121]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[120]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[120]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[119]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[119]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[118]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[118]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[117]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[117]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[116]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[116]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[115]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[115]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[114]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[114]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[113]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[113]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[112]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[112]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[111]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[111]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[110]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[110]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[109]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[109]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[108]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[108]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[107]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[107]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[106]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[106]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[105]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[105]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[104]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[104]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[103]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[103]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[102]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[102]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[101]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[101]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(din[100]), .clocked_on(wr_clk), .data_in(1'b0), .enable(
        1'b0), .Q(wrdata_d1[100]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[99]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[99]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[99]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[98]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[98]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[98]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[97]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[97]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[97]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[96]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[96]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[95]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[95]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[94]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[94]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[93]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[93]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[92]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[92]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[91]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[91]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[90]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[90]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[89]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[89]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[88]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[88]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[87]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[87]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[86]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[86]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[85]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[85]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[84]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[84]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[83]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[83]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[82]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[82]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[81]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[81]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[80]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[80]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[79]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[79]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[78]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[78]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[77]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[77]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[76]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[76]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[75]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[75]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[74]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[74]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[73]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[73]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[72]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[72]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[71]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[71]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[70]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[70]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[69]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[69]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[68]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[68]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[67]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[67]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[66]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[66]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[65]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[65]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[64]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[64]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[63]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[63]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[62]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[62]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[61]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[61]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[60]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[60]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[59]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[59]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[58]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[58]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[57]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[57]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[56]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[56]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[55]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[55]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[54]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[54]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[53]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[53]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[52]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[52]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[51]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[51]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[50]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[50]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[49]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[49]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[48]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[48]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[47]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[47]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[46]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[46]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[45]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[45]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[44]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[44]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[43]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[43]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[42]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[42]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[41]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[41]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[40]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[40]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[39]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[39]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[38]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[38]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[37]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[37]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[36]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[36]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[35]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[35]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[34]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[34]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[33]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[33]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[32]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[32]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[31]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[31]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[30]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[30]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[29]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[29]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[28]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[28]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[27]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[27]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[26]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[26]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[25]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[25]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[24]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[24]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[23]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[23]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[22]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[22]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[21]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[21]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[20]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[20]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[19]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[19]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[18]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[18]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[17]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[17]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[16]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[16]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[15]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[15]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[14]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[14]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[13]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[13]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[12]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[12]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[11]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[11]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[10]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[10]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[9]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[8]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[7]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[6]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[5]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[4]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[3]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[2]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[1]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \wrdata_d1_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        din[0]), .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(
        wrdata_d1[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  wr_en_d1_reg ( .clear(1'b0), .preset(1'b0), .next_state(wr_en), 
        .clocked_on(wr_clk), .data_in(1'b0), .enable(1'b0), .Q(wr_en_d1), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N989) );
  \**SEQGEN**  \rdptr_d1_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        rd_adr[3]), .clocked_on(rd_clk), .data_in(1'b0), .enable(1'b0), .Q(
        rdptr_d1[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \rdptr_d1_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        rd_adr[2]), .clocked_on(rd_clk), .data_in(1'b0), .enable(1'b0), .Q(
        rdptr_d1[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \rdptr_d1_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        rd_adr[1]), .clocked_on(rd_clk), .data_in(1'b0), .enable(1'b0), .Q(
        rdptr_d1[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  \rdptr_d1_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        rd_adr[0]), .clocked_on(rd_clk), .data_in(1'b0), .enable(1'b0), .Q(
        rdptr_d1[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(N989) );
  \**SEQGEN**  ren_d1_reg ( .clear(1'b0), .preset(1'b0), .next_state(read_en), 
        .clocked_on(rd_clk), .data_in(1'b0), .enable(1'b0), .Q(ren_d1), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N989) );
  \**SEQGEN**  \dout_reg[159]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N421), .enable(N360), .Q(dout[159]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[158]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N420), .enable(N360), .Q(dout[158]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[157]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N419), .enable(N360), .Q(dout[157]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[156]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N418), .enable(N360), .Q(dout[156]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[155]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N417), .enable(N360), .Q(dout[155]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[154]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N416), .enable(N360), .Q(dout[154]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[153]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N415), .enable(N360), .Q(dout[153]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[152]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N414), .enable(N360), .Q(dout[152]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[151]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N413), .enable(N360), .Q(dout[151]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[150]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N412), .enable(N360), .Q(dout[150]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[149]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N411), .enable(N360), .Q(dout[149]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[148]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N410), .enable(N360), .Q(dout[148]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[147]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N409), .enable(N360), .Q(dout[147]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[146]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N408), .enable(N360), .Q(dout[146]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[145]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N407), .enable(N360), .Q(dout[145]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[144]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N406), .enable(N360), .Q(dout[144]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[143]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N405), .enable(N360), .Q(dout[143]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[142]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N404), .enable(N360), .Q(dout[142]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[141]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N403), .enable(N360), .Q(dout[141]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[140]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N402), .enable(N360), .Q(dout[140]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[139]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N401), .enable(N360), .Q(dout[139]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[138]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N400), .enable(N360), .Q(dout[138]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[137]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N399), .enable(N360), .Q(dout[137]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[136]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N398), .enable(N360), .Q(dout[136]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[135]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N397), .enable(N360), .Q(dout[135]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[134]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N396), .enable(N360), .Q(dout[134]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[133]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N395), .enable(N360), .Q(dout[133]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[132]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N394), .enable(N360), .Q(dout[132]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[131]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N393), .enable(N360), .Q(dout[131]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[130]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N392), .enable(N360), .Q(dout[130]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[129]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N391), .enable(N360), .Q(dout[129]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[128]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N390), .enable(N360), .Q(dout[128]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[127]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N389), .enable(N360), .Q(dout[127]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[126]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N388), .enable(N360), .Q(dout[126]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[125]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N387), .enable(N360), .Q(dout[125]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[124]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N386), .enable(N360), .Q(dout[124]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[123]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N385), .enable(N360), .Q(dout[123]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[122]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N384), .enable(N360), .Q(dout[122]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[121]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N383), .enable(N360), .Q(dout[121]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[120]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N382), .enable(N360), .Q(dout[120]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[119]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N381), .enable(N360), .Q(dout[119]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[118]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N380), .enable(N360), .Q(dout[118]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[117]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N379), .enable(N360), .Q(dout[117]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[116]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N378), .enable(N360), .Q(dout[116]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[115]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N377), .enable(N360), .Q(dout[115]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[114]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N376), .enable(N360), .Q(dout[114]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[113]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N375), .enable(N360), .Q(dout[113]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[112]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N374), .enable(N360), .Q(dout[112]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[111]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N373), .enable(N360), .Q(dout[111]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[110]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N372), .enable(N360), .Q(dout[110]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[109]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N371), .enable(N360), .Q(dout[109]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[108]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N370), .enable(N360), .Q(dout[108]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[107]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N369), .enable(N360), .Q(dout[107]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[106]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N368), .enable(N360), .Q(dout[106]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[105]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N367), .enable(N360), .Q(dout[105]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[104]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N366), .enable(N360), .Q(dout[104]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[103]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N365), .enable(N360), .Q(dout[103]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[102]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N364), .enable(N360), .Q(dout[102]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[101]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N363), .enable(N360), .Q(dout[101]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[100]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), .clocked_on(1'b0), .data_in(N362), .enable(N360), .Q(dout[100]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[99]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N361), .enable(N360), .Q(dout[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[98]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N359), .enable(N260), .Q(dout[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[97]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N358), .enable(N260), .Q(dout[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N357), .enable(N260), .Q(dout[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N356), .enable(N260), .Q(dout[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N355), .enable(N260), .Q(dout[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N354), .enable(N260), .Q(dout[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N353), .enable(N260), .Q(dout[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N352), .enable(N260), .Q(dout[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N351), .enable(N260), .Q(dout[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N350), .enable(N260), .Q(dout[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N349), .enable(N260), .Q(dout[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N348), .enable(N260), .Q(dout[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N347), .enable(N260), .Q(dout[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N346), .enable(N260), .Q(dout[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N345), .enable(N260), .Q(dout[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N344), .enable(N260), .Q(dout[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N343), .enable(N260), .Q(dout[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N342), .enable(N260), .Q(dout[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N341), .enable(N260), .Q(dout[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N340), .enable(N260), .Q(dout[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N339), .enable(N260), .Q(dout[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N338), .enable(N260), .Q(dout[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N337), .enable(N260), .Q(dout[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N336), .enable(N260), .Q(dout[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N335), .enable(N260), .Q(dout[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N334), .enable(N260), .Q(dout[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N333), .enable(N260), .Q(dout[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N332), .enable(N260), .Q(dout[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N331), .enable(N260), .Q(dout[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N330), .enable(N260), .Q(dout[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N329), .enable(N260), .Q(dout[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N328), .enable(N260), .Q(dout[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N327), .enable(N260), .Q(dout[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N326), .enable(N260), .Q(dout[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N325), .enable(N260), .Q(dout[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N324), .enable(N260), .Q(dout[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N323), .enable(N260), .Q(dout[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N322), .enable(N260), .Q(dout[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N321), .enable(N260), .Q(dout[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N320), .enable(N260), .Q(dout[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N319), .enable(N260), .Q(dout[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N318), .enable(N260), .Q(dout[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N317), .enable(N260), .Q(dout[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N316), .enable(N260), .Q(dout[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N315), .enable(N260), .Q(dout[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N314), .enable(N260), .Q(dout[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N313), .enable(N260), .Q(dout[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N312), .enable(N260), .Q(dout[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N311), .enable(N260), .Q(dout[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N310), .enable(N260), .Q(dout[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N309), .enable(N260), .Q(dout[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N308), .enable(N260), .Q(dout[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N307), .enable(N260), .Q(dout[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N306), .enable(N260), .Q(dout[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N305), .enable(N260), .Q(dout[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N304), .enable(N260), .Q(dout[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N303), .enable(N260), .Q(dout[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N302), .enable(N260), .Q(dout[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N301), .enable(N260), .Q(dout[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N300), .enable(N260), .Q(dout[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N299), .enable(N260), .Q(dout[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N298), .enable(N260), .Q(dout[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N297), .enable(N260), .Q(dout[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N296), .enable(N260), .Q(dout[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N295), .enable(N260), .Q(dout[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N294), .enable(N260), .Q(dout[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N293), .enable(N260), .Q(dout[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N292), .enable(N260), .Q(dout[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N291), .enable(N260), .Q(dout[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N290), .enable(N260), .Q(dout[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N289), .enable(N260), .Q(dout[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N288), .enable(N260), .Q(dout[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N287), .enable(N260), .Q(dout[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N286), .enable(N260), .Q(dout[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N285), .enable(N260), .Q(dout[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N284), .enable(N260), .Q(dout[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N283), .enable(N260), .Q(dout[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N282), .enable(N260), .Q(dout[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N281), .enable(N260), .Q(dout[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N280), .enable(N260), .Q(dout[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N279), .enable(N260), .Q(dout[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N278), .enable(N260), .Q(dout[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N277), .enable(N260), .Q(dout[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N276), .enable(N260), .Q(dout[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N275), .enable(N260), .Q(dout[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N274), .enable(N260), .Q(dout[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N273), .enable(N260), .Q(dout[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N272), .enable(N260), .Q(dout[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N271), .enable(N260), .Q(dout[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N270), .enable(N260), .Q(dout[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N269), .enable(N260), .Q(dout[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N268), .enable(N260), .Q(dout[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N267), .enable(N260), .Q(dout[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N266), .enable(N260), .Q(dout[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N265), .enable(N260), .Q(dout[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N264), .enable(N260), .Q(dout[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N263), .enable(N260), .Q(dout[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N262), .enable(N260), .Q(dout[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \dout_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N261), .enable(N260), .Q(dout[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N988), 
        .Q(\inq_ary[15][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N988), 
        .Q(\inq_ary[15][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N988), 
        .Q(\inq_ary[15][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N988), 
        .Q(\inq_ary[15][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N988), 
        .Q(\inq_ary[15][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N988), 
        .Q(\inq_ary[15][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N988), 
        .Q(\inq_ary[15][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N988), 
        .Q(\inq_ary[15][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N988), 
        .Q(\inq_ary[15][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N988), 
        .Q(\inq_ary[15][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N988), 
        .Q(\inq_ary[15][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N988), 
        .Q(\inq_ary[15][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N988), 
        .Q(\inq_ary[15][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N988), 
        .Q(\inq_ary[15][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N988), 
        .Q(\inq_ary[15][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N988), 
        .Q(\inq_ary[15][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N988), 
        .Q(\inq_ary[15][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N988), 
        .Q(\inq_ary[15][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N988), 
        .Q(\inq_ary[15][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N988), 
        .Q(\inq_ary[15][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N988), 
        .Q(\inq_ary[15][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N988), 
        .Q(\inq_ary[15][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N988), 
        .Q(\inq_ary[15][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N988), 
        .Q(\inq_ary[15][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N988), 
        .Q(\inq_ary[15][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N988), 
        .Q(\inq_ary[15][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N988), 
        .Q(\inq_ary[15][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N988), 
        .Q(\inq_ary[15][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N988), 
        .Q(\inq_ary[15][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N988), 
        .Q(\inq_ary[15][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N988), 
        .Q(\inq_ary[15][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N988), 
        .Q(\inq_ary[15][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N988), 
        .Q(\inq_ary[15][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N988), 
        .Q(\inq_ary[15][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N988), 
        .Q(\inq_ary[15][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N988), 
        .Q(\inq_ary[15][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N988), 
        .Q(\inq_ary[15][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N988), 
        .Q(\inq_ary[15][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N988), 
        .Q(\inq_ary[15][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N988), 
        .Q(\inq_ary[15][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N988), 
        .Q(\inq_ary[15][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N988), 
        .Q(\inq_ary[15][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N988), 
        .Q(\inq_ary[15][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N988), 
        .Q(\inq_ary[15][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N988), 
        .Q(\inq_ary[15][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N988), 
        .Q(\inq_ary[15][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N988), 
        .Q(\inq_ary[15][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N988), 
        .Q(\inq_ary[15][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N988), 
        .Q(\inq_ary[15][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N988), 
        .Q(\inq_ary[15][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N988), 
        .Q(\inq_ary[15][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N988), 
        .Q(\inq_ary[15][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N988), 
        .Q(\inq_ary[15][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N988), 
        .Q(\inq_ary[15][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N988), 
        .Q(\inq_ary[15][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N988), 
        .Q(\inq_ary[15][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N988), 
        .Q(\inq_ary[15][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N988), 
        .Q(\inq_ary[15][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N988), 
        .Q(\inq_ary[15][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N988), 
        .Q(\inq_ary[15][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N988), 
        .Q(\inq_ary[15][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N987), 
        .Q(\inq_ary[15][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N987), 
        .Q(\inq_ary[15][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N987), 
        .Q(\inq_ary[15][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N987), 
        .Q(\inq_ary[15][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N987), 
        .Q(\inq_ary[15][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N987), 
        .Q(\inq_ary[15][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N987), 
        .Q(\inq_ary[15][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N987), 
        .Q(\inq_ary[15][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N987), 
        .Q(\inq_ary[15][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N987), 
        .Q(\inq_ary[15][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N987), 
        .Q(\inq_ary[15][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N987), 
        .Q(\inq_ary[15][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N987), 
        .Q(\inq_ary[15][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N987), 
        .Q(\inq_ary[15][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N987), 
        .Q(\inq_ary[15][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N987), 
        .Q(\inq_ary[15][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N987), 
        .Q(\inq_ary[15][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N987), 
        .Q(\inq_ary[15][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N987), 
        .Q(\inq_ary[15][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N987), 
        .Q(\inq_ary[15][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N987), 
        .Q(\inq_ary[15][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N987), 
        .Q(\inq_ary[15][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N987), 
        .Q(\inq_ary[15][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N987), 
        .Q(\inq_ary[15][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N987), 
        .Q(\inq_ary[15][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N987), 
        .Q(\inq_ary[15][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N987), 
        .Q(\inq_ary[15][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N987), 
        .Q(\inq_ary[15][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N987), 
        .Q(\inq_ary[15][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N987), 
        .Q(\inq_ary[15][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N987), 
        .Q(\inq_ary[15][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N987), 
        .Q(\inq_ary[15][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N987), 
        .Q(\inq_ary[15][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N987), 
        .Q(\inq_ary[15][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N987), 
        .Q(\inq_ary[15][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N987), 
        .Q(\inq_ary[15][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N987), 
        .Q(\inq_ary[15][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N987), 
        .Q(\inq_ary[15][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N987), 
        .Q(\inq_ary[15][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N987), 
        .Q(\inq_ary[15][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N987), 
        .Q(\inq_ary[15][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N987), 
        .Q(\inq_ary[15][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N987), 
        .Q(\inq_ary[15][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N987), 
        .Q(\inq_ary[15][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N987), 
        .Q(\inq_ary[15][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N987), 
        .Q(\inq_ary[15][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N987), 
        .Q(\inq_ary[15][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N987), 
        .Q(\inq_ary[15][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N987), 
        .Q(\inq_ary[15][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N987), 
        .Q(\inq_ary[15][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N987), 
        .Q(\inq_ary[15][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N987), 
        .Q(\inq_ary[15][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N987), 
        .Q(\inq_ary[15][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N987), 
        .Q(\inq_ary[15][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N987), 
        .Q(\inq_ary[15][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N987), 
        .Q(\inq_ary[15][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N987), 
        .Q(\inq_ary[15][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N987), 
        .Q(\inq_ary[15][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N987), 
        .Q(\inq_ary[15][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N987), 
        .Q(\inq_ary[15][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N987), 
        .Q(\inq_ary[15][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N987), 
        .Q(\inq_ary[15][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N987), 
        .Q(\inq_ary[15][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N987), 
        .Q(\inq_ary[15][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N987), 
        .Q(\inq_ary[15][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N987), 
        .Q(\inq_ary[15][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N987), 
        .Q(\inq_ary[15][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N987), 
        .Q(\inq_ary[15][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N987), 
        .Q(\inq_ary[15][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N987), 
        .Q(\inq_ary[15][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N987), 
        .Q(\inq_ary[15][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N987), 
        .Q(\inq_ary[15][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N987), 
        .Q(\inq_ary[15][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N987), 
        .Q(\inq_ary[15][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N987), 
        .Q(\inq_ary[15][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N987), 
        .Q(\inq_ary[15][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N987), 
        .Q(\inq_ary[15][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N987), 
        .Q(\inq_ary[15][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N987), 
        .Q(\inq_ary[15][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N987), 
        .Q(\inq_ary[15][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N987), 
        .Q(\inq_ary[15][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N987), 
        .Q(\inq_ary[15][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N987), 
        .Q(\inq_ary[15][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N987), 
        .Q(\inq_ary[15][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N987), 
        .Q(\inq_ary[15][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N987), 
        .Q(\inq_ary[15][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N987), 
        .Q(\inq_ary[15][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N987), 
        .Q(\inq_ary[15][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N987), 
        .Q(\inq_ary[15][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N987), 
        .Q(\inq_ary[15][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N987), 
        .Q(\inq_ary[15][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N987), 
        .Q(\inq_ary[15][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N987), 
        .Q(\inq_ary[15][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N987), 
        .Q(\inq_ary[15][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N987), 
        .Q(\inq_ary[15][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N987), 
        .Q(\inq_ary[15][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N987), 
        .Q(\inq_ary[15][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N987), 
        .Q(\inq_ary[15][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[15][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N987), 
        .Q(\inq_ary[15][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N986), 
        .Q(\inq_ary[14][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N986), 
        .Q(\inq_ary[14][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N986), 
        .Q(\inq_ary[14][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N986), 
        .Q(\inq_ary[14][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N986), 
        .Q(\inq_ary[14][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N986), 
        .Q(\inq_ary[14][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N986), 
        .Q(\inq_ary[14][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N986), 
        .Q(\inq_ary[14][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N986), 
        .Q(\inq_ary[14][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N986), 
        .Q(\inq_ary[14][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N986), 
        .Q(\inq_ary[14][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N986), 
        .Q(\inq_ary[14][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N986), 
        .Q(\inq_ary[14][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N986), 
        .Q(\inq_ary[14][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N986), 
        .Q(\inq_ary[14][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N986), 
        .Q(\inq_ary[14][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N986), 
        .Q(\inq_ary[14][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N986), 
        .Q(\inq_ary[14][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N986), 
        .Q(\inq_ary[14][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N986), 
        .Q(\inq_ary[14][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N986), 
        .Q(\inq_ary[14][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N986), 
        .Q(\inq_ary[14][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N986), 
        .Q(\inq_ary[14][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N986), 
        .Q(\inq_ary[14][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N986), 
        .Q(\inq_ary[14][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N986), 
        .Q(\inq_ary[14][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N986), 
        .Q(\inq_ary[14][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N986), 
        .Q(\inq_ary[14][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N986), 
        .Q(\inq_ary[14][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N986), 
        .Q(\inq_ary[14][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N986), 
        .Q(\inq_ary[14][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N986), 
        .Q(\inq_ary[14][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N986), 
        .Q(\inq_ary[14][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N986), 
        .Q(\inq_ary[14][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N986), 
        .Q(\inq_ary[14][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N986), 
        .Q(\inq_ary[14][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N986), 
        .Q(\inq_ary[14][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N986), 
        .Q(\inq_ary[14][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N986), 
        .Q(\inq_ary[14][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N986), 
        .Q(\inq_ary[14][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N986), 
        .Q(\inq_ary[14][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N986), 
        .Q(\inq_ary[14][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N986), 
        .Q(\inq_ary[14][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N986), 
        .Q(\inq_ary[14][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N986), 
        .Q(\inq_ary[14][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N986), 
        .Q(\inq_ary[14][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N986), 
        .Q(\inq_ary[14][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N986), 
        .Q(\inq_ary[14][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N986), 
        .Q(\inq_ary[14][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N986), 
        .Q(\inq_ary[14][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N986), 
        .Q(\inq_ary[14][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N986), 
        .Q(\inq_ary[14][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N986), 
        .Q(\inq_ary[14][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N986), 
        .Q(\inq_ary[14][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N986), 
        .Q(\inq_ary[14][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N986), 
        .Q(\inq_ary[14][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N986), 
        .Q(\inq_ary[14][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N986), 
        .Q(\inq_ary[14][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N986), 
        .Q(\inq_ary[14][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N986), 
        .Q(\inq_ary[14][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N986), 
        .Q(\inq_ary[14][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N985), 
        .Q(\inq_ary[14][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N985), 
        .Q(\inq_ary[14][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N985), 
        .Q(\inq_ary[14][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N985), 
        .Q(\inq_ary[14][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N985), 
        .Q(\inq_ary[14][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N985), 
        .Q(\inq_ary[14][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N985), 
        .Q(\inq_ary[14][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N985), 
        .Q(\inq_ary[14][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N985), 
        .Q(\inq_ary[14][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N985), 
        .Q(\inq_ary[14][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N985), 
        .Q(\inq_ary[14][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N985), 
        .Q(\inq_ary[14][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N985), 
        .Q(\inq_ary[14][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N985), 
        .Q(\inq_ary[14][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N985), 
        .Q(\inq_ary[14][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N985), 
        .Q(\inq_ary[14][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N985), 
        .Q(\inq_ary[14][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N985), 
        .Q(\inq_ary[14][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N985), 
        .Q(\inq_ary[14][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N985), 
        .Q(\inq_ary[14][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N985), 
        .Q(\inq_ary[14][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N985), 
        .Q(\inq_ary[14][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N985), 
        .Q(\inq_ary[14][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N985), 
        .Q(\inq_ary[14][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N985), 
        .Q(\inq_ary[14][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N985), 
        .Q(\inq_ary[14][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N985), 
        .Q(\inq_ary[14][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N985), 
        .Q(\inq_ary[14][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N985), 
        .Q(\inq_ary[14][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N985), 
        .Q(\inq_ary[14][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N985), 
        .Q(\inq_ary[14][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N985), 
        .Q(\inq_ary[14][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N985), 
        .Q(\inq_ary[14][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N985), 
        .Q(\inq_ary[14][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N985), 
        .Q(\inq_ary[14][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N985), 
        .Q(\inq_ary[14][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N985), 
        .Q(\inq_ary[14][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N985), 
        .Q(\inq_ary[14][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N985), 
        .Q(\inq_ary[14][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N985), 
        .Q(\inq_ary[14][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N985), 
        .Q(\inq_ary[14][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N985), 
        .Q(\inq_ary[14][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N985), 
        .Q(\inq_ary[14][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N985), 
        .Q(\inq_ary[14][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N985), 
        .Q(\inq_ary[14][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N985), 
        .Q(\inq_ary[14][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N985), 
        .Q(\inq_ary[14][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N985), 
        .Q(\inq_ary[14][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N985), 
        .Q(\inq_ary[14][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N985), 
        .Q(\inq_ary[14][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N985), 
        .Q(\inq_ary[14][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N985), 
        .Q(\inq_ary[14][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N985), 
        .Q(\inq_ary[14][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N985), 
        .Q(\inq_ary[14][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N985), 
        .Q(\inq_ary[14][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N985), 
        .Q(\inq_ary[14][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N985), 
        .Q(\inq_ary[14][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N985), 
        .Q(\inq_ary[14][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N985), 
        .Q(\inq_ary[14][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N985), 
        .Q(\inq_ary[14][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N985), 
        .Q(\inq_ary[14][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N985), 
        .Q(\inq_ary[14][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N985), 
        .Q(\inq_ary[14][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N985), 
        .Q(\inq_ary[14][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N985), 
        .Q(\inq_ary[14][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N985), 
        .Q(\inq_ary[14][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N985), 
        .Q(\inq_ary[14][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N985), 
        .Q(\inq_ary[14][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N985), 
        .Q(\inq_ary[14][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N985), 
        .Q(\inq_ary[14][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N985), 
        .Q(\inq_ary[14][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N985), 
        .Q(\inq_ary[14][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N985), 
        .Q(\inq_ary[14][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N985), 
        .Q(\inq_ary[14][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N985), 
        .Q(\inq_ary[14][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N985), 
        .Q(\inq_ary[14][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N985), 
        .Q(\inq_ary[14][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N985), 
        .Q(\inq_ary[14][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N985), 
        .Q(\inq_ary[14][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N985), 
        .Q(\inq_ary[14][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N985), 
        .Q(\inq_ary[14][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N985), 
        .Q(\inq_ary[14][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N985), 
        .Q(\inq_ary[14][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N985), 
        .Q(\inq_ary[14][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N985), 
        .Q(\inq_ary[14][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N985), 
        .Q(\inq_ary[14][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N985), 
        .Q(\inq_ary[14][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N985), 
        .Q(\inq_ary[14][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N985), 
        .Q(\inq_ary[14][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N985), 
        .Q(\inq_ary[14][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N985), 
        .Q(\inq_ary[14][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N985), 
        .Q(\inq_ary[14][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N985), 
        .Q(\inq_ary[14][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N985), 
        .Q(\inq_ary[14][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N985), 
        .Q(\inq_ary[14][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N985), 
        .Q(\inq_ary[14][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N985), 
        .Q(\inq_ary[14][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N985), 
        .Q(\inq_ary[14][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[14][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N985), 
        .Q(\inq_ary[14][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N984), 
        .Q(\inq_ary[13][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N984), 
        .Q(\inq_ary[13][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N984), 
        .Q(\inq_ary[13][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N984), 
        .Q(\inq_ary[13][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N984), 
        .Q(\inq_ary[13][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N984), 
        .Q(\inq_ary[13][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N984), 
        .Q(\inq_ary[13][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N984), 
        .Q(\inq_ary[13][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N984), 
        .Q(\inq_ary[13][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N984), 
        .Q(\inq_ary[13][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N984), 
        .Q(\inq_ary[13][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N984), 
        .Q(\inq_ary[13][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N984), 
        .Q(\inq_ary[13][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N984), 
        .Q(\inq_ary[13][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N984), 
        .Q(\inq_ary[13][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N984), 
        .Q(\inq_ary[13][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N984), 
        .Q(\inq_ary[13][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N984), 
        .Q(\inq_ary[13][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N984), 
        .Q(\inq_ary[13][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N984), 
        .Q(\inq_ary[13][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N984), 
        .Q(\inq_ary[13][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N984), 
        .Q(\inq_ary[13][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N984), 
        .Q(\inq_ary[13][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N984), 
        .Q(\inq_ary[13][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N984), 
        .Q(\inq_ary[13][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N984), 
        .Q(\inq_ary[13][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N984), 
        .Q(\inq_ary[13][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N984), 
        .Q(\inq_ary[13][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N984), 
        .Q(\inq_ary[13][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N984), 
        .Q(\inq_ary[13][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N984), 
        .Q(\inq_ary[13][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N984), 
        .Q(\inq_ary[13][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N984), 
        .Q(\inq_ary[13][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N984), 
        .Q(\inq_ary[13][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N984), 
        .Q(\inq_ary[13][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N984), 
        .Q(\inq_ary[13][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N984), 
        .Q(\inq_ary[13][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N984), 
        .Q(\inq_ary[13][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N984), 
        .Q(\inq_ary[13][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N984), 
        .Q(\inq_ary[13][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N984), 
        .Q(\inq_ary[13][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N984), 
        .Q(\inq_ary[13][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N984), 
        .Q(\inq_ary[13][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N984), 
        .Q(\inq_ary[13][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N984), 
        .Q(\inq_ary[13][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N984), 
        .Q(\inq_ary[13][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N984), 
        .Q(\inq_ary[13][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N984), 
        .Q(\inq_ary[13][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N984), 
        .Q(\inq_ary[13][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N984), 
        .Q(\inq_ary[13][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N984), 
        .Q(\inq_ary[13][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N984), 
        .Q(\inq_ary[13][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N984), 
        .Q(\inq_ary[13][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N984), 
        .Q(\inq_ary[13][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N984), 
        .Q(\inq_ary[13][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N984), 
        .Q(\inq_ary[13][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N984), 
        .Q(\inq_ary[13][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N984), 
        .Q(\inq_ary[13][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N984), 
        .Q(\inq_ary[13][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N984), 
        .Q(\inq_ary[13][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N984), 
        .Q(\inq_ary[13][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N983), 
        .Q(\inq_ary[13][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N983), 
        .Q(\inq_ary[13][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N983), 
        .Q(\inq_ary[13][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N983), 
        .Q(\inq_ary[13][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N983), 
        .Q(\inq_ary[13][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N983), 
        .Q(\inq_ary[13][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N983), 
        .Q(\inq_ary[13][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N983), 
        .Q(\inq_ary[13][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N983), 
        .Q(\inq_ary[13][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N983), 
        .Q(\inq_ary[13][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N983), 
        .Q(\inq_ary[13][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N983), 
        .Q(\inq_ary[13][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N983), 
        .Q(\inq_ary[13][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N983), 
        .Q(\inq_ary[13][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N983), 
        .Q(\inq_ary[13][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N983), 
        .Q(\inq_ary[13][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N983), 
        .Q(\inq_ary[13][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N983), 
        .Q(\inq_ary[13][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N983), 
        .Q(\inq_ary[13][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N983), 
        .Q(\inq_ary[13][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N983), 
        .Q(\inq_ary[13][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N983), 
        .Q(\inq_ary[13][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N983), 
        .Q(\inq_ary[13][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N983), 
        .Q(\inq_ary[13][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N983), 
        .Q(\inq_ary[13][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N983), 
        .Q(\inq_ary[13][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N983), 
        .Q(\inq_ary[13][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N983), 
        .Q(\inq_ary[13][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N983), 
        .Q(\inq_ary[13][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N983), 
        .Q(\inq_ary[13][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N983), 
        .Q(\inq_ary[13][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N983), 
        .Q(\inq_ary[13][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N983), 
        .Q(\inq_ary[13][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N983), 
        .Q(\inq_ary[13][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N983), 
        .Q(\inq_ary[13][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N983), 
        .Q(\inq_ary[13][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N983), 
        .Q(\inq_ary[13][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N983), 
        .Q(\inq_ary[13][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N983), 
        .Q(\inq_ary[13][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N983), 
        .Q(\inq_ary[13][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N983), 
        .Q(\inq_ary[13][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N983), 
        .Q(\inq_ary[13][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N983), 
        .Q(\inq_ary[13][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N983), 
        .Q(\inq_ary[13][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N983), 
        .Q(\inq_ary[13][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N983), 
        .Q(\inq_ary[13][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N983), 
        .Q(\inq_ary[13][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N983), 
        .Q(\inq_ary[13][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N983), 
        .Q(\inq_ary[13][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N983), 
        .Q(\inq_ary[13][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N983), 
        .Q(\inq_ary[13][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N983), 
        .Q(\inq_ary[13][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N983), 
        .Q(\inq_ary[13][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N983), 
        .Q(\inq_ary[13][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N983), 
        .Q(\inq_ary[13][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N983), 
        .Q(\inq_ary[13][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N983), 
        .Q(\inq_ary[13][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N983), 
        .Q(\inq_ary[13][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N983), 
        .Q(\inq_ary[13][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N983), 
        .Q(\inq_ary[13][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N983), 
        .Q(\inq_ary[13][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N983), 
        .Q(\inq_ary[13][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N983), 
        .Q(\inq_ary[13][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N983), 
        .Q(\inq_ary[13][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N983), 
        .Q(\inq_ary[13][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N983), 
        .Q(\inq_ary[13][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N983), 
        .Q(\inq_ary[13][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N983), 
        .Q(\inq_ary[13][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N983), 
        .Q(\inq_ary[13][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N983), 
        .Q(\inq_ary[13][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N983), 
        .Q(\inq_ary[13][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N983), 
        .Q(\inq_ary[13][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N983), 
        .Q(\inq_ary[13][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N983), 
        .Q(\inq_ary[13][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N983), 
        .Q(\inq_ary[13][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N983), 
        .Q(\inq_ary[13][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N983), 
        .Q(\inq_ary[13][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N983), 
        .Q(\inq_ary[13][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N983), 
        .Q(\inq_ary[13][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N983), 
        .Q(\inq_ary[13][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N983), 
        .Q(\inq_ary[13][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N983), 
        .Q(\inq_ary[13][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N983), 
        .Q(\inq_ary[13][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N983), 
        .Q(\inq_ary[13][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N983), 
        .Q(\inq_ary[13][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N983), 
        .Q(\inq_ary[13][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N983), 
        .Q(\inq_ary[13][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N983), 
        .Q(\inq_ary[13][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N983), 
        .Q(\inq_ary[13][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N983), 
        .Q(\inq_ary[13][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N983), 
        .Q(\inq_ary[13][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N983), 
        .Q(\inq_ary[13][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N983), 
        .Q(\inq_ary[13][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N983), 
        .Q(\inq_ary[13][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N983), 
        .Q(\inq_ary[13][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N983), 
        .Q(\inq_ary[13][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N983), 
        .Q(\inq_ary[13][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N983), 
        .Q(\inq_ary[13][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[13][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N983), 
        .Q(\inq_ary[13][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N982), 
        .Q(\inq_ary[12][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N982), 
        .Q(\inq_ary[12][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N982), 
        .Q(\inq_ary[12][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N982), 
        .Q(\inq_ary[12][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N982), 
        .Q(\inq_ary[12][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N982), 
        .Q(\inq_ary[12][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N982), 
        .Q(\inq_ary[12][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N982), 
        .Q(\inq_ary[12][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N982), 
        .Q(\inq_ary[12][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N982), 
        .Q(\inq_ary[12][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N982), 
        .Q(\inq_ary[12][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N982), 
        .Q(\inq_ary[12][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N982), 
        .Q(\inq_ary[12][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N982), 
        .Q(\inq_ary[12][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N982), 
        .Q(\inq_ary[12][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N982), 
        .Q(\inq_ary[12][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N982), 
        .Q(\inq_ary[12][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N982), 
        .Q(\inq_ary[12][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N982), 
        .Q(\inq_ary[12][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N982), 
        .Q(\inq_ary[12][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N982), 
        .Q(\inq_ary[12][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N982), 
        .Q(\inq_ary[12][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N982), 
        .Q(\inq_ary[12][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N982), 
        .Q(\inq_ary[12][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N982), 
        .Q(\inq_ary[12][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N982), 
        .Q(\inq_ary[12][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N982), 
        .Q(\inq_ary[12][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N982), 
        .Q(\inq_ary[12][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N982), 
        .Q(\inq_ary[12][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N982), 
        .Q(\inq_ary[12][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N982), 
        .Q(\inq_ary[12][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N982), 
        .Q(\inq_ary[12][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N982), 
        .Q(\inq_ary[12][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N982), 
        .Q(\inq_ary[12][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N982), 
        .Q(\inq_ary[12][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N982), 
        .Q(\inq_ary[12][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N982), 
        .Q(\inq_ary[12][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N982), 
        .Q(\inq_ary[12][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N982), 
        .Q(\inq_ary[12][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N982), 
        .Q(\inq_ary[12][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N982), 
        .Q(\inq_ary[12][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N982), 
        .Q(\inq_ary[12][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N982), 
        .Q(\inq_ary[12][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N982), 
        .Q(\inq_ary[12][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N982), 
        .Q(\inq_ary[12][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N982), 
        .Q(\inq_ary[12][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N982), 
        .Q(\inq_ary[12][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N982), 
        .Q(\inq_ary[12][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N982), 
        .Q(\inq_ary[12][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N982), 
        .Q(\inq_ary[12][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N982), 
        .Q(\inq_ary[12][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N982), 
        .Q(\inq_ary[12][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N982), 
        .Q(\inq_ary[12][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N982), 
        .Q(\inq_ary[12][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N982), 
        .Q(\inq_ary[12][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N982), 
        .Q(\inq_ary[12][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N982), 
        .Q(\inq_ary[12][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N982), 
        .Q(\inq_ary[12][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N982), 
        .Q(\inq_ary[12][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N982), 
        .Q(\inq_ary[12][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N982), 
        .Q(\inq_ary[12][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N981), 
        .Q(\inq_ary[12][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N981), 
        .Q(\inq_ary[12][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N981), 
        .Q(\inq_ary[12][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N981), 
        .Q(\inq_ary[12][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N981), 
        .Q(\inq_ary[12][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N981), 
        .Q(\inq_ary[12][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N981), 
        .Q(\inq_ary[12][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N981), 
        .Q(\inq_ary[12][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N981), 
        .Q(\inq_ary[12][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N981), 
        .Q(\inq_ary[12][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N981), 
        .Q(\inq_ary[12][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N981), 
        .Q(\inq_ary[12][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N981), 
        .Q(\inq_ary[12][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N981), 
        .Q(\inq_ary[12][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N981), 
        .Q(\inq_ary[12][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N981), 
        .Q(\inq_ary[12][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N981), 
        .Q(\inq_ary[12][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N981), 
        .Q(\inq_ary[12][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N981), 
        .Q(\inq_ary[12][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N981), 
        .Q(\inq_ary[12][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N981), 
        .Q(\inq_ary[12][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N981), 
        .Q(\inq_ary[12][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N981), 
        .Q(\inq_ary[12][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N981), 
        .Q(\inq_ary[12][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N981), 
        .Q(\inq_ary[12][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N981), 
        .Q(\inq_ary[12][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N981), 
        .Q(\inq_ary[12][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N981), 
        .Q(\inq_ary[12][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N981), 
        .Q(\inq_ary[12][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N981), 
        .Q(\inq_ary[12][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N981), 
        .Q(\inq_ary[12][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N981), 
        .Q(\inq_ary[12][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N981), 
        .Q(\inq_ary[12][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N981), 
        .Q(\inq_ary[12][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N981), 
        .Q(\inq_ary[12][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N981), 
        .Q(\inq_ary[12][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N981), 
        .Q(\inq_ary[12][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N981), 
        .Q(\inq_ary[12][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N981), 
        .Q(\inq_ary[12][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N981), 
        .Q(\inq_ary[12][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N981), 
        .Q(\inq_ary[12][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N981), 
        .Q(\inq_ary[12][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N981), 
        .Q(\inq_ary[12][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N981), 
        .Q(\inq_ary[12][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N981), 
        .Q(\inq_ary[12][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N981), 
        .Q(\inq_ary[12][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N981), 
        .Q(\inq_ary[12][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N981), 
        .Q(\inq_ary[12][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N981), 
        .Q(\inq_ary[12][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N981), 
        .Q(\inq_ary[12][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N981), 
        .Q(\inq_ary[12][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N981), 
        .Q(\inq_ary[12][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N981), 
        .Q(\inq_ary[12][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N981), 
        .Q(\inq_ary[12][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N981), 
        .Q(\inq_ary[12][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N981), 
        .Q(\inq_ary[12][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N981), 
        .Q(\inq_ary[12][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N981), 
        .Q(\inq_ary[12][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N981), 
        .Q(\inq_ary[12][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N981), 
        .Q(\inq_ary[12][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N981), 
        .Q(\inq_ary[12][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N981), 
        .Q(\inq_ary[12][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N981), 
        .Q(\inq_ary[12][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N981), 
        .Q(\inq_ary[12][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N981), 
        .Q(\inq_ary[12][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N981), 
        .Q(\inq_ary[12][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N981), 
        .Q(\inq_ary[12][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N981), 
        .Q(\inq_ary[12][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N981), 
        .Q(\inq_ary[12][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N981), 
        .Q(\inq_ary[12][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N981), 
        .Q(\inq_ary[12][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N981), 
        .Q(\inq_ary[12][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N981), 
        .Q(\inq_ary[12][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N981), 
        .Q(\inq_ary[12][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N981), 
        .Q(\inq_ary[12][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N981), 
        .Q(\inq_ary[12][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N981), 
        .Q(\inq_ary[12][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N981), 
        .Q(\inq_ary[12][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N981), 
        .Q(\inq_ary[12][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N981), 
        .Q(\inq_ary[12][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N981), 
        .Q(\inq_ary[12][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N981), 
        .Q(\inq_ary[12][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N981), 
        .Q(\inq_ary[12][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N981), 
        .Q(\inq_ary[12][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N981), 
        .Q(\inq_ary[12][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N981), 
        .Q(\inq_ary[12][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N981), 
        .Q(\inq_ary[12][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N981), 
        .Q(\inq_ary[12][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N981), 
        .Q(\inq_ary[12][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N981), 
        .Q(\inq_ary[12][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N981), 
        .Q(\inq_ary[12][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N981), 
        .Q(\inq_ary[12][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N981), 
        .Q(\inq_ary[12][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N981), 
        .Q(\inq_ary[12][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N981), 
        .Q(\inq_ary[12][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N981), 
        .Q(\inq_ary[12][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N981), 
        .Q(\inq_ary[12][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N981), 
        .Q(\inq_ary[12][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[12][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N981), 
        .Q(\inq_ary[12][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N980), 
        .Q(\inq_ary[11][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N980), 
        .Q(\inq_ary[11][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N980), 
        .Q(\inq_ary[11][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N980), 
        .Q(\inq_ary[11][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N980), 
        .Q(\inq_ary[11][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N980), 
        .Q(\inq_ary[11][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N980), 
        .Q(\inq_ary[11][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N980), 
        .Q(\inq_ary[11][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N980), 
        .Q(\inq_ary[11][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N980), 
        .Q(\inq_ary[11][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N980), 
        .Q(\inq_ary[11][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N980), 
        .Q(\inq_ary[11][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N980), 
        .Q(\inq_ary[11][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N980), 
        .Q(\inq_ary[11][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N980), 
        .Q(\inq_ary[11][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N980), 
        .Q(\inq_ary[11][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N980), 
        .Q(\inq_ary[11][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N980), 
        .Q(\inq_ary[11][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N980), 
        .Q(\inq_ary[11][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N980), 
        .Q(\inq_ary[11][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N980), 
        .Q(\inq_ary[11][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N980), 
        .Q(\inq_ary[11][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N980), 
        .Q(\inq_ary[11][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N980), 
        .Q(\inq_ary[11][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N980), 
        .Q(\inq_ary[11][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N980), 
        .Q(\inq_ary[11][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N980), 
        .Q(\inq_ary[11][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N980), 
        .Q(\inq_ary[11][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N980), 
        .Q(\inq_ary[11][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N980), 
        .Q(\inq_ary[11][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N980), 
        .Q(\inq_ary[11][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N980), 
        .Q(\inq_ary[11][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N980), 
        .Q(\inq_ary[11][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N980), 
        .Q(\inq_ary[11][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N980), 
        .Q(\inq_ary[11][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N980), 
        .Q(\inq_ary[11][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N980), 
        .Q(\inq_ary[11][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N980), 
        .Q(\inq_ary[11][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N980), 
        .Q(\inq_ary[11][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N980), 
        .Q(\inq_ary[11][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N980), 
        .Q(\inq_ary[11][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N980), 
        .Q(\inq_ary[11][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N980), 
        .Q(\inq_ary[11][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N980), 
        .Q(\inq_ary[11][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N980), 
        .Q(\inq_ary[11][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N980), 
        .Q(\inq_ary[11][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N980), 
        .Q(\inq_ary[11][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N980), 
        .Q(\inq_ary[11][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N980), 
        .Q(\inq_ary[11][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N980), 
        .Q(\inq_ary[11][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N980), 
        .Q(\inq_ary[11][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N980), 
        .Q(\inq_ary[11][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N980), 
        .Q(\inq_ary[11][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N980), 
        .Q(\inq_ary[11][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N980), 
        .Q(\inq_ary[11][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N980), 
        .Q(\inq_ary[11][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N980), 
        .Q(\inq_ary[11][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N980), 
        .Q(\inq_ary[11][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N980), 
        .Q(\inq_ary[11][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N980), 
        .Q(\inq_ary[11][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N980), 
        .Q(\inq_ary[11][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N979), 
        .Q(\inq_ary[11][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N979), 
        .Q(\inq_ary[11][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N979), 
        .Q(\inq_ary[11][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N979), 
        .Q(\inq_ary[11][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N979), 
        .Q(\inq_ary[11][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N979), 
        .Q(\inq_ary[11][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N979), 
        .Q(\inq_ary[11][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N979), 
        .Q(\inq_ary[11][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N979), 
        .Q(\inq_ary[11][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N979), 
        .Q(\inq_ary[11][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N979), 
        .Q(\inq_ary[11][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N979), 
        .Q(\inq_ary[11][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N979), 
        .Q(\inq_ary[11][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N979), 
        .Q(\inq_ary[11][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N979), 
        .Q(\inq_ary[11][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N979), 
        .Q(\inq_ary[11][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N979), 
        .Q(\inq_ary[11][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N979), 
        .Q(\inq_ary[11][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N979), 
        .Q(\inq_ary[11][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N979), 
        .Q(\inq_ary[11][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N979), 
        .Q(\inq_ary[11][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N979), 
        .Q(\inq_ary[11][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N979), 
        .Q(\inq_ary[11][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N979), 
        .Q(\inq_ary[11][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N979), 
        .Q(\inq_ary[11][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N979), 
        .Q(\inq_ary[11][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N979), 
        .Q(\inq_ary[11][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N979), 
        .Q(\inq_ary[11][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N979), 
        .Q(\inq_ary[11][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N979), 
        .Q(\inq_ary[11][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N979), 
        .Q(\inq_ary[11][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N979), 
        .Q(\inq_ary[11][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N979), 
        .Q(\inq_ary[11][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N979), 
        .Q(\inq_ary[11][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N979), 
        .Q(\inq_ary[11][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N979), 
        .Q(\inq_ary[11][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N979), 
        .Q(\inq_ary[11][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N979), 
        .Q(\inq_ary[11][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N979), 
        .Q(\inq_ary[11][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N979), 
        .Q(\inq_ary[11][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N979), 
        .Q(\inq_ary[11][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N979), 
        .Q(\inq_ary[11][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N979), 
        .Q(\inq_ary[11][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N979), 
        .Q(\inq_ary[11][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N979), 
        .Q(\inq_ary[11][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N979), 
        .Q(\inq_ary[11][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N979), 
        .Q(\inq_ary[11][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N979), 
        .Q(\inq_ary[11][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N979), 
        .Q(\inq_ary[11][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N979), 
        .Q(\inq_ary[11][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N979), 
        .Q(\inq_ary[11][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N979), 
        .Q(\inq_ary[11][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N979), 
        .Q(\inq_ary[11][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N979), 
        .Q(\inq_ary[11][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N979), 
        .Q(\inq_ary[11][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N979), 
        .Q(\inq_ary[11][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N979), 
        .Q(\inq_ary[11][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N979), 
        .Q(\inq_ary[11][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N979), 
        .Q(\inq_ary[11][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N979), 
        .Q(\inq_ary[11][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N979), 
        .Q(\inq_ary[11][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N979), 
        .Q(\inq_ary[11][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N979), 
        .Q(\inq_ary[11][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N979), 
        .Q(\inq_ary[11][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N979), 
        .Q(\inq_ary[11][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N979), 
        .Q(\inq_ary[11][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N979), 
        .Q(\inq_ary[11][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N979), 
        .Q(\inq_ary[11][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N979), 
        .Q(\inq_ary[11][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N979), 
        .Q(\inq_ary[11][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N979), 
        .Q(\inq_ary[11][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N979), 
        .Q(\inq_ary[11][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N979), 
        .Q(\inq_ary[11][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N979), 
        .Q(\inq_ary[11][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N979), 
        .Q(\inq_ary[11][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N979), 
        .Q(\inq_ary[11][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N979), 
        .Q(\inq_ary[11][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N979), 
        .Q(\inq_ary[11][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N979), 
        .Q(\inq_ary[11][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N979), 
        .Q(\inq_ary[11][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N979), 
        .Q(\inq_ary[11][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N979), 
        .Q(\inq_ary[11][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N979), 
        .Q(\inq_ary[11][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N979), 
        .Q(\inq_ary[11][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N979), 
        .Q(\inq_ary[11][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N979), 
        .Q(\inq_ary[11][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N979), 
        .Q(\inq_ary[11][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N979), 
        .Q(\inq_ary[11][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N979), 
        .Q(\inq_ary[11][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N979), 
        .Q(\inq_ary[11][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N979), 
        .Q(\inq_ary[11][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N979), 
        .Q(\inq_ary[11][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N979), 
        .Q(\inq_ary[11][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N979), 
        .Q(\inq_ary[11][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N979), 
        .Q(\inq_ary[11][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N979), 
        .Q(\inq_ary[11][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N979), 
        .Q(\inq_ary[11][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N979), 
        .Q(\inq_ary[11][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[11][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N979), 
        .Q(\inq_ary[11][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N978), 
        .Q(\inq_ary[10][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N978), 
        .Q(\inq_ary[10][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N978), 
        .Q(\inq_ary[10][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N978), 
        .Q(\inq_ary[10][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N978), 
        .Q(\inq_ary[10][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N978), 
        .Q(\inq_ary[10][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N978), 
        .Q(\inq_ary[10][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N978), 
        .Q(\inq_ary[10][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N978), 
        .Q(\inq_ary[10][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N978), 
        .Q(\inq_ary[10][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N978), 
        .Q(\inq_ary[10][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N978), 
        .Q(\inq_ary[10][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N978), 
        .Q(\inq_ary[10][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N978), 
        .Q(\inq_ary[10][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N978), 
        .Q(\inq_ary[10][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N978), 
        .Q(\inq_ary[10][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N978), 
        .Q(\inq_ary[10][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N978), 
        .Q(\inq_ary[10][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N978), 
        .Q(\inq_ary[10][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N978), 
        .Q(\inq_ary[10][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N978), 
        .Q(\inq_ary[10][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N978), 
        .Q(\inq_ary[10][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N978), 
        .Q(\inq_ary[10][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N978), 
        .Q(\inq_ary[10][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N978), 
        .Q(\inq_ary[10][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N978), 
        .Q(\inq_ary[10][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N978), 
        .Q(\inq_ary[10][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N978), 
        .Q(\inq_ary[10][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N978), 
        .Q(\inq_ary[10][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N978), 
        .Q(\inq_ary[10][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N978), 
        .Q(\inq_ary[10][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N978), 
        .Q(\inq_ary[10][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N978), 
        .Q(\inq_ary[10][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N978), 
        .Q(\inq_ary[10][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N978), 
        .Q(\inq_ary[10][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N978), 
        .Q(\inq_ary[10][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N978), 
        .Q(\inq_ary[10][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N978), 
        .Q(\inq_ary[10][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N978), 
        .Q(\inq_ary[10][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N978), 
        .Q(\inq_ary[10][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N978), 
        .Q(\inq_ary[10][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N978), 
        .Q(\inq_ary[10][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N978), 
        .Q(\inq_ary[10][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N978), 
        .Q(\inq_ary[10][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N978), 
        .Q(\inq_ary[10][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N978), 
        .Q(\inq_ary[10][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N978), 
        .Q(\inq_ary[10][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N978), 
        .Q(\inq_ary[10][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N978), 
        .Q(\inq_ary[10][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N978), 
        .Q(\inq_ary[10][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N978), 
        .Q(\inq_ary[10][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N978), 
        .Q(\inq_ary[10][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N978), 
        .Q(\inq_ary[10][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N978), 
        .Q(\inq_ary[10][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N978), 
        .Q(\inq_ary[10][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N978), 
        .Q(\inq_ary[10][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N978), 
        .Q(\inq_ary[10][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N978), 
        .Q(\inq_ary[10][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N978), 
        .Q(\inq_ary[10][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N978), 
        .Q(\inq_ary[10][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N978), 
        .Q(\inq_ary[10][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N977), 
        .Q(\inq_ary[10][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N977), 
        .Q(\inq_ary[10][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N977), 
        .Q(\inq_ary[10][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N977), 
        .Q(\inq_ary[10][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N977), 
        .Q(\inq_ary[10][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N977), 
        .Q(\inq_ary[10][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N977), 
        .Q(\inq_ary[10][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N977), 
        .Q(\inq_ary[10][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N977), 
        .Q(\inq_ary[10][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N977), 
        .Q(\inq_ary[10][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N977), 
        .Q(\inq_ary[10][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N977), 
        .Q(\inq_ary[10][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N977), 
        .Q(\inq_ary[10][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N977), 
        .Q(\inq_ary[10][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N977), 
        .Q(\inq_ary[10][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N977), 
        .Q(\inq_ary[10][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N977), 
        .Q(\inq_ary[10][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N977), 
        .Q(\inq_ary[10][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N977), 
        .Q(\inq_ary[10][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N977), 
        .Q(\inq_ary[10][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N977), 
        .Q(\inq_ary[10][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N977), 
        .Q(\inq_ary[10][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N977), 
        .Q(\inq_ary[10][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N977), 
        .Q(\inq_ary[10][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N977), 
        .Q(\inq_ary[10][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N977), 
        .Q(\inq_ary[10][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N977), 
        .Q(\inq_ary[10][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N977), 
        .Q(\inq_ary[10][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N977), 
        .Q(\inq_ary[10][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N977), 
        .Q(\inq_ary[10][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N977), 
        .Q(\inq_ary[10][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N977), 
        .Q(\inq_ary[10][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N977), 
        .Q(\inq_ary[10][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N977), 
        .Q(\inq_ary[10][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N977), 
        .Q(\inq_ary[10][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N977), 
        .Q(\inq_ary[10][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N977), 
        .Q(\inq_ary[10][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N977), 
        .Q(\inq_ary[10][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N977), 
        .Q(\inq_ary[10][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N977), 
        .Q(\inq_ary[10][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N977), 
        .Q(\inq_ary[10][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N977), 
        .Q(\inq_ary[10][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N977), 
        .Q(\inq_ary[10][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N977), 
        .Q(\inq_ary[10][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N977), 
        .Q(\inq_ary[10][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N977), 
        .Q(\inq_ary[10][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N977), 
        .Q(\inq_ary[10][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N977), 
        .Q(\inq_ary[10][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N977), 
        .Q(\inq_ary[10][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N977), 
        .Q(\inq_ary[10][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N977), 
        .Q(\inq_ary[10][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N977), 
        .Q(\inq_ary[10][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N977), 
        .Q(\inq_ary[10][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N977), 
        .Q(\inq_ary[10][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N977), 
        .Q(\inq_ary[10][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N977), 
        .Q(\inq_ary[10][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N977), 
        .Q(\inq_ary[10][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N977), 
        .Q(\inq_ary[10][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N977), 
        .Q(\inq_ary[10][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N977), 
        .Q(\inq_ary[10][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N977), 
        .Q(\inq_ary[10][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N977), 
        .Q(\inq_ary[10][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N977), 
        .Q(\inq_ary[10][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N977), 
        .Q(\inq_ary[10][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N977), 
        .Q(\inq_ary[10][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N977), 
        .Q(\inq_ary[10][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N977), 
        .Q(\inq_ary[10][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N977), 
        .Q(\inq_ary[10][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N977), 
        .Q(\inq_ary[10][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N977), 
        .Q(\inq_ary[10][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N977), 
        .Q(\inq_ary[10][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N977), 
        .Q(\inq_ary[10][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N977), 
        .Q(\inq_ary[10][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N977), 
        .Q(\inq_ary[10][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N977), 
        .Q(\inq_ary[10][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N977), 
        .Q(\inq_ary[10][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N977), 
        .Q(\inq_ary[10][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N977), 
        .Q(\inq_ary[10][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N977), 
        .Q(\inq_ary[10][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N977), 
        .Q(\inq_ary[10][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N977), 
        .Q(\inq_ary[10][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N977), 
        .Q(\inq_ary[10][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N977), 
        .Q(\inq_ary[10][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N977), 
        .Q(\inq_ary[10][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N977), 
        .Q(\inq_ary[10][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N977), 
        .Q(\inq_ary[10][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N977), 
        .Q(\inq_ary[10][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N977), 
        .Q(\inq_ary[10][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N977), 
        .Q(\inq_ary[10][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][9]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N977), 
        .Q(\inq_ary[10][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][8]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N977), 
        .Q(\inq_ary[10][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][7]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N977), 
        .Q(\inq_ary[10][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][6]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N977), 
        .Q(\inq_ary[10][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][5]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N977), 
        .Q(\inq_ary[10][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][4]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N977), 
        .Q(\inq_ary[10][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][3]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N977), 
        .Q(\inq_ary[10][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][2]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N977), 
        .Q(\inq_ary[10][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][1]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N977), 
        .Q(\inq_ary[10][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[10][0]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N977), 
        .Q(\inq_ary[10][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N976), 
        .Q(\inq_ary[9][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N976), 
        .Q(\inq_ary[9][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N976), 
        .Q(\inq_ary[9][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N976), 
        .Q(\inq_ary[9][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N976), 
        .Q(\inq_ary[9][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N976), 
        .Q(\inq_ary[9][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N976), 
        .Q(\inq_ary[9][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N976), 
        .Q(\inq_ary[9][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N976), 
        .Q(\inq_ary[9][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N976), 
        .Q(\inq_ary[9][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N976), 
        .Q(\inq_ary[9][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N976), 
        .Q(\inq_ary[9][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N976), 
        .Q(\inq_ary[9][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N976), 
        .Q(\inq_ary[9][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N976), 
        .Q(\inq_ary[9][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N976), 
        .Q(\inq_ary[9][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N976), 
        .Q(\inq_ary[9][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N976), 
        .Q(\inq_ary[9][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N976), 
        .Q(\inq_ary[9][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N976), 
        .Q(\inq_ary[9][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N976), 
        .Q(\inq_ary[9][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N976), 
        .Q(\inq_ary[9][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N976), 
        .Q(\inq_ary[9][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N976), 
        .Q(\inq_ary[9][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N976), 
        .Q(\inq_ary[9][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N976), 
        .Q(\inq_ary[9][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N976), 
        .Q(\inq_ary[9][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N976), 
        .Q(\inq_ary[9][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N976), 
        .Q(\inq_ary[9][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N976), 
        .Q(\inq_ary[9][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N976), 
        .Q(\inq_ary[9][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N976), 
        .Q(\inq_ary[9][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N976), 
        .Q(\inq_ary[9][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N976), 
        .Q(\inq_ary[9][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N976), 
        .Q(\inq_ary[9][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N976), 
        .Q(\inq_ary[9][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N976), 
        .Q(\inq_ary[9][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N976), 
        .Q(\inq_ary[9][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N976), 
        .Q(\inq_ary[9][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N976), 
        .Q(\inq_ary[9][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N976), 
        .Q(\inq_ary[9][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N976), 
        .Q(\inq_ary[9][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N976), 
        .Q(\inq_ary[9][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N976), 
        .Q(\inq_ary[9][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N976), 
        .Q(\inq_ary[9][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N976), 
        .Q(\inq_ary[9][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N976), 
        .Q(\inq_ary[9][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N976), 
        .Q(\inq_ary[9][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N976), 
        .Q(\inq_ary[9][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N976), 
        .Q(\inq_ary[9][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N976), 
        .Q(\inq_ary[9][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N976), 
        .Q(\inq_ary[9][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N976), 
        .Q(\inq_ary[9][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N976), 
        .Q(\inq_ary[9][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N976), 
        .Q(\inq_ary[9][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N976), 
        .Q(\inq_ary[9][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N976), 
        .Q(\inq_ary[9][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N976), 
        .Q(\inq_ary[9][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N976), 
        .Q(\inq_ary[9][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N976), 
        .Q(\inq_ary[9][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N976), 
        .Q(\inq_ary[9][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N975), 
        .Q(\inq_ary[9][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N975), 
        .Q(\inq_ary[9][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N975), 
        .Q(\inq_ary[9][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N975), 
        .Q(\inq_ary[9][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N975), 
        .Q(\inq_ary[9][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N975), 
        .Q(\inq_ary[9][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N975), 
        .Q(\inq_ary[9][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N975), 
        .Q(\inq_ary[9][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N975), 
        .Q(\inq_ary[9][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N975), 
        .Q(\inq_ary[9][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N975), 
        .Q(\inq_ary[9][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N975), 
        .Q(\inq_ary[9][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N975), 
        .Q(\inq_ary[9][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N975), 
        .Q(\inq_ary[9][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N975), 
        .Q(\inq_ary[9][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N975), 
        .Q(\inq_ary[9][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N975), 
        .Q(\inq_ary[9][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N975), 
        .Q(\inq_ary[9][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N975), 
        .Q(\inq_ary[9][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N975), 
        .Q(\inq_ary[9][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N975), 
        .Q(\inq_ary[9][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N975), 
        .Q(\inq_ary[9][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N975), 
        .Q(\inq_ary[9][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N975), 
        .Q(\inq_ary[9][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N975), 
        .Q(\inq_ary[9][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N975), 
        .Q(\inq_ary[9][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N975), 
        .Q(\inq_ary[9][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N975), 
        .Q(\inq_ary[9][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N975), 
        .Q(\inq_ary[9][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N975), 
        .Q(\inq_ary[9][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N975), 
        .Q(\inq_ary[9][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N975), 
        .Q(\inq_ary[9][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N975), 
        .Q(\inq_ary[9][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N975), 
        .Q(\inq_ary[9][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N975), 
        .Q(\inq_ary[9][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N975), 
        .Q(\inq_ary[9][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N975), 
        .Q(\inq_ary[9][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N975), 
        .Q(\inq_ary[9][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N975), 
        .Q(\inq_ary[9][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N975), 
        .Q(\inq_ary[9][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N975), 
        .Q(\inq_ary[9][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N975), 
        .Q(\inq_ary[9][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N975), 
        .Q(\inq_ary[9][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N975), 
        .Q(\inq_ary[9][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N975), 
        .Q(\inq_ary[9][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N975), 
        .Q(\inq_ary[9][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N975), 
        .Q(\inq_ary[9][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N975), 
        .Q(\inq_ary[9][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N975), 
        .Q(\inq_ary[9][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N975), 
        .Q(\inq_ary[9][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N975), 
        .Q(\inq_ary[9][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N975), 
        .Q(\inq_ary[9][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N975), 
        .Q(\inq_ary[9][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N975), 
        .Q(\inq_ary[9][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N975), 
        .Q(\inq_ary[9][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N975), 
        .Q(\inq_ary[9][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N975), 
        .Q(\inq_ary[9][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N975), 
        .Q(\inq_ary[9][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N975), 
        .Q(\inq_ary[9][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N975), 
        .Q(\inq_ary[9][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N975), 
        .Q(\inq_ary[9][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N975), 
        .Q(\inq_ary[9][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N975), 
        .Q(\inq_ary[9][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N975), 
        .Q(\inq_ary[9][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N975), 
        .Q(\inq_ary[9][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N975), 
        .Q(\inq_ary[9][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N975), 
        .Q(\inq_ary[9][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N975), 
        .Q(\inq_ary[9][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N975), 
        .Q(\inq_ary[9][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N975), 
        .Q(\inq_ary[9][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N975), 
        .Q(\inq_ary[9][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N975), 
        .Q(\inq_ary[9][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N975), 
        .Q(\inq_ary[9][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N975), 
        .Q(\inq_ary[9][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N975), 
        .Q(\inq_ary[9][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N975), 
        .Q(\inq_ary[9][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N975), 
        .Q(\inq_ary[9][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N975), 
        .Q(\inq_ary[9][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N975), 
        .Q(\inq_ary[9][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N975), 
        .Q(\inq_ary[9][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N975), 
        .Q(\inq_ary[9][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N975), 
        .Q(\inq_ary[9][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N975), 
        .Q(\inq_ary[9][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N975), 
        .Q(\inq_ary[9][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N975), 
        .Q(\inq_ary[9][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N975), 
        .Q(\inq_ary[9][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N975), 
        .Q(\inq_ary[9][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N975), 
        .Q(\inq_ary[9][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N975), 
        .Q(\inq_ary[9][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N975), .Q(
        \inq_ary[9][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N975), .Q(
        \inq_ary[9][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N975), .Q(
        \inq_ary[9][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N975), .Q(
        \inq_ary[9][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N975), .Q(
        \inq_ary[9][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N975), .Q(
        \inq_ary[9][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N975), .Q(
        \inq_ary[9][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N975), .Q(
        \inq_ary[9][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N975), .Q(
        \inq_ary[9][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[9][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N975), .Q(
        \inq_ary[9][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N974), 
        .Q(\inq_ary[8][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N974), 
        .Q(\inq_ary[8][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N974), 
        .Q(\inq_ary[8][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N974), 
        .Q(\inq_ary[8][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N974), 
        .Q(\inq_ary[8][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N974), 
        .Q(\inq_ary[8][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N974), 
        .Q(\inq_ary[8][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N974), 
        .Q(\inq_ary[8][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N974), 
        .Q(\inq_ary[8][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N974), 
        .Q(\inq_ary[8][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N974), 
        .Q(\inq_ary[8][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N974), 
        .Q(\inq_ary[8][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N974), 
        .Q(\inq_ary[8][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N974), 
        .Q(\inq_ary[8][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N974), 
        .Q(\inq_ary[8][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N974), 
        .Q(\inq_ary[8][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N974), 
        .Q(\inq_ary[8][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N974), 
        .Q(\inq_ary[8][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N974), 
        .Q(\inq_ary[8][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N974), 
        .Q(\inq_ary[8][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N974), 
        .Q(\inq_ary[8][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N974), 
        .Q(\inq_ary[8][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N974), 
        .Q(\inq_ary[8][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N974), 
        .Q(\inq_ary[8][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N974), 
        .Q(\inq_ary[8][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N974), 
        .Q(\inq_ary[8][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N974), 
        .Q(\inq_ary[8][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N974), 
        .Q(\inq_ary[8][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N974), 
        .Q(\inq_ary[8][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N974), 
        .Q(\inq_ary[8][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N974), 
        .Q(\inq_ary[8][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N974), 
        .Q(\inq_ary[8][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N974), 
        .Q(\inq_ary[8][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N974), 
        .Q(\inq_ary[8][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N974), 
        .Q(\inq_ary[8][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N974), 
        .Q(\inq_ary[8][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N974), 
        .Q(\inq_ary[8][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N974), 
        .Q(\inq_ary[8][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N974), 
        .Q(\inq_ary[8][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N974), 
        .Q(\inq_ary[8][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N974), 
        .Q(\inq_ary[8][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N974), 
        .Q(\inq_ary[8][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N974), 
        .Q(\inq_ary[8][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N974), 
        .Q(\inq_ary[8][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N974), 
        .Q(\inq_ary[8][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N974), 
        .Q(\inq_ary[8][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N974), 
        .Q(\inq_ary[8][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N974), 
        .Q(\inq_ary[8][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N974), 
        .Q(\inq_ary[8][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N974), 
        .Q(\inq_ary[8][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N974), 
        .Q(\inq_ary[8][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N974), 
        .Q(\inq_ary[8][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N974), 
        .Q(\inq_ary[8][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N974), 
        .Q(\inq_ary[8][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N974), 
        .Q(\inq_ary[8][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N974), 
        .Q(\inq_ary[8][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N974), 
        .Q(\inq_ary[8][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N974), 
        .Q(\inq_ary[8][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N974), 
        .Q(\inq_ary[8][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N974), 
        .Q(\inq_ary[8][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N974), 
        .Q(\inq_ary[8][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N973), 
        .Q(\inq_ary[8][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N973), 
        .Q(\inq_ary[8][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N973), 
        .Q(\inq_ary[8][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N973), 
        .Q(\inq_ary[8][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N973), 
        .Q(\inq_ary[8][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N973), 
        .Q(\inq_ary[8][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N973), 
        .Q(\inq_ary[8][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N973), 
        .Q(\inq_ary[8][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N973), 
        .Q(\inq_ary[8][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N973), 
        .Q(\inq_ary[8][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N973), 
        .Q(\inq_ary[8][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N973), 
        .Q(\inq_ary[8][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N973), 
        .Q(\inq_ary[8][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N973), 
        .Q(\inq_ary[8][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N973), 
        .Q(\inq_ary[8][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N973), 
        .Q(\inq_ary[8][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N973), 
        .Q(\inq_ary[8][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N973), 
        .Q(\inq_ary[8][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N973), 
        .Q(\inq_ary[8][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N973), 
        .Q(\inq_ary[8][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N973), 
        .Q(\inq_ary[8][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N973), 
        .Q(\inq_ary[8][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N973), 
        .Q(\inq_ary[8][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N973), 
        .Q(\inq_ary[8][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N973), 
        .Q(\inq_ary[8][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N973), 
        .Q(\inq_ary[8][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N973), 
        .Q(\inq_ary[8][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N973), 
        .Q(\inq_ary[8][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N973), 
        .Q(\inq_ary[8][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N973), 
        .Q(\inq_ary[8][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N973), 
        .Q(\inq_ary[8][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N973), 
        .Q(\inq_ary[8][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N973), 
        .Q(\inq_ary[8][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N973), 
        .Q(\inq_ary[8][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N973), 
        .Q(\inq_ary[8][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N973), 
        .Q(\inq_ary[8][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N973), 
        .Q(\inq_ary[8][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N973), 
        .Q(\inq_ary[8][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N973), 
        .Q(\inq_ary[8][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N973), 
        .Q(\inq_ary[8][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N973), 
        .Q(\inq_ary[8][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N973), 
        .Q(\inq_ary[8][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N973), 
        .Q(\inq_ary[8][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N973), 
        .Q(\inq_ary[8][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N973), 
        .Q(\inq_ary[8][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N973), 
        .Q(\inq_ary[8][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N973), 
        .Q(\inq_ary[8][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N973), 
        .Q(\inq_ary[8][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N973), 
        .Q(\inq_ary[8][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N973), 
        .Q(\inq_ary[8][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N973), 
        .Q(\inq_ary[8][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N973), 
        .Q(\inq_ary[8][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N973), 
        .Q(\inq_ary[8][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N973), 
        .Q(\inq_ary[8][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N973), 
        .Q(\inq_ary[8][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N973), 
        .Q(\inq_ary[8][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N973), 
        .Q(\inq_ary[8][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N973), 
        .Q(\inq_ary[8][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N973), 
        .Q(\inq_ary[8][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N973), 
        .Q(\inq_ary[8][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N973), 
        .Q(\inq_ary[8][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N973), 
        .Q(\inq_ary[8][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N973), 
        .Q(\inq_ary[8][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N973), 
        .Q(\inq_ary[8][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N973), 
        .Q(\inq_ary[8][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N973), 
        .Q(\inq_ary[8][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N973), 
        .Q(\inq_ary[8][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N973), 
        .Q(\inq_ary[8][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N973), 
        .Q(\inq_ary[8][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N973), 
        .Q(\inq_ary[8][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N973), 
        .Q(\inq_ary[8][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N973), 
        .Q(\inq_ary[8][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N973), 
        .Q(\inq_ary[8][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N973), 
        .Q(\inq_ary[8][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N973), 
        .Q(\inq_ary[8][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N973), 
        .Q(\inq_ary[8][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N973), 
        .Q(\inq_ary[8][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N973), 
        .Q(\inq_ary[8][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N973), 
        .Q(\inq_ary[8][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N973), 
        .Q(\inq_ary[8][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N973), 
        .Q(\inq_ary[8][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N973), 
        .Q(\inq_ary[8][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N973), 
        .Q(\inq_ary[8][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N973), 
        .Q(\inq_ary[8][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N973), 
        .Q(\inq_ary[8][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N973), 
        .Q(\inq_ary[8][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N973), 
        .Q(\inq_ary[8][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N973), 
        .Q(\inq_ary[8][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N973), 
        .Q(\inq_ary[8][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N973), .Q(
        \inq_ary[8][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N973), .Q(
        \inq_ary[8][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N973), .Q(
        \inq_ary[8][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N973), .Q(
        \inq_ary[8][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N973), .Q(
        \inq_ary[8][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N973), .Q(
        \inq_ary[8][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N973), .Q(
        \inq_ary[8][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N973), .Q(
        \inq_ary[8][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N973), .Q(
        \inq_ary[8][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[8][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N973), .Q(
        \inq_ary[8][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N972), 
        .Q(\inq_ary[7][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N972), 
        .Q(\inq_ary[7][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N972), 
        .Q(\inq_ary[7][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N972), 
        .Q(\inq_ary[7][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N972), 
        .Q(\inq_ary[7][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N972), 
        .Q(\inq_ary[7][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N972), 
        .Q(\inq_ary[7][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N972), 
        .Q(\inq_ary[7][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N972), 
        .Q(\inq_ary[7][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N972), 
        .Q(\inq_ary[7][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N972), 
        .Q(\inq_ary[7][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N972), 
        .Q(\inq_ary[7][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N972), 
        .Q(\inq_ary[7][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N972), 
        .Q(\inq_ary[7][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N972), 
        .Q(\inq_ary[7][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N972), 
        .Q(\inq_ary[7][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N972), 
        .Q(\inq_ary[7][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N972), 
        .Q(\inq_ary[7][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N972), 
        .Q(\inq_ary[7][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N972), 
        .Q(\inq_ary[7][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N972), 
        .Q(\inq_ary[7][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N972), 
        .Q(\inq_ary[7][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N972), 
        .Q(\inq_ary[7][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N972), 
        .Q(\inq_ary[7][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N972), 
        .Q(\inq_ary[7][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N972), 
        .Q(\inq_ary[7][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N972), 
        .Q(\inq_ary[7][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N972), 
        .Q(\inq_ary[7][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N972), 
        .Q(\inq_ary[7][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N972), 
        .Q(\inq_ary[7][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N972), 
        .Q(\inq_ary[7][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N972), 
        .Q(\inq_ary[7][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N972), 
        .Q(\inq_ary[7][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N972), 
        .Q(\inq_ary[7][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N972), 
        .Q(\inq_ary[7][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N972), 
        .Q(\inq_ary[7][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N972), 
        .Q(\inq_ary[7][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N972), 
        .Q(\inq_ary[7][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N972), 
        .Q(\inq_ary[7][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N972), 
        .Q(\inq_ary[7][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N972), 
        .Q(\inq_ary[7][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N972), 
        .Q(\inq_ary[7][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N972), 
        .Q(\inq_ary[7][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N972), 
        .Q(\inq_ary[7][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N972), 
        .Q(\inq_ary[7][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N972), 
        .Q(\inq_ary[7][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N972), 
        .Q(\inq_ary[7][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N972), 
        .Q(\inq_ary[7][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N972), 
        .Q(\inq_ary[7][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N972), 
        .Q(\inq_ary[7][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N972), 
        .Q(\inq_ary[7][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N972), 
        .Q(\inq_ary[7][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N972), 
        .Q(\inq_ary[7][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N972), 
        .Q(\inq_ary[7][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N972), 
        .Q(\inq_ary[7][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N972), 
        .Q(\inq_ary[7][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N972), 
        .Q(\inq_ary[7][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N972), 
        .Q(\inq_ary[7][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N972), 
        .Q(\inq_ary[7][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N972), 
        .Q(\inq_ary[7][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N972), 
        .Q(\inq_ary[7][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N971), 
        .Q(\inq_ary[7][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N971), 
        .Q(\inq_ary[7][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N971), 
        .Q(\inq_ary[7][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N971), 
        .Q(\inq_ary[7][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N971), 
        .Q(\inq_ary[7][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N971), 
        .Q(\inq_ary[7][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N971), 
        .Q(\inq_ary[7][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N971), 
        .Q(\inq_ary[7][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N971), 
        .Q(\inq_ary[7][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N971), 
        .Q(\inq_ary[7][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N971), 
        .Q(\inq_ary[7][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N971), 
        .Q(\inq_ary[7][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N971), 
        .Q(\inq_ary[7][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N971), 
        .Q(\inq_ary[7][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N971), 
        .Q(\inq_ary[7][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N971), 
        .Q(\inq_ary[7][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N971), 
        .Q(\inq_ary[7][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N971), 
        .Q(\inq_ary[7][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N971), 
        .Q(\inq_ary[7][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N971), 
        .Q(\inq_ary[7][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N971), 
        .Q(\inq_ary[7][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N971), 
        .Q(\inq_ary[7][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N971), 
        .Q(\inq_ary[7][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N971), 
        .Q(\inq_ary[7][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N971), 
        .Q(\inq_ary[7][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N971), 
        .Q(\inq_ary[7][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N971), 
        .Q(\inq_ary[7][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N971), 
        .Q(\inq_ary[7][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N971), 
        .Q(\inq_ary[7][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N971), 
        .Q(\inq_ary[7][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N971), 
        .Q(\inq_ary[7][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N971), 
        .Q(\inq_ary[7][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N971), 
        .Q(\inq_ary[7][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N971), 
        .Q(\inq_ary[7][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N971), 
        .Q(\inq_ary[7][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N971), 
        .Q(\inq_ary[7][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N971), 
        .Q(\inq_ary[7][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N971), 
        .Q(\inq_ary[7][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N971), 
        .Q(\inq_ary[7][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N971), 
        .Q(\inq_ary[7][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N971), 
        .Q(\inq_ary[7][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N971), 
        .Q(\inq_ary[7][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N971), 
        .Q(\inq_ary[7][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N971), 
        .Q(\inq_ary[7][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N971), 
        .Q(\inq_ary[7][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N971), 
        .Q(\inq_ary[7][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N971), 
        .Q(\inq_ary[7][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N971), 
        .Q(\inq_ary[7][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N971), 
        .Q(\inq_ary[7][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N971), 
        .Q(\inq_ary[7][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N971), 
        .Q(\inq_ary[7][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N971), 
        .Q(\inq_ary[7][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N971), 
        .Q(\inq_ary[7][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N971), 
        .Q(\inq_ary[7][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N971), 
        .Q(\inq_ary[7][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N971), 
        .Q(\inq_ary[7][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N971), 
        .Q(\inq_ary[7][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N971), 
        .Q(\inq_ary[7][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N971), 
        .Q(\inq_ary[7][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N971), 
        .Q(\inq_ary[7][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N971), 
        .Q(\inq_ary[7][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N971), 
        .Q(\inq_ary[7][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N971), 
        .Q(\inq_ary[7][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N971), 
        .Q(\inq_ary[7][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N971), 
        .Q(\inq_ary[7][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N971), 
        .Q(\inq_ary[7][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N971), 
        .Q(\inq_ary[7][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N971), 
        .Q(\inq_ary[7][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N971), 
        .Q(\inq_ary[7][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N971), 
        .Q(\inq_ary[7][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N971), 
        .Q(\inq_ary[7][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N971), 
        .Q(\inq_ary[7][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N971), 
        .Q(\inq_ary[7][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N971), 
        .Q(\inq_ary[7][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N971), 
        .Q(\inq_ary[7][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N971), 
        .Q(\inq_ary[7][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N971), 
        .Q(\inq_ary[7][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N971), 
        .Q(\inq_ary[7][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N971), 
        .Q(\inq_ary[7][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N971), 
        .Q(\inq_ary[7][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N971), 
        .Q(\inq_ary[7][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N971), 
        .Q(\inq_ary[7][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N971), 
        .Q(\inq_ary[7][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N971), 
        .Q(\inq_ary[7][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N971), 
        .Q(\inq_ary[7][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N971), 
        .Q(\inq_ary[7][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N971), 
        .Q(\inq_ary[7][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N971), 
        .Q(\inq_ary[7][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N971), 
        .Q(\inq_ary[7][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N971), .Q(
        \inq_ary[7][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N971), .Q(
        \inq_ary[7][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N971), .Q(
        \inq_ary[7][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N971), .Q(
        \inq_ary[7][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N971), .Q(
        \inq_ary[7][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N971), .Q(
        \inq_ary[7][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N971), .Q(
        \inq_ary[7][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N971), .Q(
        \inq_ary[7][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N971), .Q(
        \inq_ary[7][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[7][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N971), .Q(
        \inq_ary[7][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N970), 
        .Q(\inq_ary[6][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N970), 
        .Q(\inq_ary[6][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N970), 
        .Q(\inq_ary[6][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N970), 
        .Q(\inq_ary[6][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N970), 
        .Q(\inq_ary[6][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N970), 
        .Q(\inq_ary[6][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N970), 
        .Q(\inq_ary[6][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N970), 
        .Q(\inq_ary[6][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N970), 
        .Q(\inq_ary[6][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N970), 
        .Q(\inq_ary[6][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N970), 
        .Q(\inq_ary[6][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N970), 
        .Q(\inq_ary[6][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N970), 
        .Q(\inq_ary[6][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N970), 
        .Q(\inq_ary[6][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N970), 
        .Q(\inq_ary[6][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N970), 
        .Q(\inq_ary[6][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N970), 
        .Q(\inq_ary[6][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N970), 
        .Q(\inq_ary[6][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N970), 
        .Q(\inq_ary[6][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N970), 
        .Q(\inq_ary[6][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N970), 
        .Q(\inq_ary[6][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N970), 
        .Q(\inq_ary[6][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N970), 
        .Q(\inq_ary[6][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N970), 
        .Q(\inq_ary[6][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N970), 
        .Q(\inq_ary[6][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N970), 
        .Q(\inq_ary[6][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N970), 
        .Q(\inq_ary[6][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N970), 
        .Q(\inq_ary[6][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N970), 
        .Q(\inq_ary[6][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N970), 
        .Q(\inq_ary[6][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N970), 
        .Q(\inq_ary[6][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N970), 
        .Q(\inq_ary[6][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N970), 
        .Q(\inq_ary[6][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N970), 
        .Q(\inq_ary[6][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N970), 
        .Q(\inq_ary[6][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N970), 
        .Q(\inq_ary[6][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N970), 
        .Q(\inq_ary[6][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N970), 
        .Q(\inq_ary[6][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N970), 
        .Q(\inq_ary[6][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N970), 
        .Q(\inq_ary[6][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N970), 
        .Q(\inq_ary[6][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N970), 
        .Q(\inq_ary[6][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N970), 
        .Q(\inq_ary[6][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N970), 
        .Q(\inq_ary[6][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N970), 
        .Q(\inq_ary[6][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N970), 
        .Q(\inq_ary[6][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N970), 
        .Q(\inq_ary[6][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N970), 
        .Q(\inq_ary[6][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N970), 
        .Q(\inq_ary[6][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N970), 
        .Q(\inq_ary[6][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N970), 
        .Q(\inq_ary[6][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N970), 
        .Q(\inq_ary[6][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N970), 
        .Q(\inq_ary[6][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N970), 
        .Q(\inq_ary[6][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N970), 
        .Q(\inq_ary[6][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N970), 
        .Q(\inq_ary[6][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N970), 
        .Q(\inq_ary[6][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N970), 
        .Q(\inq_ary[6][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N970), 
        .Q(\inq_ary[6][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N970), 
        .Q(\inq_ary[6][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N970), 
        .Q(\inq_ary[6][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N969), 
        .Q(\inq_ary[6][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N969), 
        .Q(\inq_ary[6][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N969), 
        .Q(\inq_ary[6][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N969), 
        .Q(\inq_ary[6][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N969), 
        .Q(\inq_ary[6][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N969), 
        .Q(\inq_ary[6][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N969), 
        .Q(\inq_ary[6][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N969), 
        .Q(\inq_ary[6][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N969), 
        .Q(\inq_ary[6][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N969), 
        .Q(\inq_ary[6][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N969), 
        .Q(\inq_ary[6][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N969), 
        .Q(\inq_ary[6][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N969), 
        .Q(\inq_ary[6][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N969), 
        .Q(\inq_ary[6][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N969), 
        .Q(\inq_ary[6][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N969), 
        .Q(\inq_ary[6][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N969), 
        .Q(\inq_ary[6][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N969), 
        .Q(\inq_ary[6][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N969), 
        .Q(\inq_ary[6][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N969), 
        .Q(\inq_ary[6][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N969), 
        .Q(\inq_ary[6][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N969), 
        .Q(\inq_ary[6][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N969), 
        .Q(\inq_ary[6][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N969), 
        .Q(\inq_ary[6][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N969), 
        .Q(\inq_ary[6][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N969), 
        .Q(\inq_ary[6][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N969), 
        .Q(\inq_ary[6][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N969), 
        .Q(\inq_ary[6][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N969), 
        .Q(\inq_ary[6][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N969), 
        .Q(\inq_ary[6][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N969), 
        .Q(\inq_ary[6][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N969), 
        .Q(\inq_ary[6][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N969), 
        .Q(\inq_ary[6][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N969), 
        .Q(\inq_ary[6][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N969), 
        .Q(\inq_ary[6][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N969), 
        .Q(\inq_ary[6][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N969), 
        .Q(\inq_ary[6][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N969), 
        .Q(\inq_ary[6][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N969), 
        .Q(\inq_ary[6][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N969), 
        .Q(\inq_ary[6][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N969), 
        .Q(\inq_ary[6][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N969), 
        .Q(\inq_ary[6][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N969), 
        .Q(\inq_ary[6][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N969), 
        .Q(\inq_ary[6][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N969), 
        .Q(\inq_ary[6][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N969), 
        .Q(\inq_ary[6][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N969), 
        .Q(\inq_ary[6][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N969), 
        .Q(\inq_ary[6][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N969), 
        .Q(\inq_ary[6][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N969), 
        .Q(\inq_ary[6][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N969), 
        .Q(\inq_ary[6][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N969), 
        .Q(\inq_ary[6][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N969), 
        .Q(\inq_ary[6][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N969), 
        .Q(\inq_ary[6][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N969), 
        .Q(\inq_ary[6][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N969), 
        .Q(\inq_ary[6][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N969), 
        .Q(\inq_ary[6][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N969), 
        .Q(\inq_ary[6][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N969), 
        .Q(\inq_ary[6][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N969), 
        .Q(\inq_ary[6][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N969), 
        .Q(\inq_ary[6][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N969), 
        .Q(\inq_ary[6][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N969), 
        .Q(\inq_ary[6][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N969), 
        .Q(\inq_ary[6][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N969), 
        .Q(\inq_ary[6][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N969), 
        .Q(\inq_ary[6][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N969), 
        .Q(\inq_ary[6][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N969), 
        .Q(\inq_ary[6][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N969), 
        .Q(\inq_ary[6][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N969), 
        .Q(\inq_ary[6][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N969), 
        .Q(\inq_ary[6][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N969), 
        .Q(\inq_ary[6][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N969), 
        .Q(\inq_ary[6][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N969), 
        .Q(\inq_ary[6][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N969), 
        .Q(\inq_ary[6][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N969), 
        .Q(\inq_ary[6][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N969), 
        .Q(\inq_ary[6][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N969), 
        .Q(\inq_ary[6][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N969), 
        .Q(\inq_ary[6][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N969), 
        .Q(\inq_ary[6][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N969), 
        .Q(\inq_ary[6][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N969), 
        .Q(\inq_ary[6][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N969), 
        .Q(\inq_ary[6][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N969), 
        .Q(\inq_ary[6][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N969), 
        .Q(\inq_ary[6][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N969), 
        .Q(\inq_ary[6][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N969), 
        .Q(\inq_ary[6][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N969), 
        .Q(\inq_ary[6][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N969), 
        .Q(\inq_ary[6][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N969), .Q(
        \inq_ary[6][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N969), .Q(
        \inq_ary[6][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N969), .Q(
        \inq_ary[6][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N969), .Q(
        \inq_ary[6][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N969), .Q(
        \inq_ary[6][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N969), .Q(
        \inq_ary[6][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N969), .Q(
        \inq_ary[6][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N969), .Q(
        \inq_ary[6][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N969), .Q(
        \inq_ary[6][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[6][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N969), .Q(
        \inq_ary[6][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N968), 
        .Q(\inq_ary[5][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N968), 
        .Q(\inq_ary[5][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N968), 
        .Q(\inq_ary[5][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N968), 
        .Q(\inq_ary[5][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N968), 
        .Q(\inq_ary[5][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N968), 
        .Q(\inq_ary[5][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N968), 
        .Q(\inq_ary[5][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N968), 
        .Q(\inq_ary[5][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N968), 
        .Q(\inq_ary[5][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N968), 
        .Q(\inq_ary[5][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N968), 
        .Q(\inq_ary[5][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N968), 
        .Q(\inq_ary[5][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N968), 
        .Q(\inq_ary[5][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N968), 
        .Q(\inq_ary[5][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N968), 
        .Q(\inq_ary[5][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N968), 
        .Q(\inq_ary[5][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N968), 
        .Q(\inq_ary[5][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N968), 
        .Q(\inq_ary[5][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N968), 
        .Q(\inq_ary[5][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N968), 
        .Q(\inq_ary[5][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N968), 
        .Q(\inq_ary[5][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N968), 
        .Q(\inq_ary[5][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N968), 
        .Q(\inq_ary[5][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N968), 
        .Q(\inq_ary[5][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N968), 
        .Q(\inq_ary[5][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N968), 
        .Q(\inq_ary[5][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N968), 
        .Q(\inq_ary[5][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N968), 
        .Q(\inq_ary[5][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N968), 
        .Q(\inq_ary[5][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N968), 
        .Q(\inq_ary[5][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N968), 
        .Q(\inq_ary[5][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N968), 
        .Q(\inq_ary[5][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N968), 
        .Q(\inq_ary[5][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N968), 
        .Q(\inq_ary[5][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N968), 
        .Q(\inq_ary[5][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N968), 
        .Q(\inq_ary[5][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N968), 
        .Q(\inq_ary[5][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N968), 
        .Q(\inq_ary[5][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N968), 
        .Q(\inq_ary[5][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N968), 
        .Q(\inq_ary[5][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N968), 
        .Q(\inq_ary[5][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N968), 
        .Q(\inq_ary[5][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N968), 
        .Q(\inq_ary[5][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N968), 
        .Q(\inq_ary[5][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N968), 
        .Q(\inq_ary[5][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N968), 
        .Q(\inq_ary[5][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N968), 
        .Q(\inq_ary[5][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N968), 
        .Q(\inq_ary[5][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N968), 
        .Q(\inq_ary[5][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N968), 
        .Q(\inq_ary[5][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N968), 
        .Q(\inq_ary[5][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N968), 
        .Q(\inq_ary[5][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N968), 
        .Q(\inq_ary[5][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N968), 
        .Q(\inq_ary[5][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N968), 
        .Q(\inq_ary[5][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N968), 
        .Q(\inq_ary[5][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N968), 
        .Q(\inq_ary[5][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N968), 
        .Q(\inq_ary[5][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N968), 
        .Q(\inq_ary[5][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N968), 
        .Q(\inq_ary[5][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N968), 
        .Q(\inq_ary[5][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N967), 
        .Q(\inq_ary[5][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N967), 
        .Q(\inq_ary[5][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N967), 
        .Q(\inq_ary[5][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N967), 
        .Q(\inq_ary[5][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N967), 
        .Q(\inq_ary[5][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N967), 
        .Q(\inq_ary[5][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N967), 
        .Q(\inq_ary[5][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N967), 
        .Q(\inq_ary[5][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N967), 
        .Q(\inq_ary[5][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N967), 
        .Q(\inq_ary[5][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N967), 
        .Q(\inq_ary[5][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N967), 
        .Q(\inq_ary[5][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N967), 
        .Q(\inq_ary[5][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N967), 
        .Q(\inq_ary[5][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N967), 
        .Q(\inq_ary[5][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N967), 
        .Q(\inq_ary[5][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N967), 
        .Q(\inq_ary[5][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N967), 
        .Q(\inq_ary[5][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N967), 
        .Q(\inq_ary[5][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N967), 
        .Q(\inq_ary[5][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N967), 
        .Q(\inq_ary[5][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N967), 
        .Q(\inq_ary[5][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N967), 
        .Q(\inq_ary[5][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N967), 
        .Q(\inq_ary[5][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N967), 
        .Q(\inq_ary[5][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N967), 
        .Q(\inq_ary[5][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N967), 
        .Q(\inq_ary[5][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N967), 
        .Q(\inq_ary[5][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N967), 
        .Q(\inq_ary[5][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N967), 
        .Q(\inq_ary[5][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N967), 
        .Q(\inq_ary[5][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N967), 
        .Q(\inq_ary[5][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N967), 
        .Q(\inq_ary[5][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N967), 
        .Q(\inq_ary[5][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N967), 
        .Q(\inq_ary[5][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N967), 
        .Q(\inq_ary[5][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N967), 
        .Q(\inq_ary[5][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N967), 
        .Q(\inq_ary[5][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N967), 
        .Q(\inq_ary[5][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N967), 
        .Q(\inq_ary[5][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N967), 
        .Q(\inq_ary[5][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N967), 
        .Q(\inq_ary[5][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N967), 
        .Q(\inq_ary[5][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N967), 
        .Q(\inq_ary[5][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N967), 
        .Q(\inq_ary[5][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N967), 
        .Q(\inq_ary[5][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N967), 
        .Q(\inq_ary[5][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N967), 
        .Q(\inq_ary[5][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N967), 
        .Q(\inq_ary[5][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N967), 
        .Q(\inq_ary[5][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N967), 
        .Q(\inq_ary[5][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N967), 
        .Q(\inq_ary[5][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N967), 
        .Q(\inq_ary[5][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N967), 
        .Q(\inq_ary[5][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N967), 
        .Q(\inq_ary[5][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N967), 
        .Q(\inq_ary[5][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N967), 
        .Q(\inq_ary[5][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N967), 
        .Q(\inq_ary[5][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N967), 
        .Q(\inq_ary[5][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N967), 
        .Q(\inq_ary[5][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N967), 
        .Q(\inq_ary[5][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N967), 
        .Q(\inq_ary[5][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N967), 
        .Q(\inq_ary[5][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N967), 
        .Q(\inq_ary[5][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N967), 
        .Q(\inq_ary[5][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N967), 
        .Q(\inq_ary[5][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N967), 
        .Q(\inq_ary[5][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N967), 
        .Q(\inq_ary[5][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N967), 
        .Q(\inq_ary[5][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N967), 
        .Q(\inq_ary[5][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N967), 
        .Q(\inq_ary[5][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N967), 
        .Q(\inq_ary[5][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N967), 
        .Q(\inq_ary[5][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N967), 
        .Q(\inq_ary[5][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N967), 
        .Q(\inq_ary[5][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N967), 
        .Q(\inq_ary[5][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N967), 
        .Q(\inq_ary[5][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N967), 
        .Q(\inq_ary[5][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N967), 
        .Q(\inq_ary[5][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N967), 
        .Q(\inq_ary[5][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N967), 
        .Q(\inq_ary[5][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N967), 
        .Q(\inq_ary[5][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N967), 
        .Q(\inq_ary[5][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N967), 
        .Q(\inq_ary[5][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N967), 
        .Q(\inq_ary[5][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N967), 
        .Q(\inq_ary[5][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N967), 
        .Q(\inq_ary[5][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N967), 
        .Q(\inq_ary[5][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N967), 
        .Q(\inq_ary[5][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N967), .Q(
        \inq_ary[5][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N967), .Q(
        \inq_ary[5][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N967), .Q(
        \inq_ary[5][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N967), .Q(
        \inq_ary[5][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N967), .Q(
        \inq_ary[5][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N967), .Q(
        \inq_ary[5][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N967), .Q(
        \inq_ary[5][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N967), .Q(
        \inq_ary[5][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N967), .Q(
        \inq_ary[5][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[5][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N967), .Q(
        \inq_ary[5][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N966), 
        .Q(\inq_ary[4][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N966), 
        .Q(\inq_ary[4][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N966), 
        .Q(\inq_ary[4][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N966), 
        .Q(\inq_ary[4][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N966), 
        .Q(\inq_ary[4][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N966), 
        .Q(\inq_ary[4][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N966), 
        .Q(\inq_ary[4][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N966), 
        .Q(\inq_ary[4][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N966), 
        .Q(\inq_ary[4][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N966), 
        .Q(\inq_ary[4][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N966), 
        .Q(\inq_ary[4][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N966), 
        .Q(\inq_ary[4][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N966), 
        .Q(\inq_ary[4][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N966), 
        .Q(\inq_ary[4][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N966), 
        .Q(\inq_ary[4][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N966), 
        .Q(\inq_ary[4][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N966), 
        .Q(\inq_ary[4][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N966), 
        .Q(\inq_ary[4][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N966), 
        .Q(\inq_ary[4][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N966), 
        .Q(\inq_ary[4][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N966), 
        .Q(\inq_ary[4][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N966), 
        .Q(\inq_ary[4][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N966), 
        .Q(\inq_ary[4][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N966), 
        .Q(\inq_ary[4][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N966), 
        .Q(\inq_ary[4][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N966), 
        .Q(\inq_ary[4][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N966), 
        .Q(\inq_ary[4][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N966), 
        .Q(\inq_ary[4][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N966), 
        .Q(\inq_ary[4][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N966), 
        .Q(\inq_ary[4][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N966), 
        .Q(\inq_ary[4][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N966), 
        .Q(\inq_ary[4][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N966), 
        .Q(\inq_ary[4][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N966), 
        .Q(\inq_ary[4][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N966), 
        .Q(\inq_ary[4][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N966), 
        .Q(\inq_ary[4][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N966), 
        .Q(\inq_ary[4][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N966), 
        .Q(\inq_ary[4][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N966), 
        .Q(\inq_ary[4][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N966), 
        .Q(\inq_ary[4][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N966), 
        .Q(\inq_ary[4][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N966), 
        .Q(\inq_ary[4][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N966), 
        .Q(\inq_ary[4][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N966), 
        .Q(\inq_ary[4][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N966), 
        .Q(\inq_ary[4][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N966), 
        .Q(\inq_ary[4][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N966), 
        .Q(\inq_ary[4][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N966), 
        .Q(\inq_ary[4][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N966), 
        .Q(\inq_ary[4][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N966), 
        .Q(\inq_ary[4][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N966), 
        .Q(\inq_ary[4][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N966), 
        .Q(\inq_ary[4][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N966), 
        .Q(\inq_ary[4][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N966), 
        .Q(\inq_ary[4][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N966), 
        .Q(\inq_ary[4][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N966), 
        .Q(\inq_ary[4][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N966), 
        .Q(\inq_ary[4][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N966), 
        .Q(\inq_ary[4][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N966), 
        .Q(\inq_ary[4][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N966), 
        .Q(\inq_ary[4][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N966), 
        .Q(\inq_ary[4][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N965), 
        .Q(\inq_ary[4][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N965), 
        .Q(\inq_ary[4][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N965), 
        .Q(\inq_ary[4][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N965), 
        .Q(\inq_ary[4][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N965), 
        .Q(\inq_ary[4][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N965), 
        .Q(\inq_ary[4][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N965), 
        .Q(\inq_ary[4][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N965), 
        .Q(\inq_ary[4][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N965), 
        .Q(\inq_ary[4][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N965), 
        .Q(\inq_ary[4][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N965), 
        .Q(\inq_ary[4][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N965), 
        .Q(\inq_ary[4][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N965), 
        .Q(\inq_ary[4][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N965), 
        .Q(\inq_ary[4][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N965), 
        .Q(\inq_ary[4][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N965), 
        .Q(\inq_ary[4][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N965), 
        .Q(\inq_ary[4][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N965), 
        .Q(\inq_ary[4][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N965), 
        .Q(\inq_ary[4][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N965), 
        .Q(\inq_ary[4][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N965), 
        .Q(\inq_ary[4][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N965), 
        .Q(\inq_ary[4][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N965), 
        .Q(\inq_ary[4][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N965), 
        .Q(\inq_ary[4][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N965), 
        .Q(\inq_ary[4][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N965), 
        .Q(\inq_ary[4][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N965), 
        .Q(\inq_ary[4][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N965), 
        .Q(\inq_ary[4][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N965), 
        .Q(\inq_ary[4][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N965), 
        .Q(\inq_ary[4][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N965), 
        .Q(\inq_ary[4][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N965), 
        .Q(\inq_ary[4][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N965), 
        .Q(\inq_ary[4][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N965), 
        .Q(\inq_ary[4][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N965), 
        .Q(\inq_ary[4][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N965), 
        .Q(\inq_ary[4][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N965), 
        .Q(\inq_ary[4][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N965), 
        .Q(\inq_ary[4][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N965), 
        .Q(\inq_ary[4][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N965), 
        .Q(\inq_ary[4][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N965), 
        .Q(\inq_ary[4][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N965), 
        .Q(\inq_ary[4][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N965), 
        .Q(\inq_ary[4][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N965), 
        .Q(\inq_ary[4][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N965), 
        .Q(\inq_ary[4][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N965), 
        .Q(\inq_ary[4][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N965), 
        .Q(\inq_ary[4][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N965), 
        .Q(\inq_ary[4][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N965), 
        .Q(\inq_ary[4][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N965), 
        .Q(\inq_ary[4][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N965), 
        .Q(\inq_ary[4][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N965), 
        .Q(\inq_ary[4][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N965), 
        .Q(\inq_ary[4][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N965), 
        .Q(\inq_ary[4][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N965), 
        .Q(\inq_ary[4][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N965), 
        .Q(\inq_ary[4][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N965), 
        .Q(\inq_ary[4][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N965), 
        .Q(\inq_ary[4][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N965), 
        .Q(\inq_ary[4][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N965), 
        .Q(\inq_ary[4][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N965), 
        .Q(\inq_ary[4][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N965), 
        .Q(\inq_ary[4][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N965), 
        .Q(\inq_ary[4][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N965), 
        .Q(\inq_ary[4][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N965), 
        .Q(\inq_ary[4][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N965), 
        .Q(\inq_ary[4][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N965), 
        .Q(\inq_ary[4][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N965), 
        .Q(\inq_ary[4][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N965), 
        .Q(\inq_ary[4][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N965), 
        .Q(\inq_ary[4][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N965), 
        .Q(\inq_ary[4][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N965), 
        .Q(\inq_ary[4][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N965), 
        .Q(\inq_ary[4][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N965), 
        .Q(\inq_ary[4][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N965), 
        .Q(\inq_ary[4][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N965), 
        .Q(\inq_ary[4][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N965), 
        .Q(\inq_ary[4][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N965), 
        .Q(\inq_ary[4][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N965), 
        .Q(\inq_ary[4][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N965), 
        .Q(\inq_ary[4][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N965), 
        .Q(\inq_ary[4][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N965), 
        .Q(\inq_ary[4][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N965), 
        .Q(\inq_ary[4][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N965), 
        .Q(\inq_ary[4][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N965), 
        .Q(\inq_ary[4][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N965), 
        .Q(\inq_ary[4][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N965), 
        .Q(\inq_ary[4][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N965), 
        .Q(\inq_ary[4][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N965), 
        .Q(\inq_ary[4][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N965), .Q(
        \inq_ary[4][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N965), .Q(
        \inq_ary[4][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N965), .Q(
        \inq_ary[4][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N965), .Q(
        \inq_ary[4][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N965), .Q(
        \inq_ary[4][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N965), .Q(
        \inq_ary[4][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N965), .Q(
        \inq_ary[4][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N965), .Q(
        \inq_ary[4][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N965), .Q(
        \inq_ary[4][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[4][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N965), .Q(
        \inq_ary[4][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N964), 
        .Q(\inq_ary[3][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N964), 
        .Q(\inq_ary[3][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N964), 
        .Q(\inq_ary[3][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N964), 
        .Q(\inq_ary[3][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N964), 
        .Q(\inq_ary[3][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N964), 
        .Q(\inq_ary[3][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N964), 
        .Q(\inq_ary[3][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N964), 
        .Q(\inq_ary[3][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N964), 
        .Q(\inq_ary[3][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N964), 
        .Q(\inq_ary[3][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N964), 
        .Q(\inq_ary[3][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N964), 
        .Q(\inq_ary[3][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N964), 
        .Q(\inq_ary[3][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N964), 
        .Q(\inq_ary[3][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N964), 
        .Q(\inq_ary[3][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N964), 
        .Q(\inq_ary[3][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N964), 
        .Q(\inq_ary[3][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N964), 
        .Q(\inq_ary[3][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N964), 
        .Q(\inq_ary[3][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N964), 
        .Q(\inq_ary[3][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N964), 
        .Q(\inq_ary[3][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N964), 
        .Q(\inq_ary[3][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N964), 
        .Q(\inq_ary[3][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N964), 
        .Q(\inq_ary[3][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N964), 
        .Q(\inq_ary[3][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N964), 
        .Q(\inq_ary[3][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N964), 
        .Q(\inq_ary[3][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N964), 
        .Q(\inq_ary[3][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N964), 
        .Q(\inq_ary[3][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N964), 
        .Q(\inq_ary[3][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N964), 
        .Q(\inq_ary[3][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N964), 
        .Q(\inq_ary[3][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N964), 
        .Q(\inq_ary[3][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N964), 
        .Q(\inq_ary[3][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N964), 
        .Q(\inq_ary[3][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N964), 
        .Q(\inq_ary[3][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N964), 
        .Q(\inq_ary[3][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N964), 
        .Q(\inq_ary[3][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N964), 
        .Q(\inq_ary[3][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N964), 
        .Q(\inq_ary[3][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N964), 
        .Q(\inq_ary[3][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N964), 
        .Q(\inq_ary[3][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N964), 
        .Q(\inq_ary[3][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N964), 
        .Q(\inq_ary[3][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N964), 
        .Q(\inq_ary[3][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N964), 
        .Q(\inq_ary[3][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N964), 
        .Q(\inq_ary[3][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N964), 
        .Q(\inq_ary[3][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N964), 
        .Q(\inq_ary[3][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N964), 
        .Q(\inq_ary[3][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N964), 
        .Q(\inq_ary[3][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N964), 
        .Q(\inq_ary[3][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N964), 
        .Q(\inq_ary[3][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N964), 
        .Q(\inq_ary[3][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N964), 
        .Q(\inq_ary[3][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N964), 
        .Q(\inq_ary[3][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N964), 
        .Q(\inq_ary[3][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N964), 
        .Q(\inq_ary[3][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N964), 
        .Q(\inq_ary[3][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N964), 
        .Q(\inq_ary[3][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N964), 
        .Q(\inq_ary[3][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N963), 
        .Q(\inq_ary[3][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N963), 
        .Q(\inq_ary[3][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N963), 
        .Q(\inq_ary[3][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N963), 
        .Q(\inq_ary[3][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N963), 
        .Q(\inq_ary[3][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N963), 
        .Q(\inq_ary[3][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N963), 
        .Q(\inq_ary[3][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N963), 
        .Q(\inq_ary[3][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N963), 
        .Q(\inq_ary[3][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N963), 
        .Q(\inq_ary[3][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N963), 
        .Q(\inq_ary[3][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N963), 
        .Q(\inq_ary[3][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N963), 
        .Q(\inq_ary[3][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N963), 
        .Q(\inq_ary[3][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N963), 
        .Q(\inq_ary[3][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N963), 
        .Q(\inq_ary[3][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N963), 
        .Q(\inq_ary[3][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N963), 
        .Q(\inq_ary[3][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N963), 
        .Q(\inq_ary[3][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N963), 
        .Q(\inq_ary[3][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N963), 
        .Q(\inq_ary[3][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N963), 
        .Q(\inq_ary[3][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N963), 
        .Q(\inq_ary[3][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N963), 
        .Q(\inq_ary[3][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N963), 
        .Q(\inq_ary[3][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N963), 
        .Q(\inq_ary[3][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N963), 
        .Q(\inq_ary[3][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N963), 
        .Q(\inq_ary[3][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N963), 
        .Q(\inq_ary[3][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N963), 
        .Q(\inq_ary[3][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N963), 
        .Q(\inq_ary[3][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N963), 
        .Q(\inq_ary[3][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N963), 
        .Q(\inq_ary[3][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N963), 
        .Q(\inq_ary[3][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N963), 
        .Q(\inq_ary[3][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N963), 
        .Q(\inq_ary[3][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N963), 
        .Q(\inq_ary[3][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N963), 
        .Q(\inq_ary[3][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N963), 
        .Q(\inq_ary[3][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N963), 
        .Q(\inq_ary[3][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N963), 
        .Q(\inq_ary[3][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N963), 
        .Q(\inq_ary[3][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N963), 
        .Q(\inq_ary[3][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N963), 
        .Q(\inq_ary[3][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N963), 
        .Q(\inq_ary[3][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N963), 
        .Q(\inq_ary[3][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N963), 
        .Q(\inq_ary[3][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N963), 
        .Q(\inq_ary[3][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N963), 
        .Q(\inq_ary[3][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N963), 
        .Q(\inq_ary[3][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N963), 
        .Q(\inq_ary[3][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N963), 
        .Q(\inq_ary[3][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N963), 
        .Q(\inq_ary[3][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N963), 
        .Q(\inq_ary[3][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N963), 
        .Q(\inq_ary[3][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N963), 
        .Q(\inq_ary[3][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N963), 
        .Q(\inq_ary[3][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N963), 
        .Q(\inq_ary[3][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N963), 
        .Q(\inq_ary[3][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N963), 
        .Q(\inq_ary[3][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N963), 
        .Q(\inq_ary[3][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N963), 
        .Q(\inq_ary[3][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N963), 
        .Q(\inq_ary[3][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N963), 
        .Q(\inq_ary[3][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N963), 
        .Q(\inq_ary[3][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N963), 
        .Q(\inq_ary[3][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N963), 
        .Q(\inq_ary[3][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N963), 
        .Q(\inq_ary[3][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N963), 
        .Q(\inq_ary[3][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N963), 
        .Q(\inq_ary[3][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N963), 
        .Q(\inq_ary[3][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N963), 
        .Q(\inq_ary[3][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N963), 
        .Q(\inq_ary[3][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N963), 
        .Q(\inq_ary[3][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N963), 
        .Q(\inq_ary[3][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N963), 
        .Q(\inq_ary[3][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N963), 
        .Q(\inq_ary[3][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N963), 
        .Q(\inq_ary[3][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N963), 
        .Q(\inq_ary[3][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N963), 
        .Q(\inq_ary[3][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N963), 
        .Q(\inq_ary[3][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N963), 
        .Q(\inq_ary[3][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N963), 
        .Q(\inq_ary[3][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N963), 
        .Q(\inq_ary[3][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N963), 
        .Q(\inq_ary[3][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N963), 
        .Q(\inq_ary[3][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N963), 
        .Q(\inq_ary[3][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N963), 
        .Q(\inq_ary[3][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N963), 
        .Q(\inq_ary[3][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N963), .Q(
        \inq_ary[3][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N963), .Q(
        \inq_ary[3][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N963), .Q(
        \inq_ary[3][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N963), .Q(
        \inq_ary[3][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N963), .Q(
        \inq_ary[3][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N963), .Q(
        \inq_ary[3][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N963), .Q(
        \inq_ary[3][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N963), .Q(
        \inq_ary[3][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N963), .Q(
        \inq_ary[3][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[3][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N963), .Q(
        \inq_ary[3][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N962), 
        .Q(\inq_ary[2][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N962), 
        .Q(\inq_ary[2][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N962), 
        .Q(\inq_ary[2][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N962), 
        .Q(\inq_ary[2][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N962), 
        .Q(\inq_ary[2][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N962), 
        .Q(\inq_ary[2][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N962), 
        .Q(\inq_ary[2][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N962), 
        .Q(\inq_ary[2][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N962), 
        .Q(\inq_ary[2][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N962), 
        .Q(\inq_ary[2][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N962), 
        .Q(\inq_ary[2][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N962), 
        .Q(\inq_ary[2][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N962), 
        .Q(\inq_ary[2][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N962), 
        .Q(\inq_ary[2][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N962), 
        .Q(\inq_ary[2][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N962), 
        .Q(\inq_ary[2][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N962), 
        .Q(\inq_ary[2][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N962), 
        .Q(\inq_ary[2][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N962), 
        .Q(\inq_ary[2][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N962), 
        .Q(\inq_ary[2][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N962), 
        .Q(\inq_ary[2][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N962), 
        .Q(\inq_ary[2][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N962), 
        .Q(\inq_ary[2][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N962), 
        .Q(\inq_ary[2][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N962), 
        .Q(\inq_ary[2][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N962), 
        .Q(\inq_ary[2][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N962), 
        .Q(\inq_ary[2][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N962), 
        .Q(\inq_ary[2][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N962), 
        .Q(\inq_ary[2][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N962), 
        .Q(\inq_ary[2][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N962), 
        .Q(\inq_ary[2][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N962), 
        .Q(\inq_ary[2][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N962), 
        .Q(\inq_ary[2][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N962), 
        .Q(\inq_ary[2][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N962), 
        .Q(\inq_ary[2][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N962), 
        .Q(\inq_ary[2][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N962), 
        .Q(\inq_ary[2][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N962), 
        .Q(\inq_ary[2][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N962), 
        .Q(\inq_ary[2][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N962), 
        .Q(\inq_ary[2][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N962), 
        .Q(\inq_ary[2][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N962), 
        .Q(\inq_ary[2][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N962), 
        .Q(\inq_ary[2][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N962), 
        .Q(\inq_ary[2][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N962), 
        .Q(\inq_ary[2][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N962), 
        .Q(\inq_ary[2][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N962), 
        .Q(\inq_ary[2][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N962), 
        .Q(\inq_ary[2][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N962), 
        .Q(\inq_ary[2][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N962), 
        .Q(\inq_ary[2][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N962), 
        .Q(\inq_ary[2][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N962), 
        .Q(\inq_ary[2][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N962), 
        .Q(\inq_ary[2][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N962), 
        .Q(\inq_ary[2][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N962), 
        .Q(\inq_ary[2][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N962), 
        .Q(\inq_ary[2][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N962), 
        .Q(\inq_ary[2][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N962), 
        .Q(\inq_ary[2][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N962), 
        .Q(\inq_ary[2][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N962), 
        .Q(\inq_ary[2][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N962), 
        .Q(\inq_ary[2][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N961), 
        .Q(\inq_ary[2][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N961), 
        .Q(\inq_ary[2][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N961), 
        .Q(\inq_ary[2][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N961), 
        .Q(\inq_ary[2][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N961), 
        .Q(\inq_ary[2][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N961), 
        .Q(\inq_ary[2][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N961), 
        .Q(\inq_ary[2][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N961), 
        .Q(\inq_ary[2][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N961), 
        .Q(\inq_ary[2][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N961), 
        .Q(\inq_ary[2][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N961), 
        .Q(\inq_ary[2][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N961), 
        .Q(\inq_ary[2][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N961), 
        .Q(\inq_ary[2][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N961), 
        .Q(\inq_ary[2][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N961), 
        .Q(\inq_ary[2][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N961), 
        .Q(\inq_ary[2][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N961), 
        .Q(\inq_ary[2][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N961), 
        .Q(\inq_ary[2][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N961), 
        .Q(\inq_ary[2][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N961), 
        .Q(\inq_ary[2][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N961), 
        .Q(\inq_ary[2][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N961), 
        .Q(\inq_ary[2][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N961), 
        .Q(\inq_ary[2][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N961), 
        .Q(\inq_ary[2][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N961), 
        .Q(\inq_ary[2][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N961), 
        .Q(\inq_ary[2][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N961), 
        .Q(\inq_ary[2][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N961), 
        .Q(\inq_ary[2][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N961), 
        .Q(\inq_ary[2][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N961), 
        .Q(\inq_ary[2][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N961), 
        .Q(\inq_ary[2][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N961), 
        .Q(\inq_ary[2][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N961), 
        .Q(\inq_ary[2][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N961), 
        .Q(\inq_ary[2][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N961), 
        .Q(\inq_ary[2][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N961), 
        .Q(\inq_ary[2][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N961), 
        .Q(\inq_ary[2][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N961), 
        .Q(\inq_ary[2][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N961), 
        .Q(\inq_ary[2][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N961), 
        .Q(\inq_ary[2][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N961), 
        .Q(\inq_ary[2][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N961), 
        .Q(\inq_ary[2][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N961), 
        .Q(\inq_ary[2][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N961), 
        .Q(\inq_ary[2][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N961), 
        .Q(\inq_ary[2][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N961), 
        .Q(\inq_ary[2][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N961), 
        .Q(\inq_ary[2][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N961), 
        .Q(\inq_ary[2][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N961), 
        .Q(\inq_ary[2][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N961), 
        .Q(\inq_ary[2][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N961), 
        .Q(\inq_ary[2][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N961), 
        .Q(\inq_ary[2][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N961), 
        .Q(\inq_ary[2][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N961), 
        .Q(\inq_ary[2][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N961), 
        .Q(\inq_ary[2][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N961), 
        .Q(\inq_ary[2][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N961), 
        .Q(\inq_ary[2][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N961), 
        .Q(\inq_ary[2][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N961), 
        .Q(\inq_ary[2][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N961), 
        .Q(\inq_ary[2][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N961), 
        .Q(\inq_ary[2][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N961), 
        .Q(\inq_ary[2][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N961), 
        .Q(\inq_ary[2][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N961), 
        .Q(\inq_ary[2][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N961), 
        .Q(\inq_ary[2][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N961), 
        .Q(\inq_ary[2][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N961), 
        .Q(\inq_ary[2][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N961), 
        .Q(\inq_ary[2][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N961), 
        .Q(\inq_ary[2][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N961), 
        .Q(\inq_ary[2][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N961), 
        .Q(\inq_ary[2][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N961), 
        .Q(\inq_ary[2][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N961), 
        .Q(\inq_ary[2][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N961), 
        .Q(\inq_ary[2][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N961), 
        .Q(\inq_ary[2][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N961), 
        .Q(\inq_ary[2][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N961), 
        .Q(\inq_ary[2][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N961), 
        .Q(\inq_ary[2][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N961), 
        .Q(\inq_ary[2][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N961), 
        .Q(\inq_ary[2][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N961), 
        .Q(\inq_ary[2][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N961), 
        .Q(\inq_ary[2][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N961), 
        .Q(\inq_ary[2][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N961), 
        .Q(\inq_ary[2][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N961), 
        .Q(\inq_ary[2][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N961), 
        .Q(\inq_ary[2][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N961), 
        .Q(\inq_ary[2][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N961), 
        .Q(\inq_ary[2][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N961), 
        .Q(\inq_ary[2][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N961), .Q(
        \inq_ary[2][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N961), .Q(
        \inq_ary[2][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N961), .Q(
        \inq_ary[2][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N961), .Q(
        \inq_ary[2][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N961), .Q(
        \inq_ary[2][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N961), .Q(
        \inq_ary[2][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N961), .Q(
        \inq_ary[2][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N961), .Q(
        \inq_ary[2][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N961), .Q(
        \inq_ary[2][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[2][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N961), .Q(
        \inq_ary[2][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N960), 
        .Q(\inq_ary[1][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N960), 
        .Q(\inq_ary[1][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N960), 
        .Q(\inq_ary[1][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N960), 
        .Q(\inq_ary[1][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N960), 
        .Q(\inq_ary[1][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N960), 
        .Q(\inq_ary[1][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N960), 
        .Q(\inq_ary[1][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N960), 
        .Q(\inq_ary[1][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N960), 
        .Q(\inq_ary[1][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N960), 
        .Q(\inq_ary[1][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N960), 
        .Q(\inq_ary[1][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N960), 
        .Q(\inq_ary[1][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N960), 
        .Q(\inq_ary[1][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N960), 
        .Q(\inq_ary[1][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N960), 
        .Q(\inq_ary[1][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N960), 
        .Q(\inq_ary[1][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N960), 
        .Q(\inq_ary[1][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N960), 
        .Q(\inq_ary[1][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N960), 
        .Q(\inq_ary[1][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N960), 
        .Q(\inq_ary[1][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N960), 
        .Q(\inq_ary[1][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N960), 
        .Q(\inq_ary[1][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N960), 
        .Q(\inq_ary[1][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N960), 
        .Q(\inq_ary[1][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N960), 
        .Q(\inq_ary[1][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N960), 
        .Q(\inq_ary[1][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N960), 
        .Q(\inq_ary[1][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N960), 
        .Q(\inq_ary[1][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N960), 
        .Q(\inq_ary[1][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N960), 
        .Q(\inq_ary[1][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N960), 
        .Q(\inq_ary[1][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N960), 
        .Q(\inq_ary[1][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N960), 
        .Q(\inq_ary[1][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N960), 
        .Q(\inq_ary[1][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N960), 
        .Q(\inq_ary[1][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N960), 
        .Q(\inq_ary[1][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N960), 
        .Q(\inq_ary[1][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N960), 
        .Q(\inq_ary[1][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N960), 
        .Q(\inq_ary[1][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N960), 
        .Q(\inq_ary[1][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N960), 
        .Q(\inq_ary[1][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N960), 
        .Q(\inq_ary[1][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N960), 
        .Q(\inq_ary[1][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N960), 
        .Q(\inq_ary[1][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N960), 
        .Q(\inq_ary[1][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N960), 
        .Q(\inq_ary[1][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N960), 
        .Q(\inq_ary[1][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N960), 
        .Q(\inq_ary[1][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N960), 
        .Q(\inq_ary[1][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N960), 
        .Q(\inq_ary[1][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N960), 
        .Q(\inq_ary[1][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N960), 
        .Q(\inq_ary[1][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N960), 
        .Q(\inq_ary[1][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N960), 
        .Q(\inq_ary[1][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N960), 
        .Q(\inq_ary[1][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N960), 
        .Q(\inq_ary[1][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N960), 
        .Q(\inq_ary[1][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N960), 
        .Q(\inq_ary[1][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N960), 
        .Q(\inq_ary[1][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N960), 
        .Q(\inq_ary[1][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N960), 
        .Q(\inq_ary[1][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N959), 
        .Q(\inq_ary[1][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N959), 
        .Q(\inq_ary[1][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N959), 
        .Q(\inq_ary[1][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N959), 
        .Q(\inq_ary[1][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N959), 
        .Q(\inq_ary[1][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N959), 
        .Q(\inq_ary[1][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N959), 
        .Q(\inq_ary[1][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N959), 
        .Q(\inq_ary[1][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N959), 
        .Q(\inq_ary[1][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N959), 
        .Q(\inq_ary[1][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N959), 
        .Q(\inq_ary[1][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N959), 
        .Q(\inq_ary[1][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N959), 
        .Q(\inq_ary[1][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N959), 
        .Q(\inq_ary[1][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N959), 
        .Q(\inq_ary[1][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N959), 
        .Q(\inq_ary[1][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N959), 
        .Q(\inq_ary[1][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N959), 
        .Q(\inq_ary[1][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N959), 
        .Q(\inq_ary[1][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N959), 
        .Q(\inq_ary[1][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N959), 
        .Q(\inq_ary[1][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N959), 
        .Q(\inq_ary[1][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N959), 
        .Q(\inq_ary[1][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N959), 
        .Q(\inq_ary[1][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N959), 
        .Q(\inq_ary[1][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N959), 
        .Q(\inq_ary[1][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N959), 
        .Q(\inq_ary[1][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N959), 
        .Q(\inq_ary[1][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N959), 
        .Q(\inq_ary[1][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N959), 
        .Q(\inq_ary[1][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N959), 
        .Q(\inq_ary[1][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N959), 
        .Q(\inq_ary[1][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N959), 
        .Q(\inq_ary[1][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N959), 
        .Q(\inq_ary[1][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N959), 
        .Q(\inq_ary[1][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N959), 
        .Q(\inq_ary[1][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N959), 
        .Q(\inq_ary[1][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N959), 
        .Q(\inq_ary[1][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N959), 
        .Q(\inq_ary[1][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N959), 
        .Q(\inq_ary[1][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N959), 
        .Q(\inq_ary[1][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N959), 
        .Q(\inq_ary[1][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N959), 
        .Q(\inq_ary[1][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N959), 
        .Q(\inq_ary[1][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N959), 
        .Q(\inq_ary[1][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N959), 
        .Q(\inq_ary[1][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N959), 
        .Q(\inq_ary[1][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N959), 
        .Q(\inq_ary[1][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N959), 
        .Q(\inq_ary[1][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N959), 
        .Q(\inq_ary[1][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N959), 
        .Q(\inq_ary[1][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N959), 
        .Q(\inq_ary[1][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N959), 
        .Q(\inq_ary[1][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N959), 
        .Q(\inq_ary[1][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N959), 
        .Q(\inq_ary[1][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N959), 
        .Q(\inq_ary[1][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N959), 
        .Q(\inq_ary[1][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N959), 
        .Q(\inq_ary[1][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N959), 
        .Q(\inq_ary[1][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N959), 
        .Q(\inq_ary[1][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N959), 
        .Q(\inq_ary[1][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N959), 
        .Q(\inq_ary[1][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N959), 
        .Q(\inq_ary[1][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N959), 
        .Q(\inq_ary[1][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N959), 
        .Q(\inq_ary[1][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N959), 
        .Q(\inq_ary[1][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N959), 
        .Q(\inq_ary[1][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N959), 
        .Q(\inq_ary[1][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N959), 
        .Q(\inq_ary[1][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N959), 
        .Q(\inq_ary[1][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N959), 
        .Q(\inq_ary[1][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N959), 
        .Q(\inq_ary[1][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N959), 
        .Q(\inq_ary[1][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N959), 
        .Q(\inq_ary[1][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N959), 
        .Q(\inq_ary[1][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N959), 
        .Q(\inq_ary[1][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N959), 
        .Q(\inq_ary[1][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N959), 
        .Q(\inq_ary[1][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N959), 
        .Q(\inq_ary[1][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N959), 
        .Q(\inq_ary[1][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N959), 
        .Q(\inq_ary[1][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N959), 
        .Q(\inq_ary[1][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N959), 
        .Q(\inq_ary[1][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N959), 
        .Q(\inq_ary[1][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N959), 
        .Q(\inq_ary[1][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N959), 
        .Q(\inq_ary[1][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N959), 
        .Q(\inq_ary[1][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N959), 
        .Q(\inq_ary[1][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N959), 
        .Q(\inq_ary[1][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N959), .Q(
        \inq_ary[1][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N959), .Q(
        \inq_ary[1][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N959), .Q(
        \inq_ary[1][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N959), .Q(
        \inq_ary[1][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N959), .Q(
        \inq_ary[1][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N959), .Q(
        \inq_ary[1][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N959), .Q(
        \inq_ary[1][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N959), .Q(
        \inq_ary[1][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N959), .Q(
        \inq_ary[1][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[1][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N959), .Q(
        \inq_ary[1][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][159]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N908), .enable(N958), 
        .Q(\inq_ary[0][159] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][158]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N907), .enable(N958), 
        .Q(\inq_ary[0][158] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][157]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N906), .enable(N958), 
        .Q(\inq_ary[0][157] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][156]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N905), .enable(N958), 
        .Q(\inq_ary[0][156] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][155]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N904), .enable(N958), 
        .Q(\inq_ary[0][155] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][154]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N901), .enable(N958), 
        .Q(\inq_ary[0][154] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][153]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N898), .enable(N958), 
        .Q(\inq_ary[0][153] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][152]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N895), .enable(N958), 
        .Q(\inq_ary[0][152] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][151]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N892), .enable(N958), 
        .Q(\inq_ary[0][151] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][150]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N891), .enable(N958), 
        .Q(\inq_ary[0][150] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][149]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N890), .enable(N958), 
        .Q(\inq_ary[0][149] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][148]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N889), .enable(N958), 
        .Q(\inq_ary[0][148] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][147]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N888), .enable(N958), 
        .Q(\inq_ary[0][147] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][146]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N885), .enable(N958), 
        .Q(\inq_ary[0][146] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][145]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N882), .enable(N958), 
        .Q(\inq_ary[0][145] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][144]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N879), .enable(N958), 
        .Q(\inq_ary[0][144] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][143]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N876), .enable(N958), 
        .Q(\inq_ary[0][143] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][142]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N875), .enable(N958), 
        .Q(\inq_ary[0][142] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][141]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N874), .enable(N958), 
        .Q(\inq_ary[0][141] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][140]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N873), .enable(N958), 
        .Q(\inq_ary[0][140] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][139]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N872), .enable(N958), 
        .Q(\inq_ary[0][139] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][138]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N869), .enable(N958), 
        .Q(\inq_ary[0][138] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][137]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N866), .enable(N958), 
        .Q(\inq_ary[0][137] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][136]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N863), .enable(N958), 
        .Q(\inq_ary[0][136] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][135]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N860), .enable(N958), 
        .Q(\inq_ary[0][135] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][134]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N859), .enable(N958), 
        .Q(\inq_ary[0][134] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][133]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N858), .enable(N958), 
        .Q(\inq_ary[0][133] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][132]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N857), .enable(N958), 
        .Q(\inq_ary[0][132] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][131]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N856), .enable(N958), 
        .Q(\inq_ary[0][131] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][130]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N853), .enable(N958), 
        .Q(\inq_ary[0][130] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][129]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N850), .enable(N958), 
        .Q(\inq_ary[0][129] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][128]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N847), .enable(N958), 
        .Q(\inq_ary[0][128] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][127]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N844), .enable(N958), 
        .Q(\inq_ary[0][127] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][126]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N843), .enable(N958), 
        .Q(\inq_ary[0][126] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][125]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N842), .enable(N958), 
        .Q(\inq_ary[0][125] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][124]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N841), .enable(N958), 
        .Q(\inq_ary[0][124] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][123]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N840), .enable(N958), 
        .Q(\inq_ary[0][123] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][122]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N837), .enable(N958), 
        .Q(\inq_ary[0][122] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][121]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N834), .enable(N958), 
        .Q(\inq_ary[0][121] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][120]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N831), .enable(N958), 
        .Q(\inq_ary[0][120] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][119]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N828), .enable(N958), 
        .Q(\inq_ary[0][119] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][118]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N827), .enable(N958), 
        .Q(\inq_ary[0][118] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][117]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N826), .enable(N958), 
        .Q(\inq_ary[0][117] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][116]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N825), .enable(N958), 
        .Q(\inq_ary[0][116] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][115]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N824), .enable(N958), 
        .Q(\inq_ary[0][115] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][114]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N821), .enable(N958), 
        .Q(\inq_ary[0][114] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][113]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N818), .enable(N958), 
        .Q(\inq_ary[0][113] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][112]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N815), .enable(N958), 
        .Q(\inq_ary[0][112] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][111]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N812), .enable(N958), 
        .Q(\inq_ary[0][111] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][110]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N811), .enable(N958), 
        .Q(\inq_ary[0][110] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][109]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N810), .enable(N958), 
        .Q(\inq_ary[0][109] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][108]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N809), .enable(N958), 
        .Q(\inq_ary[0][108] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][107]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N808), .enable(N958), 
        .Q(\inq_ary[0][107] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][106]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N805), .enable(N958), 
        .Q(\inq_ary[0][106] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][105]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N802), .enable(N958), 
        .Q(\inq_ary[0][105] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][104]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N799), .enable(N958), 
        .Q(\inq_ary[0][104] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][103]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N796), .enable(N958), 
        .Q(\inq_ary[0][103] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][102]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N795), .enable(N958), 
        .Q(\inq_ary[0][102] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][101]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N794), .enable(N958), 
        .Q(\inq_ary[0][101] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][100]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N793), .enable(N958), 
        .Q(\inq_ary[0][100] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][99]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N792), .enable(N958), 
        .Q(\inq_ary[0][99] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][98]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N789), .enable(N957), 
        .Q(\inq_ary[0][98] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][97]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N786), .enable(N957), 
        .Q(\inq_ary[0][97] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][96]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N783), .enable(N957), 
        .Q(\inq_ary[0][96] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][95]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N780), .enable(N957), 
        .Q(\inq_ary[0][95] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][94]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N779), .enable(N957), 
        .Q(\inq_ary[0][94] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][93]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N778), .enable(N957), 
        .Q(\inq_ary[0][93] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][92]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N777), .enable(N957), 
        .Q(\inq_ary[0][92] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][91]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N776), .enable(N957), 
        .Q(\inq_ary[0][91] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][90]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N773), .enable(N957), 
        .Q(\inq_ary[0][90] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][89]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N770), .enable(N957), 
        .Q(\inq_ary[0][89] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][88]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N767), .enable(N957), 
        .Q(\inq_ary[0][88] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][87]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N764), .enable(N957), 
        .Q(\inq_ary[0][87] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][86]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N763), .enable(N957), 
        .Q(\inq_ary[0][86] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][85]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N762), .enable(N957), 
        .Q(\inq_ary[0][85] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][84]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N761), .enable(N957), 
        .Q(\inq_ary[0][84] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][83]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N760), .enable(N957), 
        .Q(\inq_ary[0][83] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][82]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N757), .enable(N957), 
        .Q(\inq_ary[0][82] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][81]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N754), .enable(N957), 
        .Q(\inq_ary[0][81] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][80]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N751), .enable(N957), 
        .Q(\inq_ary[0][80] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][79]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N748), .enable(N957), 
        .Q(\inq_ary[0][79] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][78]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N747), .enable(N957), 
        .Q(\inq_ary[0][78] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][77]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N746), .enable(N957), 
        .Q(\inq_ary[0][77] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][76]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N745), .enable(N957), 
        .Q(\inq_ary[0][76] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][75]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N744), .enable(N957), 
        .Q(\inq_ary[0][75] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][74]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N741), .enable(N957), 
        .Q(\inq_ary[0][74] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][73]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N738), .enable(N957), 
        .Q(\inq_ary[0][73] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][72]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N735), .enable(N957), 
        .Q(\inq_ary[0][72] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][71]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N732), .enable(N957), 
        .Q(\inq_ary[0][71] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][70]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N731), .enable(N957), 
        .Q(\inq_ary[0][70] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][69]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N730), .enable(N957), 
        .Q(\inq_ary[0][69] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][68]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N729), .enable(N957), 
        .Q(\inq_ary[0][68] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][67]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N728), .enable(N957), 
        .Q(\inq_ary[0][67] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][66]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N725), .enable(N957), 
        .Q(\inq_ary[0][66] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][65]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N722), .enable(N957), 
        .Q(\inq_ary[0][65] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][64]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N719), .enable(N957), 
        .Q(\inq_ary[0][64] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][63]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N716), .enable(N957), 
        .Q(\inq_ary[0][63] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][62]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N715), .enable(N957), 
        .Q(\inq_ary[0][62] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][61]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N714), .enable(N957), 
        .Q(\inq_ary[0][61] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][60]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N713), .enable(N957), 
        .Q(\inq_ary[0][60] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][59]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N712), .enable(N957), 
        .Q(\inq_ary[0][59] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][58]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N709), .enable(N957), 
        .Q(\inq_ary[0][58] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][57]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N706), .enable(N957), 
        .Q(\inq_ary[0][57] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][56]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N703), .enable(N957), 
        .Q(\inq_ary[0][56] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][55]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N700), .enable(N957), 
        .Q(\inq_ary[0][55] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][54]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N699), .enable(N957), 
        .Q(\inq_ary[0][54] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][53]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N698), .enable(N957), 
        .Q(\inq_ary[0][53] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][52]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N697), .enable(N957), 
        .Q(\inq_ary[0][52] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][51]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N696), .enable(N957), 
        .Q(\inq_ary[0][51] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][50]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N693), .enable(N957), 
        .Q(\inq_ary[0][50] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][49]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N690), .enable(N957), 
        .Q(\inq_ary[0][49] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][48]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N687), .enable(N957), 
        .Q(\inq_ary[0][48] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][47]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N684), .enable(N957), 
        .Q(\inq_ary[0][47] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][46]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N683), .enable(N957), 
        .Q(\inq_ary[0][46] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][45]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N682), .enable(N957), 
        .Q(\inq_ary[0][45] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][44]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N681), .enable(N957), 
        .Q(\inq_ary[0][44] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][43]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N680), .enable(N957), 
        .Q(\inq_ary[0][43] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][42]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N677), .enable(N957), 
        .Q(\inq_ary[0][42] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][41]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N674), .enable(N957), 
        .Q(\inq_ary[0][41] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][40]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N671), .enable(N957), 
        .Q(\inq_ary[0][40] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][39]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N668), .enable(N957), 
        .Q(\inq_ary[0][39] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][38]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N667), .enable(N957), 
        .Q(\inq_ary[0][38] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][37]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N666), .enable(N957), 
        .Q(\inq_ary[0][37] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][36]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N665), .enable(N957), 
        .Q(\inq_ary[0][36] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][35]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N664), .enable(N957), 
        .Q(\inq_ary[0][35] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][34]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N661), .enable(N957), 
        .Q(\inq_ary[0][34] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][33]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N658), .enable(N957), 
        .Q(\inq_ary[0][33] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][32]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N655), .enable(N957), 
        .Q(\inq_ary[0][32] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][31]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N652), .enable(N957), 
        .Q(\inq_ary[0][31] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][30]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N651), .enable(N957), 
        .Q(\inq_ary[0][30] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][29]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N650), .enable(N957), 
        .Q(\inq_ary[0][29] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][28]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N649), .enable(N957), 
        .Q(\inq_ary[0][28] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][27]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N648), .enable(N957), 
        .Q(\inq_ary[0][27] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][26]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N645), .enable(N957), 
        .Q(\inq_ary[0][26] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][25]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N642), .enable(N957), 
        .Q(\inq_ary[0][25] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][24]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N639), .enable(N957), 
        .Q(\inq_ary[0][24] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][23]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N636), .enable(N957), 
        .Q(\inq_ary[0][23] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][22]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N635), .enable(N957), 
        .Q(\inq_ary[0][22] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][21]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N634), .enable(N957), 
        .Q(\inq_ary[0][21] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][20]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N633), .enable(N957), 
        .Q(\inq_ary[0][20] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][19]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N632), .enable(N957), 
        .Q(\inq_ary[0][19] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][18]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N629), .enable(N957), 
        .Q(\inq_ary[0][18] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][17]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N626), .enable(N957), 
        .Q(\inq_ary[0][17] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][16]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N623), .enable(N957), 
        .Q(\inq_ary[0][16] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][15]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N620), .enable(N957), 
        .Q(\inq_ary[0][15] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][14]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N619), .enable(N957), 
        .Q(\inq_ary[0][14] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][13]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N618), .enable(N957), 
        .Q(\inq_ary[0][13] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][12]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N617), .enable(N957), 
        .Q(\inq_ary[0][12] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][11]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N616), .enable(N957), 
        .Q(\inq_ary[0][11] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][10]  ( .clear(1'b0), .preset(1'b0), 
        .next_state(1'b0), .clocked_on(1'b0), .data_in(N613), .enable(N957), 
        .Q(\inq_ary[0][10] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N610), .enable(N957), .Q(
        \inq_ary[0][9] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N607), .enable(N957), .Q(
        \inq_ary[0][8] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N604), .enable(N957), .Q(
        \inq_ary[0][7] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N603), .enable(N957), .Q(
        \inq_ary[0][6] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N602), .enable(N957), .Q(
        \inq_ary[0][5] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N601), .enable(N957), .Q(
        \inq_ary[0][4] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N600), .enable(N957), .Q(
        \inq_ary[0][3] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N597), .enable(N957), .Q(
        \inq_ary[0][2] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N594), .enable(N957), .Q(
        \inq_ary[0][1] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  \**SEQGEN**  \inq_ary_reg[0][0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        1'b0), .clocked_on(1'b0), .data_in(N591), .enable(N957), .Q(
        \inq_ary[0][0] ), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b0) );
  GTECH_AND2 C24306 ( .A(wrptr_d1[2]), .B(wrptr_d1[3]), .Z(N990) );
  GTECH_AND2 C24307 ( .A(N0), .B(wrptr_d1[3]), .Z(N991) );
  GTECH_NOT I_0 ( .A(wrptr_d1[2]), .Z(N0) );
  GTECH_AND2 C24308 ( .A(wrptr_d1[2]), .B(N1), .Z(N992) );
  GTECH_NOT I_1 ( .A(wrptr_d1[3]), .Z(N1) );
  GTECH_AND2 C24309 ( .A(N2), .B(N3), .Z(N993) );
  GTECH_NOT I_2 ( .A(wrptr_d1[2]), .Z(N2) );
  GTECH_NOT I_3 ( .A(wrptr_d1[3]), .Z(N3) );
  GTECH_AND2 C24310 ( .A(wrptr_d1[0]), .B(wrptr_d1[1]), .Z(N994) );
  GTECH_AND2 C24311 ( .A(N4), .B(wrptr_d1[1]), .Z(N995) );
  GTECH_NOT I_4 ( .A(wrptr_d1[0]), .Z(N4) );
  GTECH_AND2 C24312 ( .A(wrptr_d1[0]), .B(N5), .Z(N996) );
  GTECH_NOT I_5 ( .A(wrptr_d1[1]), .Z(N5) );
  GTECH_AND2 C24313 ( .A(N6), .B(N7), .Z(N997) );
  GTECH_NOT I_6 ( .A(wrptr_d1[0]), .Z(N6) );
  GTECH_NOT I_7 ( .A(wrptr_d1[1]), .Z(N7) );
  GTECH_AND2 C24314 ( .A(N990), .B(N994), .Z(N924) );
  GTECH_AND2 C24315 ( .A(N990), .B(N995), .Z(N923) );
  GTECH_AND2 C24316 ( .A(N990), .B(N996), .Z(N922) );
  GTECH_AND2 C24317 ( .A(N990), .B(N997), .Z(N921) );
  GTECH_AND2 C24318 ( .A(N991), .B(N994), .Z(N920) );
  GTECH_AND2 C24319 ( .A(N991), .B(N995), .Z(N919) );
  GTECH_AND2 C24320 ( .A(N991), .B(N996), .Z(N918) );
  GTECH_AND2 C24321 ( .A(N991), .B(N997), .Z(N917) );
  GTECH_AND2 C24322 ( .A(N992), .B(N994), .Z(N916) );
  GTECH_AND2 C24323 ( .A(N992), .B(N995), .Z(N915) );
  GTECH_AND2 C24324 ( .A(N992), .B(N996), .Z(N914) );
  GTECH_AND2 C24325 ( .A(N992), .B(N997), .Z(N913) );
  GTECH_AND2 C24326 ( .A(N993), .B(N994), .Z(N912) );
  GTECH_AND2 C24327 ( .A(N993), .B(N995), .Z(N911) );
  GTECH_AND2 C24328 ( .A(N993), .B(N996), .Z(N910) );
  GTECH_AND2 C24329 ( .A(N993), .B(N997), .Z(N909) );
  SELECT_OP C24906 ( .DATA1({ren_d1, ren_d1}), .DATA2({1'b1, 1'b1}), 
        .CONTROL1(N8), .CONTROL2(N9), .Z({N360, N260}) );
  GTECH_BUF B_0 ( .A(reset_l), .Z(N8) );
  GTECH_BUF B_1 ( .A(N259), .Z(N9) );
  SELECT_OP C24907 ( .DATA1({N99, N100, N101, N102, N103, N104, N105, N106, 
        N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, 
        N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, 
        N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, 
        N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, 
        N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, 
        N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, 
        N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
        N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
        N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
        N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, 
        N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
        N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, 
        N251, N252, N253, N254, N255, N256, N257, N258}), .DATA2({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CONTROL1(N8), .CONTROL2(N9), .Z({N421, N420, N419, N418, 
        N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, 
        N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, 
        N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, 
        N369, N368, N367, N366, N365, N364, N363, N362, N361, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261}) );
  SELECT_OP C24908 ( .DATA1(wrdata_d1[0]), .DATA2(N581), .CONTROL1(N10), 
        .CONTROL2(N590), .Z(N591) );
  GTECH_BUF B_2 ( .A(N589), .Z(N10) );
  SELECT_OP C24909 ( .DATA1(wrdata_d1[1]), .DATA2(N580), .CONTROL1(N11), 
        .CONTROL2(N593), .Z(N594) );
  GTECH_BUF B_3 ( .A(N592), .Z(N11) );
  SELECT_OP C24910 ( .DATA1(wrdata_d1[2]), .DATA2(N579), .CONTROL1(N12), 
        .CONTROL2(N596), .Z(N597) );
  GTECH_BUF B_4 ( .A(N595), .Z(N12) );
  SELECT_OP C24911 ( .DATA1(wrdata_d1[3]), .DATA2(N578), .CONTROL1(N13), 
        .CONTROL2(N599), .Z(N600) );
  GTECH_BUF B_5 ( .A(N598), .Z(N13) );
  SELECT_OP C24912 ( .DATA1(wrdata_d1[4]), .DATA2(N577), .CONTROL1(N10), 
        .CONTROL2(N590), .Z(N601) );
  SELECT_OP C24913 ( .DATA1(wrdata_d1[5]), .DATA2(N576), .CONTROL1(N11), 
        .CONTROL2(N593), .Z(N602) );
  SELECT_OP C24914 ( .DATA1(wrdata_d1[6]), .DATA2(N575), .CONTROL1(N12), 
        .CONTROL2(N596), .Z(N603) );
  SELECT_OP C24915 ( .DATA1(wrdata_d1[7]), .DATA2(N574), .CONTROL1(N13), 
        .CONTROL2(N599), .Z(N604) );
  SELECT_OP C24916 ( .DATA1(wrdata_d1[8]), .DATA2(N573), .CONTROL1(N14), 
        .CONTROL2(N606), .Z(N607) );
  GTECH_BUF B_6 ( .A(N605), .Z(N14) );
  SELECT_OP C24917 ( .DATA1(wrdata_d1[9]), .DATA2(N572), .CONTROL1(N15), 
        .CONTROL2(N609), .Z(N610) );
  GTECH_BUF B_7 ( .A(N608), .Z(N15) );
  SELECT_OP C24918 ( .DATA1(wrdata_d1[10]), .DATA2(N571), .CONTROL1(N16), 
        .CONTROL2(N612), .Z(N613) );
  GTECH_BUF B_8 ( .A(N611), .Z(N16) );
  SELECT_OP C24919 ( .DATA1(wrdata_d1[11]), .DATA2(N570), .CONTROL1(N17), 
        .CONTROL2(N615), .Z(N616) );
  GTECH_BUF B_9 ( .A(N614), .Z(N17) );
  SELECT_OP C24920 ( .DATA1(wrdata_d1[12]), .DATA2(N569), .CONTROL1(N14), 
        .CONTROL2(N606), .Z(N617) );
  SELECT_OP C24921 ( .DATA1(wrdata_d1[13]), .DATA2(N568), .CONTROL1(N15), 
        .CONTROL2(N609), .Z(N618) );
  SELECT_OP C24922 ( .DATA1(wrdata_d1[14]), .DATA2(N567), .CONTROL1(N16), 
        .CONTROL2(N612), .Z(N619) );
  SELECT_OP C24923 ( .DATA1(wrdata_d1[15]), .DATA2(N566), .CONTROL1(N17), 
        .CONTROL2(N615), .Z(N620) );
  SELECT_OP C24924 ( .DATA1(wrdata_d1[16]), .DATA2(N565), .CONTROL1(N18), 
        .CONTROL2(N622), .Z(N623) );
  GTECH_BUF B_10 ( .A(N621), .Z(N18) );
  SELECT_OP C24925 ( .DATA1(wrdata_d1[17]), .DATA2(N564), .CONTROL1(N19), 
        .CONTROL2(N625), .Z(N626) );
  GTECH_BUF B_11 ( .A(N624), .Z(N19) );
  SELECT_OP C24926 ( .DATA1(wrdata_d1[18]), .DATA2(N563), .CONTROL1(N20), 
        .CONTROL2(N628), .Z(N629) );
  GTECH_BUF B_12 ( .A(N627), .Z(N20) );
  SELECT_OP C24927 ( .DATA1(wrdata_d1[19]), .DATA2(N562), .CONTROL1(N21), 
        .CONTROL2(N631), .Z(N632) );
  GTECH_BUF B_13 ( .A(N630), .Z(N21) );
  SELECT_OP C24928 ( .DATA1(wrdata_d1[20]), .DATA2(N561), .CONTROL1(N18), 
        .CONTROL2(N622), .Z(N633) );
  SELECT_OP C24929 ( .DATA1(wrdata_d1[21]), .DATA2(N560), .CONTROL1(N19), 
        .CONTROL2(N625), .Z(N634) );
  SELECT_OP C24930 ( .DATA1(wrdata_d1[22]), .DATA2(N559), .CONTROL1(N20), 
        .CONTROL2(N628), .Z(N635) );
  SELECT_OP C24931 ( .DATA1(wrdata_d1[23]), .DATA2(N558), .CONTROL1(N21), 
        .CONTROL2(N631), .Z(N636) );
  SELECT_OP C24932 ( .DATA1(wrdata_d1[24]), .DATA2(N557), .CONTROL1(N22), 
        .CONTROL2(N638), .Z(N639) );
  GTECH_BUF B_14 ( .A(N637), .Z(N22) );
  SELECT_OP C24933 ( .DATA1(wrdata_d1[25]), .DATA2(N556), .CONTROL1(N23), 
        .CONTROL2(N641), .Z(N642) );
  GTECH_BUF B_15 ( .A(N640), .Z(N23) );
  SELECT_OP C24934 ( .DATA1(wrdata_d1[26]), .DATA2(N555), .CONTROL1(N24), 
        .CONTROL2(N644), .Z(N645) );
  GTECH_BUF B_16 ( .A(N643), .Z(N24) );
  SELECT_OP C24935 ( .DATA1(wrdata_d1[27]), .DATA2(N554), .CONTROL1(N25), 
        .CONTROL2(N647), .Z(N648) );
  GTECH_BUF B_17 ( .A(N646), .Z(N25) );
  SELECT_OP C24936 ( .DATA1(wrdata_d1[28]), .DATA2(N553), .CONTROL1(N22), 
        .CONTROL2(N638), .Z(N649) );
  SELECT_OP C24937 ( .DATA1(wrdata_d1[29]), .DATA2(N552), .CONTROL1(N23), 
        .CONTROL2(N641), .Z(N650) );
  SELECT_OP C24938 ( .DATA1(wrdata_d1[30]), .DATA2(N551), .CONTROL1(N24), 
        .CONTROL2(N644), .Z(N651) );
  SELECT_OP C24939 ( .DATA1(wrdata_d1[31]), .DATA2(N550), .CONTROL1(N25), 
        .CONTROL2(N647), .Z(N652) );
  SELECT_OP C24940 ( .DATA1(wrdata_d1[32]), .DATA2(N549), .CONTROL1(N26), 
        .CONTROL2(N654), .Z(N655) );
  GTECH_BUF B_18 ( .A(N653), .Z(N26) );
  SELECT_OP C24941 ( .DATA1(wrdata_d1[33]), .DATA2(N548), .CONTROL1(N27), 
        .CONTROL2(N657), .Z(N658) );
  GTECH_BUF B_19 ( .A(N656), .Z(N27) );
  SELECT_OP C24942 ( .DATA1(wrdata_d1[34]), .DATA2(N547), .CONTROL1(N28), 
        .CONTROL2(N660), .Z(N661) );
  GTECH_BUF B_20 ( .A(N659), .Z(N28) );
  SELECT_OP C24943 ( .DATA1(wrdata_d1[35]), .DATA2(N546), .CONTROL1(N29), 
        .CONTROL2(N663), .Z(N664) );
  GTECH_BUF B_21 ( .A(N662), .Z(N29) );
  SELECT_OP C24944 ( .DATA1(wrdata_d1[36]), .DATA2(N545), .CONTROL1(N26), 
        .CONTROL2(N654), .Z(N665) );
  SELECT_OP C24945 ( .DATA1(wrdata_d1[37]), .DATA2(N544), .CONTROL1(N27), 
        .CONTROL2(N657), .Z(N666) );
  SELECT_OP C24946 ( .DATA1(wrdata_d1[38]), .DATA2(N543), .CONTROL1(N28), 
        .CONTROL2(N660), .Z(N667) );
  SELECT_OP C24947 ( .DATA1(wrdata_d1[39]), .DATA2(N542), .CONTROL1(N29), 
        .CONTROL2(N663), .Z(N668) );
  SELECT_OP C24948 ( .DATA1(wrdata_d1[40]), .DATA2(N541), .CONTROL1(N30), 
        .CONTROL2(N670), .Z(N671) );
  GTECH_BUF B_22 ( .A(N669), .Z(N30) );
  SELECT_OP C24949 ( .DATA1(wrdata_d1[41]), .DATA2(N540), .CONTROL1(N31), 
        .CONTROL2(N673), .Z(N674) );
  GTECH_BUF B_23 ( .A(N672), .Z(N31) );
  SELECT_OP C24950 ( .DATA1(wrdata_d1[42]), .DATA2(N539), .CONTROL1(N32), 
        .CONTROL2(N676), .Z(N677) );
  GTECH_BUF B_24 ( .A(N675), .Z(N32) );
  SELECT_OP C24951 ( .DATA1(wrdata_d1[43]), .DATA2(N538), .CONTROL1(N33), 
        .CONTROL2(N679), .Z(N680) );
  GTECH_BUF B_25 ( .A(N678), .Z(N33) );
  SELECT_OP C24952 ( .DATA1(wrdata_d1[44]), .DATA2(N537), .CONTROL1(N30), 
        .CONTROL2(N670), .Z(N681) );
  SELECT_OP C24953 ( .DATA1(wrdata_d1[45]), .DATA2(N536), .CONTROL1(N31), 
        .CONTROL2(N673), .Z(N682) );
  SELECT_OP C24954 ( .DATA1(wrdata_d1[46]), .DATA2(N535), .CONTROL1(N32), 
        .CONTROL2(N676), .Z(N683) );
  SELECT_OP C24955 ( .DATA1(wrdata_d1[47]), .DATA2(N534), .CONTROL1(N33), 
        .CONTROL2(N679), .Z(N684) );
  SELECT_OP C24956 ( .DATA1(wrdata_d1[48]), .DATA2(N533), .CONTROL1(N34), 
        .CONTROL2(N686), .Z(N687) );
  GTECH_BUF B_26 ( .A(N685), .Z(N34) );
  SELECT_OP C24957 ( .DATA1(wrdata_d1[49]), .DATA2(N532), .CONTROL1(N35), 
        .CONTROL2(N689), .Z(N690) );
  GTECH_BUF B_27 ( .A(N688), .Z(N35) );
  SELECT_OP C24958 ( .DATA1(wrdata_d1[50]), .DATA2(N531), .CONTROL1(N36), 
        .CONTROL2(N692), .Z(N693) );
  GTECH_BUF B_28 ( .A(N691), .Z(N36) );
  SELECT_OP C24959 ( .DATA1(wrdata_d1[51]), .DATA2(N530), .CONTROL1(N37), 
        .CONTROL2(N695), .Z(N696) );
  GTECH_BUF B_29 ( .A(N694), .Z(N37) );
  SELECT_OP C24960 ( .DATA1(wrdata_d1[52]), .DATA2(N529), .CONTROL1(N34), 
        .CONTROL2(N686), .Z(N697) );
  SELECT_OP C24961 ( .DATA1(wrdata_d1[53]), .DATA2(N528), .CONTROL1(N35), 
        .CONTROL2(N689), .Z(N698) );
  SELECT_OP C24962 ( .DATA1(wrdata_d1[54]), .DATA2(N527), .CONTROL1(N36), 
        .CONTROL2(N692), .Z(N699) );
  SELECT_OP C24963 ( .DATA1(wrdata_d1[55]), .DATA2(N526), .CONTROL1(N37), 
        .CONTROL2(N695), .Z(N700) );
  SELECT_OP C24964 ( .DATA1(wrdata_d1[56]), .DATA2(N525), .CONTROL1(N38), 
        .CONTROL2(N702), .Z(N703) );
  GTECH_BUF B_30 ( .A(N701), .Z(N38) );
  SELECT_OP C24965 ( .DATA1(wrdata_d1[57]), .DATA2(N524), .CONTROL1(N39), 
        .CONTROL2(N705), .Z(N706) );
  GTECH_BUF B_31 ( .A(N704), .Z(N39) );
  SELECT_OP C24966 ( .DATA1(wrdata_d1[58]), .DATA2(N523), .CONTROL1(N40), 
        .CONTROL2(N708), .Z(N709) );
  GTECH_BUF B_32 ( .A(N707), .Z(N40) );
  SELECT_OP C24967 ( .DATA1(wrdata_d1[59]), .DATA2(N522), .CONTROL1(N41), 
        .CONTROL2(N711), .Z(N712) );
  GTECH_BUF B_33 ( .A(N710), .Z(N41) );
  SELECT_OP C24968 ( .DATA1(wrdata_d1[60]), .DATA2(N521), .CONTROL1(N38), 
        .CONTROL2(N702), .Z(N713) );
  SELECT_OP C24969 ( .DATA1(wrdata_d1[61]), .DATA2(N520), .CONTROL1(N39), 
        .CONTROL2(N705), .Z(N714) );
  SELECT_OP C24970 ( .DATA1(wrdata_d1[62]), .DATA2(N519), .CONTROL1(N40), 
        .CONTROL2(N708), .Z(N715) );
  SELECT_OP C24971 ( .DATA1(wrdata_d1[63]), .DATA2(N518), .CONTROL1(N41), 
        .CONTROL2(N711), .Z(N716) );
  SELECT_OP C24972 ( .DATA1(wrdata_d1[64]), .DATA2(N517), .CONTROL1(N42), 
        .CONTROL2(N718), .Z(N719) );
  GTECH_BUF B_34 ( .A(N717), .Z(N42) );
  SELECT_OP C24973 ( .DATA1(wrdata_d1[65]), .DATA2(N516), .CONTROL1(N43), 
        .CONTROL2(N721), .Z(N722) );
  GTECH_BUF B_35 ( .A(N720), .Z(N43) );
  SELECT_OP C24974 ( .DATA1(wrdata_d1[66]), .DATA2(N515), .CONTROL1(N44), 
        .CONTROL2(N724), .Z(N725) );
  GTECH_BUF B_36 ( .A(N723), .Z(N44) );
  SELECT_OP C24975 ( .DATA1(wrdata_d1[67]), .DATA2(N514), .CONTROL1(N45), 
        .CONTROL2(N727), .Z(N728) );
  GTECH_BUF B_37 ( .A(N726), .Z(N45) );
  SELECT_OP C24976 ( .DATA1(wrdata_d1[68]), .DATA2(N513), .CONTROL1(N42), 
        .CONTROL2(N718), .Z(N729) );
  SELECT_OP C24977 ( .DATA1(wrdata_d1[69]), .DATA2(N512), .CONTROL1(N43), 
        .CONTROL2(N721), .Z(N730) );
  SELECT_OP C24978 ( .DATA1(wrdata_d1[70]), .DATA2(N511), .CONTROL1(N44), 
        .CONTROL2(N724), .Z(N731) );
  SELECT_OP C24979 ( .DATA1(wrdata_d1[71]), .DATA2(N510), .CONTROL1(N45), 
        .CONTROL2(N727), .Z(N732) );
  SELECT_OP C24980 ( .DATA1(wrdata_d1[72]), .DATA2(N509), .CONTROL1(N46), 
        .CONTROL2(N734), .Z(N735) );
  GTECH_BUF B_38 ( .A(N733), .Z(N46) );
  SELECT_OP C24981 ( .DATA1(wrdata_d1[73]), .DATA2(N508), .CONTROL1(N47), 
        .CONTROL2(N737), .Z(N738) );
  GTECH_BUF B_39 ( .A(N736), .Z(N47) );
  SELECT_OP C24982 ( .DATA1(wrdata_d1[74]), .DATA2(N507), .CONTROL1(N48), 
        .CONTROL2(N740), .Z(N741) );
  GTECH_BUF B_40 ( .A(N739), .Z(N48) );
  SELECT_OP C24983 ( .DATA1(wrdata_d1[75]), .DATA2(N506), .CONTROL1(N49), 
        .CONTROL2(N743), .Z(N744) );
  GTECH_BUF B_41 ( .A(N742), .Z(N49) );
  SELECT_OP C24984 ( .DATA1(wrdata_d1[76]), .DATA2(N505), .CONTROL1(N46), 
        .CONTROL2(N734), .Z(N745) );
  SELECT_OP C24985 ( .DATA1(wrdata_d1[77]), .DATA2(N504), .CONTROL1(N47), 
        .CONTROL2(N737), .Z(N746) );
  SELECT_OP C24986 ( .DATA1(wrdata_d1[78]), .DATA2(N503), .CONTROL1(N48), 
        .CONTROL2(N740), .Z(N747) );
  SELECT_OP C24987 ( .DATA1(wrdata_d1[79]), .DATA2(N502), .CONTROL1(N49), 
        .CONTROL2(N743), .Z(N748) );
  SELECT_OP C24988 ( .DATA1(wrdata_d1[80]), .DATA2(N501), .CONTROL1(N50), 
        .CONTROL2(N750), .Z(N751) );
  GTECH_BUF B_42 ( .A(N749), .Z(N50) );
  SELECT_OP C24989 ( .DATA1(wrdata_d1[81]), .DATA2(N500), .CONTROL1(N51), 
        .CONTROL2(N753), .Z(N754) );
  GTECH_BUF B_43 ( .A(N752), .Z(N51) );
  SELECT_OP C24990 ( .DATA1(wrdata_d1[82]), .DATA2(N499), .CONTROL1(N52), 
        .CONTROL2(N756), .Z(N757) );
  GTECH_BUF B_44 ( .A(N755), .Z(N52) );
  SELECT_OP C24991 ( .DATA1(wrdata_d1[83]), .DATA2(N498), .CONTROL1(N53), 
        .CONTROL2(N759), .Z(N760) );
  GTECH_BUF B_45 ( .A(N758), .Z(N53) );
  SELECT_OP C24992 ( .DATA1(wrdata_d1[84]), .DATA2(N497), .CONTROL1(N50), 
        .CONTROL2(N750), .Z(N761) );
  SELECT_OP C24993 ( .DATA1(wrdata_d1[85]), .DATA2(N496), .CONTROL1(N51), 
        .CONTROL2(N753), .Z(N762) );
  SELECT_OP C24994 ( .DATA1(wrdata_d1[86]), .DATA2(N495), .CONTROL1(N52), 
        .CONTROL2(N756), .Z(N763) );
  SELECT_OP C24995 ( .DATA1(wrdata_d1[87]), .DATA2(N494), .CONTROL1(N53), 
        .CONTROL2(N759), .Z(N764) );
  SELECT_OP C24996 ( .DATA1(wrdata_d1[88]), .DATA2(N493), .CONTROL1(N54), 
        .CONTROL2(N766), .Z(N767) );
  GTECH_BUF B_46 ( .A(N765), .Z(N54) );
  SELECT_OP C24997 ( .DATA1(wrdata_d1[89]), .DATA2(N492), .CONTROL1(N55), 
        .CONTROL2(N769), .Z(N770) );
  GTECH_BUF B_47 ( .A(N768), .Z(N55) );
  SELECT_OP C24998 ( .DATA1(wrdata_d1[90]), .DATA2(N491), .CONTROL1(N56), 
        .CONTROL2(N772), .Z(N773) );
  GTECH_BUF B_48 ( .A(N771), .Z(N56) );
  SELECT_OP C24999 ( .DATA1(wrdata_d1[91]), .DATA2(N490), .CONTROL1(N57), 
        .CONTROL2(N775), .Z(N776) );
  GTECH_BUF B_49 ( .A(N774), .Z(N57) );
  SELECT_OP C25000 ( .DATA1(wrdata_d1[92]), .DATA2(N489), .CONTROL1(N54), 
        .CONTROL2(N766), .Z(N777) );
  SELECT_OP C25001 ( .DATA1(wrdata_d1[93]), .DATA2(N488), .CONTROL1(N55), 
        .CONTROL2(N769), .Z(N778) );
  SELECT_OP C25002 ( .DATA1(wrdata_d1[94]), .DATA2(N487), .CONTROL1(N56), 
        .CONTROL2(N772), .Z(N779) );
  SELECT_OP C25003 ( .DATA1(wrdata_d1[95]), .DATA2(N486), .CONTROL1(N57), 
        .CONTROL2(N775), .Z(N780) );
  SELECT_OP C25004 ( .DATA1(wrdata_d1[96]), .DATA2(N485), .CONTROL1(N58), 
        .CONTROL2(N782), .Z(N783) );
  GTECH_BUF B_50 ( .A(N781), .Z(N58) );
  SELECT_OP C25005 ( .DATA1(wrdata_d1[97]), .DATA2(N484), .CONTROL1(N59), 
        .CONTROL2(N785), .Z(N786) );
  GTECH_BUF B_51 ( .A(N784), .Z(N59) );
  SELECT_OP C25006 ( .DATA1(wrdata_d1[98]), .DATA2(N483), .CONTROL1(N60), 
        .CONTROL2(N788), .Z(N789) );
  GTECH_BUF B_52 ( .A(N787), .Z(N60) );
  SELECT_OP C25007 ( .DATA1(wrdata_d1[99]), .DATA2(N482), .CONTROL1(N61), 
        .CONTROL2(N791), .Z(N792) );
  GTECH_BUF B_53 ( .A(N790), .Z(N61) );
  SELECT_OP C25008 ( .DATA1(wrdata_d1[100]), .DATA2(N481), .CONTROL1(N58), 
        .CONTROL2(N782), .Z(N793) );
  SELECT_OP C25009 ( .DATA1(wrdata_d1[101]), .DATA2(N480), .CONTROL1(N59), 
        .CONTROL2(N785), .Z(N794) );
  SELECT_OP C25010 ( .DATA1(wrdata_d1[102]), .DATA2(N479), .CONTROL1(N60), 
        .CONTROL2(N788), .Z(N795) );
  SELECT_OP C25011 ( .DATA1(wrdata_d1[103]), .DATA2(N478), .CONTROL1(N61), 
        .CONTROL2(N791), .Z(N796) );
  SELECT_OP C25012 ( .DATA1(wrdata_d1[104]), .DATA2(N477), .CONTROL1(N62), 
        .CONTROL2(N798), .Z(N799) );
  GTECH_BUF B_54 ( .A(N797), .Z(N62) );
  SELECT_OP C25013 ( .DATA1(wrdata_d1[105]), .DATA2(N476), .CONTROL1(N63), 
        .CONTROL2(N801), .Z(N802) );
  GTECH_BUF B_55 ( .A(N800), .Z(N63) );
  SELECT_OP C25014 ( .DATA1(wrdata_d1[106]), .DATA2(N475), .CONTROL1(N64), 
        .CONTROL2(N804), .Z(N805) );
  GTECH_BUF B_56 ( .A(N803), .Z(N64) );
  SELECT_OP C25015 ( .DATA1(wrdata_d1[107]), .DATA2(N474), .CONTROL1(N65), 
        .CONTROL2(N807), .Z(N808) );
  GTECH_BUF B_57 ( .A(N806), .Z(N65) );
  SELECT_OP C25016 ( .DATA1(wrdata_d1[108]), .DATA2(N473), .CONTROL1(N62), 
        .CONTROL2(N798), .Z(N809) );
  SELECT_OP C25017 ( .DATA1(wrdata_d1[109]), .DATA2(N472), .CONTROL1(N63), 
        .CONTROL2(N801), .Z(N810) );
  SELECT_OP C25018 ( .DATA1(wrdata_d1[110]), .DATA2(N471), .CONTROL1(N64), 
        .CONTROL2(N804), .Z(N811) );
  SELECT_OP C25019 ( .DATA1(wrdata_d1[111]), .DATA2(N470), .CONTROL1(N65), 
        .CONTROL2(N807), .Z(N812) );
  SELECT_OP C25020 ( .DATA1(wrdata_d1[112]), .DATA2(N469), .CONTROL1(N66), 
        .CONTROL2(N814), .Z(N815) );
  GTECH_BUF B_58 ( .A(N813), .Z(N66) );
  SELECT_OP C25021 ( .DATA1(wrdata_d1[113]), .DATA2(N468), .CONTROL1(N67), 
        .CONTROL2(N817), .Z(N818) );
  GTECH_BUF B_59 ( .A(N816), .Z(N67) );
  SELECT_OP C25022 ( .DATA1(wrdata_d1[114]), .DATA2(N467), .CONTROL1(N68), 
        .CONTROL2(N820), .Z(N821) );
  GTECH_BUF B_60 ( .A(N819), .Z(N68) );
  SELECT_OP C25023 ( .DATA1(wrdata_d1[115]), .DATA2(N466), .CONTROL1(N69), 
        .CONTROL2(N823), .Z(N824) );
  GTECH_BUF B_61 ( .A(N822), .Z(N69) );
  SELECT_OP C25024 ( .DATA1(wrdata_d1[116]), .DATA2(N465), .CONTROL1(N66), 
        .CONTROL2(N814), .Z(N825) );
  SELECT_OP C25025 ( .DATA1(wrdata_d1[117]), .DATA2(N464), .CONTROL1(N67), 
        .CONTROL2(N817), .Z(N826) );
  SELECT_OP C25026 ( .DATA1(wrdata_d1[118]), .DATA2(N463), .CONTROL1(N68), 
        .CONTROL2(N820), .Z(N827) );
  SELECT_OP C25027 ( .DATA1(wrdata_d1[119]), .DATA2(N462), .CONTROL1(N69), 
        .CONTROL2(N823), .Z(N828) );
  SELECT_OP C25028 ( .DATA1(wrdata_d1[120]), .DATA2(N461), .CONTROL1(N70), 
        .CONTROL2(N830), .Z(N831) );
  GTECH_BUF B_62 ( .A(N829), .Z(N70) );
  SELECT_OP C25029 ( .DATA1(wrdata_d1[121]), .DATA2(N460), .CONTROL1(N71), 
        .CONTROL2(N833), .Z(N834) );
  GTECH_BUF B_63 ( .A(N832), .Z(N71) );
  SELECT_OP C25030 ( .DATA1(wrdata_d1[122]), .DATA2(N459), .CONTROL1(N72), 
        .CONTROL2(N836), .Z(N837) );
  GTECH_BUF B_64 ( .A(N835), .Z(N72) );
  SELECT_OP C25031 ( .DATA1(wrdata_d1[123]), .DATA2(N458), .CONTROL1(N73), 
        .CONTROL2(N839), .Z(N840) );
  GTECH_BUF B_65 ( .A(N838), .Z(N73) );
  SELECT_OP C25032 ( .DATA1(wrdata_d1[124]), .DATA2(N457), .CONTROL1(N70), 
        .CONTROL2(N830), .Z(N841) );
  SELECT_OP C25033 ( .DATA1(wrdata_d1[125]), .DATA2(N456), .CONTROL1(N71), 
        .CONTROL2(N833), .Z(N842) );
  SELECT_OP C25034 ( .DATA1(wrdata_d1[126]), .DATA2(N455), .CONTROL1(N72), 
        .CONTROL2(N836), .Z(N843) );
  SELECT_OP C25035 ( .DATA1(wrdata_d1[127]), .DATA2(N454), .CONTROL1(N73), 
        .CONTROL2(N839), .Z(N844) );
  SELECT_OP C25036 ( .DATA1(wrdata_d1[128]), .DATA2(N453), .CONTROL1(N74), 
        .CONTROL2(N846), .Z(N847) );
  GTECH_BUF B_66 ( .A(N845), .Z(N74) );
  SELECT_OP C25037 ( .DATA1(wrdata_d1[129]), .DATA2(N452), .CONTROL1(N75), 
        .CONTROL2(N849), .Z(N850) );
  GTECH_BUF B_67 ( .A(N848), .Z(N75) );
  SELECT_OP C25038 ( .DATA1(wrdata_d1[130]), .DATA2(N451), .CONTROL1(N76), 
        .CONTROL2(N852), .Z(N853) );
  GTECH_BUF B_68 ( .A(N851), .Z(N76) );
  SELECT_OP C25039 ( .DATA1(wrdata_d1[131]), .DATA2(N450), .CONTROL1(N77), 
        .CONTROL2(N855), .Z(N856) );
  GTECH_BUF B_69 ( .A(N854), .Z(N77) );
  SELECT_OP C25040 ( .DATA1(wrdata_d1[132]), .DATA2(N449), .CONTROL1(N74), 
        .CONTROL2(N846), .Z(N857) );
  SELECT_OP C25041 ( .DATA1(wrdata_d1[133]), .DATA2(N448), .CONTROL1(N75), 
        .CONTROL2(N849), .Z(N858) );
  SELECT_OP C25042 ( .DATA1(wrdata_d1[134]), .DATA2(N447), .CONTROL1(N76), 
        .CONTROL2(N852), .Z(N859) );
  SELECT_OP C25043 ( .DATA1(wrdata_d1[135]), .DATA2(N446), .CONTROL1(N77), 
        .CONTROL2(N855), .Z(N860) );
  SELECT_OP C25044 ( .DATA1(wrdata_d1[136]), .DATA2(N445), .CONTROL1(N78), 
        .CONTROL2(N862), .Z(N863) );
  GTECH_BUF B_70 ( .A(N861), .Z(N78) );
  SELECT_OP C25045 ( .DATA1(wrdata_d1[137]), .DATA2(N444), .CONTROL1(N79), 
        .CONTROL2(N865), .Z(N866) );
  GTECH_BUF B_71 ( .A(N864), .Z(N79) );
  SELECT_OP C25046 ( .DATA1(wrdata_d1[138]), .DATA2(N443), .CONTROL1(N80), 
        .CONTROL2(N868), .Z(N869) );
  GTECH_BUF B_72 ( .A(N867), .Z(N80) );
  SELECT_OP C25047 ( .DATA1(wrdata_d1[139]), .DATA2(N442), .CONTROL1(N81), 
        .CONTROL2(N871), .Z(N872) );
  GTECH_BUF B_73 ( .A(N870), .Z(N81) );
  SELECT_OP C25048 ( .DATA1(wrdata_d1[140]), .DATA2(N441), .CONTROL1(N78), 
        .CONTROL2(N862), .Z(N873) );
  SELECT_OP C25049 ( .DATA1(wrdata_d1[141]), .DATA2(N440), .CONTROL1(N79), 
        .CONTROL2(N865), .Z(N874) );
  SELECT_OP C25050 ( .DATA1(wrdata_d1[142]), .DATA2(N439), .CONTROL1(N80), 
        .CONTROL2(N868), .Z(N875) );
  SELECT_OP C25051 ( .DATA1(wrdata_d1[143]), .DATA2(N438), .CONTROL1(N81), 
        .CONTROL2(N871), .Z(N876) );
  SELECT_OP C25052 ( .DATA1(wrdata_d1[144]), .DATA2(N437), .CONTROL1(N82), 
        .CONTROL2(N878), .Z(N879) );
  GTECH_BUF B_74 ( .A(N877), .Z(N82) );
  SELECT_OP C25053 ( .DATA1(wrdata_d1[145]), .DATA2(N436), .CONTROL1(N83), 
        .CONTROL2(N881), .Z(N882) );
  GTECH_BUF B_75 ( .A(N880), .Z(N83) );
  SELECT_OP C25054 ( .DATA1(wrdata_d1[146]), .DATA2(N435), .CONTROL1(N84), 
        .CONTROL2(N884), .Z(N885) );
  GTECH_BUF B_76 ( .A(N883), .Z(N84) );
  SELECT_OP C25055 ( .DATA1(wrdata_d1[147]), .DATA2(N434), .CONTROL1(N85), 
        .CONTROL2(N887), .Z(N888) );
  GTECH_BUF B_77 ( .A(N886), .Z(N85) );
  SELECT_OP C25056 ( .DATA1(wrdata_d1[148]), .DATA2(N433), .CONTROL1(N82), 
        .CONTROL2(N878), .Z(N889) );
  SELECT_OP C25057 ( .DATA1(wrdata_d1[149]), .DATA2(N432), .CONTROL1(N83), 
        .CONTROL2(N881), .Z(N890) );
  SELECT_OP C25058 ( .DATA1(wrdata_d1[150]), .DATA2(N431), .CONTROL1(N84), 
        .CONTROL2(N884), .Z(N891) );
  SELECT_OP C25059 ( .DATA1(wrdata_d1[151]), .DATA2(N430), .CONTROL1(N85), 
        .CONTROL2(N887), .Z(N892) );
  SELECT_OP C25060 ( .DATA1(wrdata_d1[152]), .DATA2(N429), .CONTROL1(N86), 
        .CONTROL2(N894), .Z(N895) );
  GTECH_BUF B_78 ( .A(N893), .Z(N86) );
  SELECT_OP C25061 ( .DATA1(wrdata_d1[153]), .DATA2(N428), .CONTROL1(N87), 
        .CONTROL2(N897), .Z(N898) );
  GTECH_BUF B_79 ( .A(N896), .Z(N87) );
  SELECT_OP C25062 ( .DATA1(wrdata_d1[154]), .DATA2(N427), .CONTROL1(N88), 
        .CONTROL2(N900), .Z(N901) );
  GTECH_BUF B_80 ( .A(N899), .Z(N88) );
  SELECT_OP C25063 ( .DATA1(wrdata_d1[155]), .DATA2(N426), .CONTROL1(N89), 
        .CONTROL2(N903), .Z(N904) );
  GTECH_BUF B_81 ( .A(N902), .Z(N89) );
  SELECT_OP C25064 ( .DATA1(wrdata_d1[156]), .DATA2(N425), .CONTROL1(N86), 
        .CONTROL2(N894), .Z(N905) );
  SELECT_OP C25065 ( .DATA1(wrdata_d1[157]), .DATA2(N424), .CONTROL1(N87), 
        .CONTROL2(N897), .Z(N906) );
  SELECT_OP C25066 ( .DATA1(wrdata_d1[158]), .DATA2(N423), .CONTROL1(N88), 
        .CONTROL2(N900), .Z(N907) );
  SELECT_OP C25067 ( .DATA1(wrdata_d1[159]), .DATA2(N422), .CONTROL1(N89), 
        .CONTROL2(N903), .Z(N908) );
  SELECT_OP C25068 ( .DATA1({N924, N924, N923, N923, N922, N922, N921, N921, 
        N920, N920, N919, N919, N918, N918, N917, N917, N916, N916, N915, N915, 
        N914, N914, N913, N913, N912, N912, N911, N911, N910, N910, N909, N909}), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N90), 
        .CONTROL2(N588), .Z({N956, N955, N954, N953, N952, N951, N950, N949, 
        N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, 
        N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925}) );
  GTECH_BUF B_82 ( .A(N587), .Z(N90) );
  SELECT_OP C25069 ( .DATA1({N956, N955, N954, N953, N952, N951, N950, N949, 
        N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, 
        N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925}), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CONTROL1(N8), 
        .CONTROL2(N9), .Z({N988, N987, N986, N985, N984, N983, N982, N981, 
        N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957}) );
  MUX_OP C25070 ( .D0({\inq_ary[0][0] , \inq_ary[0][1] , \inq_ary[0][2] , 
        \inq_ary[0][3] , \inq_ary[0][4] , \inq_ary[0][5] , \inq_ary[0][6] , 
        \inq_ary[0][7] , \inq_ary[0][8] , \inq_ary[0][9] , \inq_ary[0][10] , 
        \inq_ary[0][11] , \inq_ary[0][12] , \inq_ary[0][13] , \inq_ary[0][14] , 
        \inq_ary[0][15] , \inq_ary[0][16] , \inq_ary[0][17] , \inq_ary[0][18] , 
        \inq_ary[0][19] , \inq_ary[0][20] , \inq_ary[0][21] , \inq_ary[0][22] , 
        \inq_ary[0][23] , \inq_ary[0][24] , \inq_ary[0][25] , \inq_ary[0][26] , 
        \inq_ary[0][27] , \inq_ary[0][28] , \inq_ary[0][29] , \inq_ary[0][30] , 
        \inq_ary[0][31] , \inq_ary[0][32] , \inq_ary[0][33] , \inq_ary[0][34] , 
        \inq_ary[0][35] , \inq_ary[0][36] , \inq_ary[0][37] , \inq_ary[0][38] , 
        \inq_ary[0][39] , \inq_ary[0][40] , \inq_ary[0][41] , \inq_ary[0][42] , 
        \inq_ary[0][43] , \inq_ary[0][44] , \inq_ary[0][45] , \inq_ary[0][46] , 
        \inq_ary[0][47] , \inq_ary[0][48] , \inq_ary[0][49] , \inq_ary[0][50] , 
        \inq_ary[0][51] , \inq_ary[0][52] , \inq_ary[0][53] , \inq_ary[0][54] , 
        \inq_ary[0][55] , \inq_ary[0][56] , \inq_ary[0][57] , \inq_ary[0][58] , 
        \inq_ary[0][59] , \inq_ary[0][60] , \inq_ary[0][61] , \inq_ary[0][62] , 
        \inq_ary[0][63] , \inq_ary[0][64] , \inq_ary[0][65] , \inq_ary[0][66] , 
        \inq_ary[0][67] , \inq_ary[0][68] , \inq_ary[0][69] , \inq_ary[0][70] , 
        \inq_ary[0][71] , \inq_ary[0][72] , \inq_ary[0][73] , \inq_ary[0][74] , 
        \inq_ary[0][75] , \inq_ary[0][76] , \inq_ary[0][77] , \inq_ary[0][78] , 
        \inq_ary[0][79] , \inq_ary[0][80] , \inq_ary[0][81] , \inq_ary[0][82] , 
        \inq_ary[0][83] , \inq_ary[0][84] , \inq_ary[0][85] , \inq_ary[0][86] , 
        \inq_ary[0][87] , \inq_ary[0][88] , \inq_ary[0][89] , \inq_ary[0][90] , 
        \inq_ary[0][91] , \inq_ary[0][92] , \inq_ary[0][93] , \inq_ary[0][94] , 
        \inq_ary[0][95] , \inq_ary[0][96] , \inq_ary[0][97] , \inq_ary[0][98] , 
        \inq_ary[0][99] , \inq_ary[0][100] , \inq_ary[0][101] , 
        \inq_ary[0][102] , \inq_ary[0][103] , \inq_ary[0][104] , 
        \inq_ary[0][105] , \inq_ary[0][106] , \inq_ary[0][107] , 
        \inq_ary[0][108] , \inq_ary[0][109] , \inq_ary[0][110] , 
        \inq_ary[0][111] , \inq_ary[0][112] , \inq_ary[0][113] , 
        \inq_ary[0][114] , \inq_ary[0][115] , \inq_ary[0][116] , 
        \inq_ary[0][117] , \inq_ary[0][118] , \inq_ary[0][119] , 
        \inq_ary[0][120] , \inq_ary[0][121] , \inq_ary[0][122] , 
        \inq_ary[0][123] , \inq_ary[0][124] , \inq_ary[0][125] , 
        \inq_ary[0][126] , \inq_ary[0][127] , \inq_ary[0][128] , 
        \inq_ary[0][129] , \inq_ary[0][130] , \inq_ary[0][131] , 
        \inq_ary[0][132] , \inq_ary[0][133] , \inq_ary[0][134] , 
        \inq_ary[0][135] , \inq_ary[0][136] , \inq_ary[0][137] , 
        \inq_ary[0][138] , \inq_ary[0][139] , \inq_ary[0][140] , 
        \inq_ary[0][141] , \inq_ary[0][142] , \inq_ary[0][143] , 
        \inq_ary[0][144] , \inq_ary[0][145] , \inq_ary[0][146] , 
        \inq_ary[0][147] , \inq_ary[0][148] , \inq_ary[0][149] , 
        \inq_ary[0][150] , \inq_ary[0][151] , \inq_ary[0][152] , 
        \inq_ary[0][153] , \inq_ary[0][154] , \inq_ary[0][155] , 
        \inq_ary[0][156] , \inq_ary[0][157] , \inq_ary[0][158] , 
        \inq_ary[0][159] }), .D1({\inq_ary[1][0] , \inq_ary[1][1] , 
        \inq_ary[1][2] , \inq_ary[1][3] , \inq_ary[1][4] , \inq_ary[1][5] , 
        \inq_ary[1][6] , \inq_ary[1][7] , \inq_ary[1][8] , \inq_ary[1][9] , 
        \inq_ary[1][10] , \inq_ary[1][11] , \inq_ary[1][12] , \inq_ary[1][13] , 
        \inq_ary[1][14] , \inq_ary[1][15] , \inq_ary[1][16] , \inq_ary[1][17] , 
        \inq_ary[1][18] , \inq_ary[1][19] , \inq_ary[1][20] , \inq_ary[1][21] , 
        \inq_ary[1][22] , \inq_ary[1][23] , \inq_ary[1][24] , \inq_ary[1][25] , 
        \inq_ary[1][26] , \inq_ary[1][27] , \inq_ary[1][28] , \inq_ary[1][29] , 
        \inq_ary[1][30] , \inq_ary[1][31] , \inq_ary[1][32] , \inq_ary[1][33] , 
        \inq_ary[1][34] , \inq_ary[1][35] , \inq_ary[1][36] , \inq_ary[1][37] , 
        \inq_ary[1][38] , \inq_ary[1][39] , \inq_ary[1][40] , \inq_ary[1][41] , 
        \inq_ary[1][42] , \inq_ary[1][43] , \inq_ary[1][44] , \inq_ary[1][45] , 
        \inq_ary[1][46] , \inq_ary[1][47] , \inq_ary[1][48] , \inq_ary[1][49] , 
        \inq_ary[1][50] , \inq_ary[1][51] , \inq_ary[1][52] , \inq_ary[1][53] , 
        \inq_ary[1][54] , \inq_ary[1][55] , \inq_ary[1][56] , \inq_ary[1][57] , 
        \inq_ary[1][58] , \inq_ary[1][59] , \inq_ary[1][60] , \inq_ary[1][61] , 
        \inq_ary[1][62] , \inq_ary[1][63] , \inq_ary[1][64] , \inq_ary[1][65] , 
        \inq_ary[1][66] , \inq_ary[1][67] , \inq_ary[1][68] , \inq_ary[1][69] , 
        \inq_ary[1][70] , \inq_ary[1][71] , \inq_ary[1][72] , \inq_ary[1][73] , 
        \inq_ary[1][74] , \inq_ary[1][75] , \inq_ary[1][76] , \inq_ary[1][77] , 
        \inq_ary[1][78] , \inq_ary[1][79] , \inq_ary[1][80] , \inq_ary[1][81] , 
        \inq_ary[1][82] , \inq_ary[1][83] , \inq_ary[1][84] , \inq_ary[1][85] , 
        \inq_ary[1][86] , \inq_ary[1][87] , \inq_ary[1][88] , \inq_ary[1][89] , 
        \inq_ary[1][90] , \inq_ary[1][91] , \inq_ary[1][92] , \inq_ary[1][93] , 
        \inq_ary[1][94] , \inq_ary[1][95] , \inq_ary[1][96] , \inq_ary[1][97] , 
        \inq_ary[1][98] , \inq_ary[1][99] , \inq_ary[1][100] , 
        \inq_ary[1][101] , \inq_ary[1][102] , \inq_ary[1][103] , 
        \inq_ary[1][104] , \inq_ary[1][105] , \inq_ary[1][106] , 
        \inq_ary[1][107] , \inq_ary[1][108] , \inq_ary[1][109] , 
        \inq_ary[1][110] , \inq_ary[1][111] , \inq_ary[1][112] , 
        \inq_ary[1][113] , \inq_ary[1][114] , \inq_ary[1][115] , 
        \inq_ary[1][116] , \inq_ary[1][117] , \inq_ary[1][118] , 
        \inq_ary[1][119] , \inq_ary[1][120] , \inq_ary[1][121] , 
        \inq_ary[1][122] , \inq_ary[1][123] , \inq_ary[1][124] , 
        \inq_ary[1][125] , \inq_ary[1][126] , \inq_ary[1][127] , 
        \inq_ary[1][128] , \inq_ary[1][129] , \inq_ary[1][130] , 
        \inq_ary[1][131] , \inq_ary[1][132] , \inq_ary[1][133] , 
        \inq_ary[1][134] , \inq_ary[1][135] , \inq_ary[1][136] , 
        \inq_ary[1][137] , \inq_ary[1][138] , \inq_ary[1][139] , 
        \inq_ary[1][140] , \inq_ary[1][141] , \inq_ary[1][142] , 
        \inq_ary[1][143] , \inq_ary[1][144] , \inq_ary[1][145] , 
        \inq_ary[1][146] , \inq_ary[1][147] , \inq_ary[1][148] , 
        \inq_ary[1][149] , \inq_ary[1][150] , \inq_ary[1][151] , 
        \inq_ary[1][152] , \inq_ary[1][153] , \inq_ary[1][154] , 
        \inq_ary[1][155] , \inq_ary[1][156] , \inq_ary[1][157] , 
        \inq_ary[1][158] , \inq_ary[1][159] }), .D2({\inq_ary[2][0] , 
        \inq_ary[2][1] , \inq_ary[2][2] , \inq_ary[2][3] , \inq_ary[2][4] , 
        \inq_ary[2][5] , \inq_ary[2][6] , \inq_ary[2][7] , \inq_ary[2][8] , 
        \inq_ary[2][9] , \inq_ary[2][10] , \inq_ary[2][11] , \inq_ary[2][12] , 
        \inq_ary[2][13] , \inq_ary[2][14] , \inq_ary[2][15] , \inq_ary[2][16] , 
        \inq_ary[2][17] , \inq_ary[2][18] , \inq_ary[2][19] , \inq_ary[2][20] , 
        \inq_ary[2][21] , \inq_ary[2][22] , \inq_ary[2][23] , \inq_ary[2][24] , 
        \inq_ary[2][25] , \inq_ary[2][26] , \inq_ary[2][27] , \inq_ary[2][28] , 
        \inq_ary[2][29] , \inq_ary[2][30] , \inq_ary[2][31] , \inq_ary[2][32] , 
        \inq_ary[2][33] , \inq_ary[2][34] , \inq_ary[2][35] , \inq_ary[2][36] , 
        \inq_ary[2][37] , \inq_ary[2][38] , \inq_ary[2][39] , \inq_ary[2][40] , 
        \inq_ary[2][41] , \inq_ary[2][42] , \inq_ary[2][43] , \inq_ary[2][44] , 
        \inq_ary[2][45] , \inq_ary[2][46] , \inq_ary[2][47] , \inq_ary[2][48] , 
        \inq_ary[2][49] , \inq_ary[2][50] , \inq_ary[2][51] , \inq_ary[2][52] , 
        \inq_ary[2][53] , \inq_ary[2][54] , \inq_ary[2][55] , \inq_ary[2][56] , 
        \inq_ary[2][57] , \inq_ary[2][58] , \inq_ary[2][59] , \inq_ary[2][60] , 
        \inq_ary[2][61] , \inq_ary[2][62] , \inq_ary[2][63] , \inq_ary[2][64] , 
        \inq_ary[2][65] , \inq_ary[2][66] , \inq_ary[2][67] , \inq_ary[2][68] , 
        \inq_ary[2][69] , \inq_ary[2][70] , \inq_ary[2][71] , \inq_ary[2][72] , 
        \inq_ary[2][73] , \inq_ary[2][74] , \inq_ary[2][75] , \inq_ary[2][76] , 
        \inq_ary[2][77] , \inq_ary[2][78] , \inq_ary[2][79] , \inq_ary[2][80] , 
        \inq_ary[2][81] , \inq_ary[2][82] , \inq_ary[2][83] , \inq_ary[2][84] , 
        \inq_ary[2][85] , \inq_ary[2][86] , \inq_ary[2][87] , \inq_ary[2][88] , 
        \inq_ary[2][89] , \inq_ary[2][90] , \inq_ary[2][91] , \inq_ary[2][92] , 
        \inq_ary[2][93] , \inq_ary[2][94] , \inq_ary[2][95] , \inq_ary[2][96] , 
        \inq_ary[2][97] , \inq_ary[2][98] , \inq_ary[2][99] , 
        \inq_ary[2][100] , \inq_ary[2][101] , \inq_ary[2][102] , 
        \inq_ary[2][103] , \inq_ary[2][104] , \inq_ary[2][105] , 
        \inq_ary[2][106] , \inq_ary[2][107] , \inq_ary[2][108] , 
        \inq_ary[2][109] , \inq_ary[2][110] , \inq_ary[2][111] , 
        \inq_ary[2][112] , \inq_ary[2][113] , \inq_ary[2][114] , 
        \inq_ary[2][115] , \inq_ary[2][116] , \inq_ary[2][117] , 
        \inq_ary[2][118] , \inq_ary[2][119] , \inq_ary[2][120] , 
        \inq_ary[2][121] , \inq_ary[2][122] , \inq_ary[2][123] , 
        \inq_ary[2][124] , \inq_ary[2][125] , \inq_ary[2][126] , 
        \inq_ary[2][127] , \inq_ary[2][128] , \inq_ary[2][129] , 
        \inq_ary[2][130] , \inq_ary[2][131] , \inq_ary[2][132] , 
        \inq_ary[2][133] , \inq_ary[2][134] , \inq_ary[2][135] , 
        \inq_ary[2][136] , \inq_ary[2][137] , \inq_ary[2][138] , 
        \inq_ary[2][139] , \inq_ary[2][140] , \inq_ary[2][141] , 
        \inq_ary[2][142] , \inq_ary[2][143] , \inq_ary[2][144] , 
        \inq_ary[2][145] , \inq_ary[2][146] , \inq_ary[2][147] , 
        \inq_ary[2][148] , \inq_ary[2][149] , \inq_ary[2][150] , 
        \inq_ary[2][151] , \inq_ary[2][152] , \inq_ary[2][153] , 
        \inq_ary[2][154] , \inq_ary[2][155] , \inq_ary[2][156] , 
        \inq_ary[2][157] , \inq_ary[2][158] , \inq_ary[2][159] }), .D3({
        \inq_ary[3][0] , \inq_ary[3][1] , \inq_ary[3][2] , \inq_ary[3][3] , 
        \inq_ary[3][4] , \inq_ary[3][5] , \inq_ary[3][6] , \inq_ary[3][7] , 
        \inq_ary[3][8] , \inq_ary[3][9] , \inq_ary[3][10] , \inq_ary[3][11] , 
        \inq_ary[3][12] , \inq_ary[3][13] , \inq_ary[3][14] , \inq_ary[3][15] , 
        \inq_ary[3][16] , \inq_ary[3][17] , \inq_ary[3][18] , \inq_ary[3][19] , 
        \inq_ary[3][20] , \inq_ary[3][21] , \inq_ary[3][22] , \inq_ary[3][23] , 
        \inq_ary[3][24] , \inq_ary[3][25] , \inq_ary[3][26] , \inq_ary[3][27] , 
        \inq_ary[3][28] , \inq_ary[3][29] , \inq_ary[3][30] , \inq_ary[3][31] , 
        \inq_ary[3][32] , \inq_ary[3][33] , \inq_ary[3][34] , \inq_ary[3][35] , 
        \inq_ary[3][36] , \inq_ary[3][37] , \inq_ary[3][38] , \inq_ary[3][39] , 
        \inq_ary[3][40] , \inq_ary[3][41] , \inq_ary[3][42] , \inq_ary[3][43] , 
        \inq_ary[3][44] , \inq_ary[3][45] , \inq_ary[3][46] , \inq_ary[3][47] , 
        \inq_ary[3][48] , \inq_ary[3][49] , \inq_ary[3][50] , \inq_ary[3][51] , 
        \inq_ary[3][52] , \inq_ary[3][53] , \inq_ary[3][54] , \inq_ary[3][55] , 
        \inq_ary[3][56] , \inq_ary[3][57] , \inq_ary[3][58] , \inq_ary[3][59] , 
        \inq_ary[3][60] , \inq_ary[3][61] , \inq_ary[3][62] , \inq_ary[3][63] , 
        \inq_ary[3][64] , \inq_ary[3][65] , \inq_ary[3][66] , \inq_ary[3][67] , 
        \inq_ary[3][68] , \inq_ary[3][69] , \inq_ary[3][70] , \inq_ary[3][71] , 
        \inq_ary[3][72] , \inq_ary[3][73] , \inq_ary[3][74] , \inq_ary[3][75] , 
        \inq_ary[3][76] , \inq_ary[3][77] , \inq_ary[3][78] , \inq_ary[3][79] , 
        \inq_ary[3][80] , \inq_ary[3][81] , \inq_ary[3][82] , \inq_ary[3][83] , 
        \inq_ary[3][84] , \inq_ary[3][85] , \inq_ary[3][86] , \inq_ary[3][87] , 
        \inq_ary[3][88] , \inq_ary[3][89] , \inq_ary[3][90] , \inq_ary[3][91] , 
        \inq_ary[3][92] , \inq_ary[3][93] , \inq_ary[3][94] , \inq_ary[3][95] , 
        \inq_ary[3][96] , \inq_ary[3][97] , \inq_ary[3][98] , \inq_ary[3][99] , 
        \inq_ary[3][100] , \inq_ary[3][101] , \inq_ary[3][102] , 
        \inq_ary[3][103] , \inq_ary[3][104] , \inq_ary[3][105] , 
        \inq_ary[3][106] , \inq_ary[3][107] , \inq_ary[3][108] , 
        \inq_ary[3][109] , \inq_ary[3][110] , \inq_ary[3][111] , 
        \inq_ary[3][112] , \inq_ary[3][113] , \inq_ary[3][114] , 
        \inq_ary[3][115] , \inq_ary[3][116] , \inq_ary[3][117] , 
        \inq_ary[3][118] , \inq_ary[3][119] , \inq_ary[3][120] , 
        \inq_ary[3][121] , \inq_ary[3][122] , \inq_ary[3][123] , 
        \inq_ary[3][124] , \inq_ary[3][125] , \inq_ary[3][126] , 
        \inq_ary[3][127] , \inq_ary[3][128] , \inq_ary[3][129] , 
        \inq_ary[3][130] , \inq_ary[3][131] , \inq_ary[3][132] , 
        \inq_ary[3][133] , \inq_ary[3][134] , \inq_ary[3][135] , 
        \inq_ary[3][136] , \inq_ary[3][137] , \inq_ary[3][138] , 
        \inq_ary[3][139] , \inq_ary[3][140] , \inq_ary[3][141] , 
        \inq_ary[3][142] , \inq_ary[3][143] , \inq_ary[3][144] , 
        \inq_ary[3][145] , \inq_ary[3][146] , \inq_ary[3][147] , 
        \inq_ary[3][148] , \inq_ary[3][149] , \inq_ary[3][150] , 
        \inq_ary[3][151] , \inq_ary[3][152] , \inq_ary[3][153] , 
        \inq_ary[3][154] , \inq_ary[3][155] , \inq_ary[3][156] , 
        \inq_ary[3][157] , \inq_ary[3][158] , \inq_ary[3][159] }), .D4({
        \inq_ary[4][0] , \inq_ary[4][1] , \inq_ary[4][2] , \inq_ary[4][3] , 
        \inq_ary[4][4] , \inq_ary[4][5] , \inq_ary[4][6] , \inq_ary[4][7] , 
        \inq_ary[4][8] , \inq_ary[4][9] , \inq_ary[4][10] , \inq_ary[4][11] , 
        \inq_ary[4][12] , \inq_ary[4][13] , \inq_ary[4][14] , \inq_ary[4][15] , 
        \inq_ary[4][16] , \inq_ary[4][17] , \inq_ary[4][18] , \inq_ary[4][19] , 
        \inq_ary[4][20] , \inq_ary[4][21] , \inq_ary[4][22] , \inq_ary[4][23] , 
        \inq_ary[4][24] , \inq_ary[4][25] , \inq_ary[4][26] , \inq_ary[4][27] , 
        \inq_ary[4][28] , \inq_ary[4][29] , \inq_ary[4][30] , \inq_ary[4][31] , 
        \inq_ary[4][32] , \inq_ary[4][33] , \inq_ary[4][34] , \inq_ary[4][35] , 
        \inq_ary[4][36] , \inq_ary[4][37] , \inq_ary[4][38] , \inq_ary[4][39] , 
        \inq_ary[4][40] , \inq_ary[4][41] , \inq_ary[4][42] , \inq_ary[4][43] , 
        \inq_ary[4][44] , \inq_ary[4][45] , \inq_ary[4][46] , \inq_ary[4][47] , 
        \inq_ary[4][48] , \inq_ary[4][49] , \inq_ary[4][50] , \inq_ary[4][51] , 
        \inq_ary[4][52] , \inq_ary[4][53] , \inq_ary[4][54] , \inq_ary[4][55] , 
        \inq_ary[4][56] , \inq_ary[4][57] , \inq_ary[4][58] , \inq_ary[4][59] , 
        \inq_ary[4][60] , \inq_ary[4][61] , \inq_ary[4][62] , \inq_ary[4][63] , 
        \inq_ary[4][64] , \inq_ary[4][65] , \inq_ary[4][66] , \inq_ary[4][67] , 
        \inq_ary[4][68] , \inq_ary[4][69] , \inq_ary[4][70] , \inq_ary[4][71] , 
        \inq_ary[4][72] , \inq_ary[4][73] , \inq_ary[4][74] , \inq_ary[4][75] , 
        \inq_ary[4][76] , \inq_ary[4][77] , \inq_ary[4][78] , \inq_ary[4][79] , 
        \inq_ary[4][80] , \inq_ary[4][81] , \inq_ary[4][82] , \inq_ary[4][83] , 
        \inq_ary[4][84] , \inq_ary[4][85] , \inq_ary[4][86] , \inq_ary[4][87] , 
        \inq_ary[4][88] , \inq_ary[4][89] , \inq_ary[4][90] , \inq_ary[4][91] , 
        \inq_ary[4][92] , \inq_ary[4][93] , \inq_ary[4][94] , \inq_ary[4][95] , 
        \inq_ary[4][96] , \inq_ary[4][97] , \inq_ary[4][98] , \inq_ary[4][99] , 
        \inq_ary[4][100] , \inq_ary[4][101] , \inq_ary[4][102] , 
        \inq_ary[4][103] , \inq_ary[4][104] , \inq_ary[4][105] , 
        \inq_ary[4][106] , \inq_ary[4][107] , \inq_ary[4][108] , 
        \inq_ary[4][109] , \inq_ary[4][110] , \inq_ary[4][111] , 
        \inq_ary[4][112] , \inq_ary[4][113] , \inq_ary[4][114] , 
        \inq_ary[4][115] , \inq_ary[4][116] , \inq_ary[4][117] , 
        \inq_ary[4][118] , \inq_ary[4][119] , \inq_ary[4][120] , 
        \inq_ary[4][121] , \inq_ary[4][122] , \inq_ary[4][123] , 
        \inq_ary[4][124] , \inq_ary[4][125] , \inq_ary[4][126] , 
        \inq_ary[4][127] , \inq_ary[4][128] , \inq_ary[4][129] , 
        \inq_ary[4][130] , \inq_ary[4][131] , \inq_ary[4][132] , 
        \inq_ary[4][133] , \inq_ary[4][134] , \inq_ary[4][135] , 
        \inq_ary[4][136] , \inq_ary[4][137] , \inq_ary[4][138] , 
        \inq_ary[4][139] , \inq_ary[4][140] , \inq_ary[4][141] , 
        \inq_ary[4][142] , \inq_ary[4][143] , \inq_ary[4][144] , 
        \inq_ary[4][145] , \inq_ary[4][146] , \inq_ary[4][147] , 
        \inq_ary[4][148] , \inq_ary[4][149] , \inq_ary[4][150] , 
        \inq_ary[4][151] , \inq_ary[4][152] , \inq_ary[4][153] , 
        \inq_ary[4][154] , \inq_ary[4][155] , \inq_ary[4][156] , 
        \inq_ary[4][157] , \inq_ary[4][158] , \inq_ary[4][159] }), .D5({
        \inq_ary[5][0] , \inq_ary[5][1] , \inq_ary[5][2] , \inq_ary[5][3] , 
        \inq_ary[5][4] , \inq_ary[5][5] , \inq_ary[5][6] , \inq_ary[5][7] , 
        \inq_ary[5][8] , \inq_ary[5][9] , \inq_ary[5][10] , \inq_ary[5][11] , 
        \inq_ary[5][12] , \inq_ary[5][13] , \inq_ary[5][14] , \inq_ary[5][15] , 
        \inq_ary[5][16] , \inq_ary[5][17] , \inq_ary[5][18] , \inq_ary[5][19] , 
        \inq_ary[5][20] , \inq_ary[5][21] , \inq_ary[5][22] , \inq_ary[5][23] , 
        \inq_ary[5][24] , \inq_ary[5][25] , \inq_ary[5][26] , \inq_ary[5][27] , 
        \inq_ary[5][28] , \inq_ary[5][29] , \inq_ary[5][30] , \inq_ary[5][31] , 
        \inq_ary[5][32] , \inq_ary[5][33] , \inq_ary[5][34] , \inq_ary[5][35] , 
        \inq_ary[5][36] , \inq_ary[5][37] , \inq_ary[5][38] , \inq_ary[5][39] , 
        \inq_ary[5][40] , \inq_ary[5][41] , \inq_ary[5][42] , \inq_ary[5][43] , 
        \inq_ary[5][44] , \inq_ary[5][45] , \inq_ary[5][46] , \inq_ary[5][47] , 
        \inq_ary[5][48] , \inq_ary[5][49] , \inq_ary[5][50] , \inq_ary[5][51] , 
        \inq_ary[5][52] , \inq_ary[5][53] , \inq_ary[5][54] , \inq_ary[5][55] , 
        \inq_ary[5][56] , \inq_ary[5][57] , \inq_ary[5][58] , \inq_ary[5][59] , 
        \inq_ary[5][60] , \inq_ary[5][61] , \inq_ary[5][62] , \inq_ary[5][63] , 
        \inq_ary[5][64] , \inq_ary[5][65] , \inq_ary[5][66] , \inq_ary[5][67] , 
        \inq_ary[5][68] , \inq_ary[5][69] , \inq_ary[5][70] , \inq_ary[5][71] , 
        \inq_ary[5][72] , \inq_ary[5][73] , \inq_ary[5][74] , \inq_ary[5][75] , 
        \inq_ary[5][76] , \inq_ary[5][77] , \inq_ary[5][78] , \inq_ary[5][79] , 
        \inq_ary[5][80] , \inq_ary[5][81] , \inq_ary[5][82] , \inq_ary[5][83] , 
        \inq_ary[5][84] , \inq_ary[5][85] , \inq_ary[5][86] , \inq_ary[5][87] , 
        \inq_ary[5][88] , \inq_ary[5][89] , \inq_ary[5][90] , \inq_ary[5][91] , 
        \inq_ary[5][92] , \inq_ary[5][93] , \inq_ary[5][94] , \inq_ary[5][95] , 
        \inq_ary[5][96] , \inq_ary[5][97] , \inq_ary[5][98] , \inq_ary[5][99] , 
        \inq_ary[5][100] , \inq_ary[5][101] , \inq_ary[5][102] , 
        \inq_ary[5][103] , \inq_ary[5][104] , \inq_ary[5][105] , 
        \inq_ary[5][106] , \inq_ary[5][107] , \inq_ary[5][108] , 
        \inq_ary[5][109] , \inq_ary[5][110] , \inq_ary[5][111] , 
        \inq_ary[5][112] , \inq_ary[5][113] , \inq_ary[5][114] , 
        \inq_ary[5][115] , \inq_ary[5][116] , \inq_ary[5][117] , 
        \inq_ary[5][118] , \inq_ary[5][119] , \inq_ary[5][120] , 
        \inq_ary[5][121] , \inq_ary[5][122] , \inq_ary[5][123] , 
        \inq_ary[5][124] , \inq_ary[5][125] , \inq_ary[5][126] , 
        \inq_ary[5][127] , \inq_ary[5][128] , \inq_ary[5][129] , 
        \inq_ary[5][130] , \inq_ary[5][131] , \inq_ary[5][132] , 
        \inq_ary[5][133] , \inq_ary[5][134] , \inq_ary[5][135] , 
        \inq_ary[5][136] , \inq_ary[5][137] , \inq_ary[5][138] , 
        \inq_ary[5][139] , \inq_ary[5][140] , \inq_ary[5][141] , 
        \inq_ary[5][142] , \inq_ary[5][143] , \inq_ary[5][144] , 
        \inq_ary[5][145] , \inq_ary[5][146] , \inq_ary[5][147] , 
        \inq_ary[5][148] , \inq_ary[5][149] , \inq_ary[5][150] , 
        \inq_ary[5][151] , \inq_ary[5][152] , \inq_ary[5][153] , 
        \inq_ary[5][154] , \inq_ary[5][155] , \inq_ary[5][156] , 
        \inq_ary[5][157] , \inq_ary[5][158] , \inq_ary[5][159] }), .D6({
        \inq_ary[6][0] , \inq_ary[6][1] , \inq_ary[6][2] , \inq_ary[6][3] , 
        \inq_ary[6][4] , \inq_ary[6][5] , \inq_ary[6][6] , \inq_ary[6][7] , 
        \inq_ary[6][8] , \inq_ary[6][9] , \inq_ary[6][10] , \inq_ary[6][11] , 
        \inq_ary[6][12] , \inq_ary[6][13] , \inq_ary[6][14] , \inq_ary[6][15] , 
        \inq_ary[6][16] , \inq_ary[6][17] , \inq_ary[6][18] , \inq_ary[6][19] , 
        \inq_ary[6][20] , \inq_ary[6][21] , \inq_ary[6][22] , \inq_ary[6][23] , 
        \inq_ary[6][24] , \inq_ary[6][25] , \inq_ary[6][26] , \inq_ary[6][27] , 
        \inq_ary[6][28] , \inq_ary[6][29] , \inq_ary[6][30] , \inq_ary[6][31] , 
        \inq_ary[6][32] , \inq_ary[6][33] , \inq_ary[6][34] , \inq_ary[6][35] , 
        \inq_ary[6][36] , \inq_ary[6][37] , \inq_ary[6][38] , \inq_ary[6][39] , 
        \inq_ary[6][40] , \inq_ary[6][41] , \inq_ary[6][42] , \inq_ary[6][43] , 
        \inq_ary[6][44] , \inq_ary[6][45] , \inq_ary[6][46] , \inq_ary[6][47] , 
        \inq_ary[6][48] , \inq_ary[6][49] , \inq_ary[6][50] , \inq_ary[6][51] , 
        \inq_ary[6][52] , \inq_ary[6][53] , \inq_ary[6][54] , \inq_ary[6][55] , 
        \inq_ary[6][56] , \inq_ary[6][57] , \inq_ary[6][58] , \inq_ary[6][59] , 
        \inq_ary[6][60] , \inq_ary[6][61] , \inq_ary[6][62] , \inq_ary[6][63] , 
        \inq_ary[6][64] , \inq_ary[6][65] , \inq_ary[6][66] , \inq_ary[6][67] , 
        \inq_ary[6][68] , \inq_ary[6][69] , \inq_ary[6][70] , \inq_ary[6][71] , 
        \inq_ary[6][72] , \inq_ary[6][73] , \inq_ary[6][74] , \inq_ary[6][75] , 
        \inq_ary[6][76] , \inq_ary[6][77] , \inq_ary[6][78] , \inq_ary[6][79] , 
        \inq_ary[6][80] , \inq_ary[6][81] , \inq_ary[6][82] , \inq_ary[6][83] , 
        \inq_ary[6][84] , \inq_ary[6][85] , \inq_ary[6][86] , \inq_ary[6][87] , 
        \inq_ary[6][88] , \inq_ary[6][89] , \inq_ary[6][90] , \inq_ary[6][91] , 
        \inq_ary[6][92] , \inq_ary[6][93] , \inq_ary[6][94] , \inq_ary[6][95] , 
        \inq_ary[6][96] , \inq_ary[6][97] , \inq_ary[6][98] , \inq_ary[6][99] , 
        \inq_ary[6][100] , \inq_ary[6][101] , \inq_ary[6][102] , 
        \inq_ary[6][103] , \inq_ary[6][104] , \inq_ary[6][105] , 
        \inq_ary[6][106] , \inq_ary[6][107] , \inq_ary[6][108] , 
        \inq_ary[6][109] , \inq_ary[6][110] , \inq_ary[6][111] , 
        \inq_ary[6][112] , \inq_ary[6][113] , \inq_ary[6][114] , 
        \inq_ary[6][115] , \inq_ary[6][116] , \inq_ary[6][117] , 
        \inq_ary[6][118] , \inq_ary[6][119] , \inq_ary[6][120] , 
        \inq_ary[6][121] , \inq_ary[6][122] , \inq_ary[6][123] , 
        \inq_ary[6][124] , \inq_ary[6][125] , \inq_ary[6][126] , 
        \inq_ary[6][127] , \inq_ary[6][128] , \inq_ary[6][129] , 
        \inq_ary[6][130] , \inq_ary[6][131] , \inq_ary[6][132] , 
        \inq_ary[6][133] , \inq_ary[6][134] , \inq_ary[6][135] , 
        \inq_ary[6][136] , \inq_ary[6][137] , \inq_ary[6][138] , 
        \inq_ary[6][139] , \inq_ary[6][140] , \inq_ary[6][141] , 
        \inq_ary[6][142] , \inq_ary[6][143] , \inq_ary[6][144] , 
        \inq_ary[6][145] , \inq_ary[6][146] , \inq_ary[6][147] , 
        \inq_ary[6][148] , \inq_ary[6][149] , \inq_ary[6][150] , 
        \inq_ary[6][151] , \inq_ary[6][152] , \inq_ary[6][153] , 
        \inq_ary[6][154] , \inq_ary[6][155] , \inq_ary[6][156] , 
        \inq_ary[6][157] , \inq_ary[6][158] , \inq_ary[6][159] }), .D7({
        \inq_ary[7][0] , \inq_ary[7][1] , \inq_ary[7][2] , \inq_ary[7][3] , 
        \inq_ary[7][4] , \inq_ary[7][5] , \inq_ary[7][6] , \inq_ary[7][7] , 
        \inq_ary[7][8] , \inq_ary[7][9] , \inq_ary[7][10] , \inq_ary[7][11] , 
        \inq_ary[7][12] , \inq_ary[7][13] , \inq_ary[7][14] , \inq_ary[7][15] , 
        \inq_ary[7][16] , \inq_ary[7][17] , \inq_ary[7][18] , \inq_ary[7][19] , 
        \inq_ary[7][20] , \inq_ary[7][21] , \inq_ary[7][22] , \inq_ary[7][23] , 
        \inq_ary[7][24] , \inq_ary[7][25] , \inq_ary[7][26] , \inq_ary[7][27] , 
        \inq_ary[7][28] , \inq_ary[7][29] , \inq_ary[7][30] , \inq_ary[7][31] , 
        \inq_ary[7][32] , \inq_ary[7][33] , \inq_ary[7][34] , \inq_ary[7][35] , 
        \inq_ary[7][36] , \inq_ary[7][37] , \inq_ary[7][38] , \inq_ary[7][39] , 
        \inq_ary[7][40] , \inq_ary[7][41] , \inq_ary[7][42] , \inq_ary[7][43] , 
        \inq_ary[7][44] , \inq_ary[7][45] , \inq_ary[7][46] , \inq_ary[7][47] , 
        \inq_ary[7][48] , \inq_ary[7][49] , \inq_ary[7][50] , \inq_ary[7][51] , 
        \inq_ary[7][52] , \inq_ary[7][53] , \inq_ary[7][54] , \inq_ary[7][55] , 
        \inq_ary[7][56] , \inq_ary[7][57] , \inq_ary[7][58] , \inq_ary[7][59] , 
        \inq_ary[7][60] , \inq_ary[7][61] , \inq_ary[7][62] , \inq_ary[7][63] , 
        \inq_ary[7][64] , \inq_ary[7][65] , \inq_ary[7][66] , \inq_ary[7][67] , 
        \inq_ary[7][68] , \inq_ary[7][69] , \inq_ary[7][70] , \inq_ary[7][71] , 
        \inq_ary[7][72] , \inq_ary[7][73] , \inq_ary[7][74] , \inq_ary[7][75] , 
        \inq_ary[7][76] , \inq_ary[7][77] , \inq_ary[7][78] , \inq_ary[7][79] , 
        \inq_ary[7][80] , \inq_ary[7][81] , \inq_ary[7][82] , \inq_ary[7][83] , 
        \inq_ary[7][84] , \inq_ary[7][85] , \inq_ary[7][86] , \inq_ary[7][87] , 
        \inq_ary[7][88] , \inq_ary[7][89] , \inq_ary[7][90] , \inq_ary[7][91] , 
        \inq_ary[7][92] , \inq_ary[7][93] , \inq_ary[7][94] , \inq_ary[7][95] , 
        \inq_ary[7][96] , \inq_ary[7][97] , \inq_ary[7][98] , \inq_ary[7][99] , 
        \inq_ary[7][100] , \inq_ary[7][101] , \inq_ary[7][102] , 
        \inq_ary[7][103] , \inq_ary[7][104] , \inq_ary[7][105] , 
        \inq_ary[7][106] , \inq_ary[7][107] , \inq_ary[7][108] , 
        \inq_ary[7][109] , \inq_ary[7][110] , \inq_ary[7][111] , 
        \inq_ary[7][112] , \inq_ary[7][113] , \inq_ary[7][114] , 
        \inq_ary[7][115] , \inq_ary[7][116] , \inq_ary[7][117] , 
        \inq_ary[7][118] , \inq_ary[7][119] , \inq_ary[7][120] , 
        \inq_ary[7][121] , \inq_ary[7][122] , \inq_ary[7][123] , 
        \inq_ary[7][124] , \inq_ary[7][125] , \inq_ary[7][126] , 
        \inq_ary[7][127] , \inq_ary[7][128] , \inq_ary[7][129] , 
        \inq_ary[7][130] , \inq_ary[7][131] , \inq_ary[7][132] , 
        \inq_ary[7][133] , \inq_ary[7][134] , \inq_ary[7][135] , 
        \inq_ary[7][136] , \inq_ary[7][137] , \inq_ary[7][138] , 
        \inq_ary[7][139] , \inq_ary[7][140] , \inq_ary[7][141] , 
        \inq_ary[7][142] , \inq_ary[7][143] , \inq_ary[7][144] , 
        \inq_ary[7][145] , \inq_ary[7][146] , \inq_ary[7][147] , 
        \inq_ary[7][148] , \inq_ary[7][149] , \inq_ary[7][150] , 
        \inq_ary[7][151] , \inq_ary[7][152] , \inq_ary[7][153] , 
        \inq_ary[7][154] , \inq_ary[7][155] , \inq_ary[7][156] , 
        \inq_ary[7][157] , \inq_ary[7][158] , \inq_ary[7][159] }), .D8({
        \inq_ary[8][0] , \inq_ary[8][1] , \inq_ary[8][2] , \inq_ary[8][3] , 
        \inq_ary[8][4] , \inq_ary[8][5] , \inq_ary[8][6] , \inq_ary[8][7] , 
        \inq_ary[8][8] , \inq_ary[8][9] , \inq_ary[8][10] , \inq_ary[8][11] , 
        \inq_ary[8][12] , \inq_ary[8][13] , \inq_ary[8][14] , \inq_ary[8][15] , 
        \inq_ary[8][16] , \inq_ary[8][17] , \inq_ary[8][18] , \inq_ary[8][19] , 
        \inq_ary[8][20] , \inq_ary[8][21] , \inq_ary[8][22] , \inq_ary[8][23] , 
        \inq_ary[8][24] , \inq_ary[8][25] , \inq_ary[8][26] , \inq_ary[8][27] , 
        \inq_ary[8][28] , \inq_ary[8][29] , \inq_ary[8][30] , \inq_ary[8][31] , 
        \inq_ary[8][32] , \inq_ary[8][33] , \inq_ary[8][34] , \inq_ary[8][35] , 
        \inq_ary[8][36] , \inq_ary[8][37] , \inq_ary[8][38] , \inq_ary[8][39] , 
        \inq_ary[8][40] , \inq_ary[8][41] , \inq_ary[8][42] , \inq_ary[8][43] , 
        \inq_ary[8][44] , \inq_ary[8][45] , \inq_ary[8][46] , \inq_ary[8][47] , 
        \inq_ary[8][48] , \inq_ary[8][49] , \inq_ary[8][50] , \inq_ary[8][51] , 
        \inq_ary[8][52] , \inq_ary[8][53] , \inq_ary[8][54] , \inq_ary[8][55] , 
        \inq_ary[8][56] , \inq_ary[8][57] , \inq_ary[8][58] , \inq_ary[8][59] , 
        \inq_ary[8][60] , \inq_ary[8][61] , \inq_ary[8][62] , \inq_ary[8][63] , 
        \inq_ary[8][64] , \inq_ary[8][65] , \inq_ary[8][66] , \inq_ary[8][67] , 
        \inq_ary[8][68] , \inq_ary[8][69] , \inq_ary[8][70] , \inq_ary[8][71] , 
        \inq_ary[8][72] , \inq_ary[8][73] , \inq_ary[8][74] , \inq_ary[8][75] , 
        \inq_ary[8][76] , \inq_ary[8][77] , \inq_ary[8][78] , \inq_ary[8][79] , 
        \inq_ary[8][80] , \inq_ary[8][81] , \inq_ary[8][82] , \inq_ary[8][83] , 
        \inq_ary[8][84] , \inq_ary[8][85] , \inq_ary[8][86] , \inq_ary[8][87] , 
        \inq_ary[8][88] , \inq_ary[8][89] , \inq_ary[8][90] , \inq_ary[8][91] , 
        \inq_ary[8][92] , \inq_ary[8][93] , \inq_ary[8][94] , \inq_ary[8][95] , 
        \inq_ary[8][96] , \inq_ary[8][97] , \inq_ary[8][98] , \inq_ary[8][99] , 
        \inq_ary[8][100] , \inq_ary[8][101] , \inq_ary[8][102] , 
        \inq_ary[8][103] , \inq_ary[8][104] , \inq_ary[8][105] , 
        \inq_ary[8][106] , \inq_ary[8][107] , \inq_ary[8][108] , 
        \inq_ary[8][109] , \inq_ary[8][110] , \inq_ary[8][111] , 
        \inq_ary[8][112] , \inq_ary[8][113] , \inq_ary[8][114] , 
        \inq_ary[8][115] , \inq_ary[8][116] , \inq_ary[8][117] , 
        \inq_ary[8][118] , \inq_ary[8][119] , \inq_ary[8][120] , 
        \inq_ary[8][121] , \inq_ary[8][122] , \inq_ary[8][123] , 
        \inq_ary[8][124] , \inq_ary[8][125] , \inq_ary[8][126] , 
        \inq_ary[8][127] , \inq_ary[8][128] , \inq_ary[8][129] , 
        \inq_ary[8][130] , \inq_ary[8][131] , \inq_ary[8][132] , 
        \inq_ary[8][133] , \inq_ary[8][134] , \inq_ary[8][135] , 
        \inq_ary[8][136] , \inq_ary[8][137] , \inq_ary[8][138] , 
        \inq_ary[8][139] , \inq_ary[8][140] , \inq_ary[8][141] , 
        \inq_ary[8][142] , \inq_ary[8][143] , \inq_ary[8][144] , 
        \inq_ary[8][145] , \inq_ary[8][146] , \inq_ary[8][147] , 
        \inq_ary[8][148] , \inq_ary[8][149] , \inq_ary[8][150] , 
        \inq_ary[8][151] , \inq_ary[8][152] , \inq_ary[8][153] , 
        \inq_ary[8][154] , \inq_ary[8][155] , \inq_ary[8][156] , 
        \inq_ary[8][157] , \inq_ary[8][158] , \inq_ary[8][159] }), .D9({
        \inq_ary[9][0] , \inq_ary[9][1] , \inq_ary[9][2] , \inq_ary[9][3] , 
        \inq_ary[9][4] , \inq_ary[9][5] , \inq_ary[9][6] , \inq_ary[9][7] , 
        \inq_ary[9][8] , \inq_ary[9][9] , \inq_ary[9][10] , \inq_ary[9][11] , 
        \inq_ary[9][12] , \inq_ary[9][13] , \inq_ary[9][14] , \inq_ary[9][15] , 
        \inq_ary[9][16] , \inq_ary[9][17] , \inq_ary[9][18] , \inq_ary[9][19] , 
        \inq_ary[9][20] , \inq_ary[9][21] , \inq_ary[9][22] , \inq_ary[9][23] , 
        \inq_ary[9][24] , \inq_ary[9][25] , \inq_ary[9][26] , \inq_ary[9][27] , 
        \inq_ary[9][28] , \inq_ary[9][29] , \inq_ary[9][30] , \inq_ary[9][31] , 
        \inq_ary[9][32] , \inq_ary[9][33] , \inq_ary[9][34] , \inq_ary[9][35] , 
        \inq_ary[9][36] , \inq_ary[9][37] , \inq_ary[9][38] , \inq_ary[9][39] , 
        \inq_ary[9][40] , \inq_ary[9][41] , \inq_ary[9][42] , \inq_ary[9][43] , 
        \inq_ary[9][44] , \inq_ary[9][45] , \inq_ary[9][46] , \inq_ary[9][47] , 
        \inq_ary[9][48] , \inq_ary[9][49] , \inq_ary[9][50] , \inq_ary[9][51] , 
        \inq_ary[9][52] , \inq_ary[9][53] , \inq_ary[9][54] , \inq_ary[9][55] , 
        \inq_ary[9][56] , \inq_ary[9][57] , \inq_ary[9][58] , \inq_ary[9][59] , 
        \inq_ary[9][60] , \inq_ary[9][61] , \inq_ary[9][62] , \inq_ary[9][63] , 
        \inq_ary[9][64] , \inq_ary[9][65] , \inq_ary[9][66] , \inq_ary[9][67] , 
        \inq_ary[9][68] , \inq_ary[9][69] , \inq_ary[9][70] , \inq_ary[9][71] , 
        \inq_ary[9][72] , \inq_ary[9][73] , \inq_ary[9][74] , \inq_ary[9][75] , 
        \inq_ary[9][76] , \inq_ary[9][77] , \inq_ary[9][78] , \inq_ary[9][79] , 
        \inq_ary[9][80] , \inq_ary[9][81] , \inq_ary[9][82] , \inq_ary[9][83] , 
        \inq_ary[9][84] , \inq_ary[9][85] , \inq_ary[9][86] , \inq_ary[9][87] , 
        \inq_ary[9][88] , \inq_ary[9][89] , \inq_ary[9][90] , \inq_ary[9][91] , 
        \inq_ary[9][92] , \inq_ary[9][93] , \inq_ary[9][94] , \inq_ary[9][95] , 
        \inq_ary[9][96] , \inq_ary[9][97] , \inq_ary[9][98] , \inq_ary[9][99] , 
        \inq_ary[9][100] , \inq_ary[9][101] , \inq_ary[9][102] , 
        \inq_ary[9][103] , \inq_ary[9][104] , \inq_ary[9][105] , 
        \inq_ary[9][106] , \inq_ary[9][107] , \inq_ary[9][108] , 
        \inq_ary[9][109] , \inq_ary[9][110] , \inq_ary[9][111] , 
        \inq_ary[9][112] , \inq_ary[9][113] , \inq_ary[9][114] , 
        \inq_ary[9][115] , \inq_ary[9][116] , \inq_ary[9][117] , 
        \inq_ary[9][118] , \inq_ary[9][119] , \inq_ary[9][120] , 
        \inq_ary[9][121] , \inq_ary[9][122] , \inq_ary[9][123] , 
        \inq_ary[9][124] , \inq_ary[9][125] , \inq_ary[9][126] , 
        \inq_ary[9][127] , \inq_ary[9][128] , \inq_ary[9][129] , 
        \inq_ary[9][130] , \inq_ary[9][131] , \inq_ary[9][132] , 
        \inq_ary[9][133] , \inq_ary[9][134] , \inq_ary[9][135] , 
        \inq_ary[9][136] , \inq_ary[9][137] , \inq_ary[9][138] , 
        \inq_ary[9][139] , \inq_ary[9][140] , \inq_ary[9][141] , 
        \inq_ary[9][142] , \inq_ary[9][143] , \inq_ary[9][144] , 
        \inq_ary[9][145] , \inq_ary[9][146] , \inq_ary[9][147] , 
        \inq_ary[9][148] , \inq_ary[9][149] , \inq_ary[9][150] , 
        \inq_ary[9][151] , \inq_ary[9][152] , \inq_ary[9][153] , 
        \inq_ary[9][154] , \inq_ary[9][155] , \inq_ary[9][156] , 
        \inq_ary[9][157] , \inq_ary[9][158] , \inq_ary[9][159] }), .D10({
        \inq_ary[10][0] , \inq_ary[10][1] , \inq_ary[10][2] , \inq_ary[10][3] , 
        \inq_ary[10][4] , \inq_ary[10][5] , \inq_ary[10][6] , \inq_ary[10][7] , 
        \inq_ary[10][8] , \inq_ary[10][9] , \inq_ary[10][10] , 
        \inq_ary[10][11] , \inq_ary[10][12] , \inq_ary[10][13] , 
        \inq_ary[10][14] , \inq_ary[10][15] , \inq_ary[10][16] , 
        \inq_ary[10][17] , \inq_ary[10][18] , \inq_ary[10][19] , 
        \inq_ary[10][20] , \inq_ary[10][21] , \inq_ary[10][22] , 
        \inq_ary[10][23] , \inq_ary[10][24] , \inq_ary[10][25] , 
        \inq_ary[10][26] , \inq_ary[10][27] , \inq_ary[10][28] , 
        \inq_ary[10][29] , \inq_ary[10][30] , \inq_ary[10][31] , 
        \inq_ary[10][32] , \inq_ary[10][33] , \inq_ary[10][34] , 
        \inq_ary[10][35] , \inq_ary[10][36] , \inq_ary[10][37] , 
        \inq_ary[10][38] , \inq_ary[10][39] , \inq_ary[10][40] , 
        \inq_ary[10][41] , \inq_ary[10][42] , \inq_ary[10][43] , 
        \inq_ary[10][44] , \inq_ary[10][45] , \inq_ary[10][46] , 
        \inq_ary[10][47] , \inq_ary[10][48] , \inq_ary[10][49] , 
        \inq_ary[10][50] , \inq_ary[10][51] , \inq_ary[10][52] , 
        \inq_ary[10][53] , \inq_ary[10][54] , \inq_ary[10][55] , 
        \inq_ary[10][56] , \inq_ary[10][57] , \inq_ary[10][58] , 
        \inq_ary[10][59] , \inq_ary[10][60] , \inq_ary[10][61] , 
        \inq_ary[10][62] , \inq_ary[10][63] , \inq_ary[10][64] , 
        \inq_ary[10][65] , \inq_ary[10][66] , \inq_ary[10][67] , 
        \inq_ary[10][68] , \inq_ary[10][69] , \inq_ary[10][70] , 
        \inq_ary[10][71] , \inq_ary[10][72] , \inq_ary[10][73] , 
        \inq_ary[10][74] , \inq_ary[10][75] , \inq_ary[10][76] , 
        \inq_ary[10][77] , \inq_ary[10][78] , \inq_ary[10][79] , 
        \inq_ary[10][80] , \inq_ary[10][81] , \inq_ary[10][82] , 
        \inq_ary[10][83] , \inq_ary[10][84] , \inq_ary[10][85] , 
        \inq_ary[10][86] , \inq_ary[10][87] , \inq_ary[10][88] , 
        \inq_ary[10][89] , \inq_ary[10][90] , \inq_ary[10][91] , 
        \inq_ary[10][92] , \inq_ary[10][93] , \inq_ary[10][94] , 
        \inq_ary[10][95] , \inq_ary[10][96] , \inq_ary[10][97] , 
        \inq_ary[10][98] , \inq_ary[10][99] , \inq_ary[10][100] , 
        \inq_ary[10][101] , \inq_ary[10][102] , \inq_ary[10][103] , 
        \inq_ary[10][104] , \inq_ary[10][105] , \inq_ary[10][106] , 
        \inq_ary[10][107] , \inq_ary[10][108] , \inq_ary[10][109] , 
        \inq_ary[10][110] , \inq_ary[10][111] , \inq_ary[10][112] , 
        \inq_ary[10][113] , \inq_ary[10][114] , \inq_ary[10][115] , 
        \inq_ary[10][116] , \inq_ary[10][117] , \inq_ary[10][118] , 
        \inq_ary[10][119] , \inq_ary[10][120] , \inq_ary[10][121] , 
        \inq_ary[10][122] , \inq_ary[10][123] , \inq_ary[10][124] , 
        \inq_ary[10][125] , \inq_ary[10][126] , \inq_ary[10][127] , 
        \inq_ary[10][128] , \inq_ary[10][129] , \inq_ary[10][130] , 
        \inq_ary[10][131] , \inq_ary[10][132] , \inq_ary[10][133] , 
        \inq_ary[10][134] , \inq_ary[10][135] , \inq_ary[10][136] , 
        \inq_ary[10][137] , \inq_ary[10][138] , \inq_ary[10][139] , 
        \inq_ary[10][140] , \inq_ary[10][141] , \inq_ary[10][142] , 
        \inq_ary[10][143] , \inq_ary[10][144] , \inq_ary[10][145] , 
        \inq_ary[10][146] , \inq_ary[10][147] , \inq_ary[10][148] , 
        \inq_ary[10][149] , \inq_ary[10][150] , \inq_ary[10][151] , 
        \inq_ary[10][152] , \inq_ary[10][153] , \inq_ary[10][154] , 
        \inq_ary[10][155] , \inq_ary[10][156] , \inq_ary[10][157] , 
        \inq_ary[10][158] , \inq_ary[10][159] }), .D11({\inq_ary[11][0] , 
        \inq_ary[11][1] , \inq_ary[11][2] , \inq_ary[11][3] , \inq_ary[11][4] , 
        \inq_ary[11][5] , \inq_ary[11][6] , \inq_ary[11][7] , \inq_ary[11][8] , 
        \inq_ary[11][9] , \inq_ary[11][10] , \inq_ary[11][11] , 
        \inq_ary[11][12] , \inq_ary[11][13] , \inq_ary[11][14] , 
        \inq_ary[11][15] , \inq_ary[11][16] , \inq_ary[11][17] , 
        \inq_ary[11][18] , \inq_ary[11][19] , \inq_ary[11][20] , 
        \inq_ary[11][21] , \inq_ary[11][22] , \inq_ary[11][23] , 
        \inq_ary[11][24] , \inq_ary[11][25] , \inq_ary[11][26] , 
        \inq_ary[11][27] , \inq_ary[11][28] , \inq_ary[11][29] , 
        \inq_ary[11][30] , \inq_ary[11][31] , \inq_ary[11][32] , 
        \inq_ary[11][33] , \inq_ary[11][34] , \inq_ary[11][35] , 
        \inq_ary[11][36] , \inq_ary[11][37] , \inq_ary[11][38] , 
        \inq_ary[11][39] , \inq_ary[11][40] , \inq_ary[11][41] , 
        \inq_ary[11][42] , \inq_ary[11][43] , \inq_ary[11][44] , 
        \inq_ary[11][45] , \inq_ary[11][46] , \inq_ary[11][47] , 
        \inq_ary[11][48] , \inq_ary[11][49] , \inq_ary[11][50] , 
        \inq_ary[11][51] , \inq_ary[11][52] , \inq_ary[11][53] , 
        \inq_ary[11][54] , \inq_ary[11][55] , \inq_ary[11][56] , 
        \inq_ary[11][57] , \inq_ary[11][58] , \inq_ary[11][59] , 
        \inq_ary[11][60] , \inq_ary[11][61] , \inq_ary[11][62] , 
        \inq_ary[11][63] , \inq_ary[11][64] , \inq_ary[11][65] , 
        \inq_ary[11][66] , \inq_ary[11][67] , \inq_ary[11][68] , 
        \inq_ary[11][69] , \inq_ary[11][70] , \inq_ary[11][71] , 
        \inq_ary[11][72] , \inq_ary[11][73] , \inq_ary[11][74] , 
        \inq_ary[11][75] , \inq_ary[11][76] , \inq_ary[11][77] , 
        \inq_ary[11][78] , \inq_ary[11][79] , \inq_ary[11][80] , 
        \inq_ary[11][81] , \inq_ary[11][82] , \inq_ary[11][83] , 
        \inq_ary[11][84] , \inq_ary[11][85] , \inq_ary[11][86] , 
        \inq_ary[11][87] , \inq_ary[11][88] , \inq_ary[11][89] , 
        \inq_ary[11][90] , \inq_ary[11][91] , \inq_ary[11][92] , 
        \inq_ary[11][93] , \inq_ary[11][94] , \inq_ary[11][95] , 
        \inq_ary[11][96] , \inq_ary[11][97] , \inq_ary[11][98] , 
        \inq_ary[11][99] , \inq_ary[11][100] , \inq_ary[11][101] , 
        \inq_ary[11][102] , \inq_ary[11][103] , \inq_ary[11][104] , 
        \inq_ary[11][105] , \inq_ary[11][106] , \inq_ary[11][107] , 
        \inq_ary[11][108] , \inq_ary[11][109] , \inq_ary[11][110] , 
        \inq_ary[11][111] , \inq_ary[11][112] , \inq_ary[11][113] , 
        \inq_ary[11][114] , \inq_ary[11][115] , \inq_ary[11][116] , 
        \inq_ary[11][117] , \inq_ary[11][118] , \inq_ary[11][119] , 
        \inq_ary[11][120] , \inq_ary[11][121] , \inq_ary[11][122] , 
        \inq_ary[11][123] , \inq_ary[11][124] , \inq_ary[11][125] , 
        \inq_ary[11][126] , \inq_ary[11][127] , \inq_ary[11][128] , 
        \inq_ary[11][129] , \inq_ary[11][130] , \inq_ary[11][131] , 
        \inq_ary[11][132] , \inq_ary[11][133] , \inq_ary[11][134] , 
        \inq_ary[11][135] , \inq_ary[11][136] , \inq_ary[11][137] , 
        \inq_ary[11][138] , \inq_ary[11][139] , \inq_ary[11][140] , 
        \inq_ary[11][141] , \inq_ary[11][142] , \inq_ary[11][143] , 
        \inq_ary[11][144] , \inq_ary[11][145] , \inq_ary[11][146] , 
        \inq_ary[11][147] , \inq_ary[11][148] , \inq_ary[11][149] , 
        \inq_ary[11][150] , \inq_ary[11][151] , \inq_ary[11][152] , 
        \inq_ary[11][153] , \inq_ary[11][154] , \inq_ary[11][155] , 
        \inq_ary[11][156] , \inq_ary[11][157] , \inq_ary[11][158] , 
        \inq_ary[11][159] }), .D12({\inq_ary[12][0] , \inq_ary[12][1] , 
        \inq_ary[12][2] , \inq_ary[12][3] , \inq_ary[12][4] , \inq_ary[12][5] , 
        \inq_ary[12][6] , \inq_ary[12][7] , \inq_ary[12][8] , \inq_ary[12][9] , 
        \inq_ary[12][10] , \inq_ary[12][11] , \inq_ary[12][12] , 
        \inq_ary[12][13] , \inq_ary[12][14] , \inq_ary[12][15] , 
        \inq_ary[12][16] , \inq_ary[12][17] , \inq_ary[12][18] , 
        \inq_ary[12][19] , \inq_ary[12][20] , \inq_ary[12][21] , 
        \inq_ary[12][22] , \inq_ary[12][23] , \inq_ary[12][24] , 
        \inq_ary[12][25] , \inq_ary[12][26] , \inq_ary[12][27] , 
        \inq_ary[12][28] , \inq_ary[12][29] , \inq_ary[12][30] , 
        \inq_ary[12][31] , \inq_ary[12][32] , \inq_ary[12][33] , 
        \inq_ary[12][34] , \inq_ary[12][35] , \inq_ary[12][36] , 
        \inq_ary[12][37] , \inq_ary[12][38] , \inq_ary[12][39] , 
        \inq_ary[12][40] , \inq_ary[12][41] , \inq_ary[12][42] , 
        \inq_ary[12][43] , \inq_ary[12][44] , \inq_ary[12][45] , 
        \inq_ary[12][46] , \inq_ary[12][47] , \inq_ary[12][48] , 
        \inq_ary[12][49] , \inq_ary[12][50] , \inq_ary[12][51] , 
        \inq_ary[12][52] , \inq_ary[12][53] , \inq_ary[12][54] , 
        \inq_ary[12][55] , \inq_ary[12][56] , \inq_ary[12][57] , 
        \inq_ary[12][58] , \inq_ary[12][59] , \inq_ary[12][60] , 
        \inq_ary[12][61] , \inq_ary[12][62] , \inq_ary[12][63] , 
        \inq_ary[12][64] , \inq_ary[12][65] , \inq_ary[12][66] , 
        \inq_ary[12][67] , \inq_ary[12][68] , \inq_ary[12][69] , 
        \inq_ary[12][70] , \inq_ary[12][71] , \inq_ary[12][72] , 
        \inq_ary[12][73] , \inq_ary[12][74] , \inq_ary[12][75] , 
        \inq_ary[12][76] , \inq_ary[12][77] , \inq_ary[12][78] , 
        \inq_ary[12][79] , \inq_ary[12][80] , \inq_ary[12][81] , 
        \inq_ary[12][82] , \inq_ary[12][83] , \inq_ary[12][84] , 
        \inq_ary[12][85] , \inq_ary[12][86] , \inq_ary[12][87] , 
        \inq_ary[12][88] , \inq_ary[12][89] , \inq_ary[12][90] , 
        \inq_ary[12][91] , \inq_ary[12][92] , \inq_ary[12][93] , 
        \inq_ary[12][94] , \inq_ary[12][95] , \inq_ary[12][96] , 
        \inq_ary[12][97] , \inq_ary[12][98] , \inq_ary[12][99] , 
        \inq_ary[12][100] , \inq_ary[12][101] , \inq_ary[12][102] , 
        \inq_ary[12][103] , \inq_ary[12][104] , \inq_ary[12][105] , 
        \inq_ary[12][106] , \inq_ary[12][107] , \inq_ary[12][108] , 
        \inq_ary[12][109] , \inq_ary[12][110] , \inq_ary[12][111] , 
        \inq_ary[12][112] , \inq_ary[12][113] , \inq_ary[12][114] , 
        \inq_ary[12][115] , \inq_ary[12][116] , \inq_ary[12][117] , 
        \inq_ary[12][118] , \inq_ary[12][119] , \inq_ary[12][120] , 
        \inq_ary[12][121] , \inq_ary[12][122] , \inq_ary[12][123] , 
        \inq_ary[12][124] , \inq_ary[12][125] , \inq_ary[12][126] , 
        \inq_ary[12][127] , \inq_ary[12][128] , \inq_ary[12][129] , 
        \inq_ary[12][130] , \inq_ary[12][131] , \inq_ary[12][132] , 
        \inq_ary[12][133] , \inq_ary[12][134] , \inq_ary[12][135] , 
        \inq_ary[12][136] , \inq_ary[12][137] , \inq_ary[12][138] , 
        \inq_ary[12][139] , \inq_ary[12][140] , \inq_ary[12][141] , 
        \inq_ary[12][142] , \inq_ary[12][143] , \inq_ary[12][144] , 
        \inq_ary[12][145] , \inq_ary[12][146] , \inq_ary[12][147] , 
        \inq_ary[12][148] , \inq_ary[12][149] , \inq_ary[12][150] , 
        \inq_ary[12][151] , \inq_ary[12][152] , \inq_ary[12][153] , 
        \inq_ary[12][154] , \inq_ary[12][155] , \inq_ary[12][156] , 
        \inq_ary[12][157] , \inq_ary[12][158] , \inq_ary[12][159] }), .D13({
        \inq_ary[13][0] , \inq_ary[13][1] , \inq_ary[13][2] , \inq_ary[13][3] , 
        \inq_ary[13][4] , \inq_ary[13][5] , \inq_ary[13][6] , \inq_ary[13][7] , 
        \inq_ary[13][8] , \inq_ary[13][9] , \inq_ary[13][10] , 
        \inq_ary[13][11] , \inq_ary[13][12] , \inq_ary[13][13] , 
        \inq_ary[13][14] , \inq_ary[13][15] , \inq_ary[13][16] , 
        \inq_ary[13][17] , \inq_ary[13][18] , \inq_ary[13][19] , 
        \inq_ary[13][20] , \inq_ary[13][21] , \inq_ary[13][22] , 
        \inq_ary[13][23] , \inq_ary[13][24] , \inq_ary[13][25] , 
        \inq_ary[13][26] , \inq_ary[13][27] , \inq_ary[13][28] , 
        \inq_ary[13][29] , \inq_ary[13][30] , \inq_ary[13][31] , 
        \inq_ary[13][32] , \inq_ary[13][33] , \inq_ary[13][34] , 
        \inq_ary[13][35] , \inq_ary[13][36] , \inq_ary[13][37] , 
        \inq_ary[13][38] , \inq_ary[13][39] , \inq_ary[13][40] , 
        \inq_ary[13][41] , \inq_ary[13][42] , \inq_ary[13][43] , 
        \inq_ary[13][44] , \inq_ary[13][45] , \inq_ary[13][46] , 
        \inq_ary[13][47] , \inq_ary[13][48] , \inq_ary[13][49] , 
        \inq_ary[13][50] , \inq_ary[13][51] , \inq_ary[13][52] , 
        \inq_ary[13][53] , \inq_ary[13][54] , \inq_ary[13][55] , 
        \inq_ary[13][56] , \inq_ary[13][57] , \inq_ary[13][58] , 
        \inq_ary[13][59] , \inq_ary[13][60] , \inq_ary[13][61] , 
        \inq_ary[13][62] , \inq_ary[13][63] , \inq_ary[13][64] , 
        \inq_ary[13][65] , \inq_ary[13][66] , \inq_ary[13][67] , 
        \inq_ary[13][68] , \inq_ary[13][69] , \inq_ary[13][70] , 
        \inq_ary[13][71] , \inq_ary[13][72] , \inq_ary[13][73] , 
        \inq_ary[13][74] , \inq_ary[13][75] , \inq_ary[13][76] , 
        \inq_ary[13][77] , \inq_ary[13][78] , \inq_ary[13][79] , 
        \inq_ary[13][80] , \inq_ary[13][81] , \inq_ary[13][82] , 
        \inq_ary[13][83] , \inq_ary[13][84] , \inq_ary[13][85] , 
        \inq_ary[13][86] , \inq_ary[13][87] , \inq_ary[13][88] , 
        \inq_ary[13][89] , \inq_ary[13][90] , \inq_ary[13][91] , 
        \inq_ary[13][92] , \inq_ary[13][93] , \inq_ary[13][94] , 
        \inq_ary[13][95] , \inq_ary[13][96] , \inq_ary[13][97] , 
        \inq_ary[13][98] , \inq_ary[13][99] , \inq_ary[13][100] , 
        \inq_ary[13][101] , \inq_ary[13][102] , \inq_ary[13][103] , 
        \inq_ary[13][104] , \inq_ary[13][105] , \inq_ary[13][106] , 
        \inq_ary[13][107] , \inq_ary[13][108] , \inq_ary[13][109] , 
        \inq_ary[13][110] , \inq_ary[13][111] , \inq_ary[13][112] , 
        \inq_ary[13][113] , \inq_ary[13][114] , \inq_ary[13][115] , 
        \inq_ary[13][116] , \inq_ary[13][117] , \inq_ary[13][118] , 
        \inq_ary[13][119] , \inq_ary[13][120] , \inq_ary[13][121] , 
        \inq_ary[13][122] , \inq_ary[13][123] , \inq_ary[13][124] , 
        \inq_ary[13][125] , \inq_ary[13][126] , \inq_ary[13][127] , 
        \inq_ary[13][128] , \inq_ary[13][129] , \inq_ary[13][130] , 
        \inq_ary[13][131] , \inq_ary[13][132] , \inq_ary[13][133] , 
        \inq_ary[13][134] , \inq_ary[13][135] , \inq_ary[13][136] , 
        \inq_ary[13][137] , \inq_ary[13][138] , \inq_ary[13][139] , 
        \inq_ary[13][140] , \inq_ary[13][141] , \inq_ary[13][142] , 
        \inq_ary[13][143] , \inq_ary[13][144] , \inq_ary[13][145] , 
        \inq_ary[13][146] , \inq_ary[13][147] , \inq_ary[13][148] , 
        \inq_ary[13][149] , \inq_ary[13][150] , \inq_ary[13][151] , 
        \inq_ary[13][152] , \inq_ary[13][153] , \inq_ary[13][154] , 
        \inq_ary[13][155] , \inq_ary[13][156] , \inq_ary[13][157] , 
        \inq_ary[13][158] , \inq_ary[13][159] }), .D14({\inq_ary[14][0] , 
        \inq_ary[14][1] , \inq_ary[14][2] , \inq_ary[14][3] , \inq_ary[14][4] , 
        \inq_ary[14][5] , \inq_ary[14][6] , \inq_ary[14][7] , \inq_ary[14][8] , 
        \inq_ary[14][9] , \inq_ary[14][10] , \inq_ary[14][11] , 
        \inq_ary[14][12] , \inq_ary[14][13] , \inq_ary[14][14] , 
        \inq_ary[14][15] , \inq_ary[14][16] , \inq_ary[14][17] , 
        \inq_ary[14][18] , \inq_ary[14][19] , \inq_ary[14][20] , 
        \inq_ary[14][21] , \inq_ary[14][22] , \inq_ary[14][23] , 
        \inq_ary[14][24] , \inq_ary[14][25] , \inq_ary[14][26] , 
        \inq_ary[14][27] , \inq_ary[14][28] , \inq_ary[14][29] , 
        \inq_ary[14][30] , \inq_ary[14][31] , \inq_ary[14][32] , 
        \inq_ary[14][33] , \inq_ary[14][34] , \inq_ary[14][35] , 
        \inq_ary[14][36] , \inq_ary[14][37] , \inq_ary[14][38] , 
        \inq_ary[14][39] , \inq_ary[14][40] , \inq_ary[14][41] , 
        \inq_ary[14][42] , \inq_ary[14][43] , \inq_ary[14][44] , 
        \inq_ary[14][45] , \inq_ary[14][46] , \inq_ary[14][47] , 
        \inq_ary[14][48] , \inq_ary[14][49] , \inq_ary[14][50] , 
        \inq_ary[14][51] , \inq_ary[14][52] , \inq_ary[14][53] , 
        \inq_ary[14][54] , \inq_ary[14][55] , \inq_ary[14][56] , 
        \inq_ary[14][57] , \inq_ary[14][58] , \inq_ary[14][59] , 
        \inq_ary[14][60] , \inq_ary[14][61] , \inq_ary[14][62] , 
        \inq_ary[14][63] , \inq_ary[14][64] , \inq_ary[14][65] , 
        \inq_ary[14][66] , \inq_ary[14][67] , \inq_ary[14][68] , 
        \inq_ary[14][69] , \inq_ary[14][70] , \inq_ary[14][71] , 
        \inq_ary[14][72] , \inq_ary[14][73] , \inq_ary[14][74] , 
        \inq_ary[14][75] , \inq_ary[14][76] , \inq_ary[14][77] , 
        \inq_ary[14][78] , \inq_ary[14][79] , \inq_ary[14][80] , 
        \inq_ary[14][81] , \inq_ary[14][82] , \inq_ary[14][83] , 
        \inq_ary[14][84] , \inq_ary[14][85] , \inq_ary[14][86] , 
        \inq_ary[14][87] , \inq_ary[14][88] , \inq_ary[14][89] , 
        \inq_ary[14][90] , \inq_ary[14][91] , \inq_ary[14][92] , 
        \inq_ary[14][93] , \inq_ary[14][94] , \inq_ary[14][95] , 
        \inq_ary[14][96] , \inq_ary[14][97] , \inq_ary[14][98] , 
        \inq_ary[14][99] , \inq_ary[14][100] , \inq_ary[14][101] , 
        \inq_ary[14][102] , \inq_ary[14][103] , \inq_ary[14][104] , 
        \inq_ary[14][105] , \inq_ary[14][106] , \inq_ary[14][107] , 
        \inq_ary[14][108] , \inq_ary[14][109] , \inq_ary[14][110] , 
        \inq_ary[14][111] , \inq_ary[14][112] , \inq_ary[14][113] , 
        \inq_ary[14][114] , \inq_ary[14][115] , \inq_ary[14][116] , 
        \inq_ary[14][117] , \inq_ary[14][118] , \inq_ary[14][119] , 
        \inq_ary[14][120] , \inq_ary[14][121] , \inq_ary[14][122] , 
        \inq_ary[14][123] , \inq_ary[14][124] , \inq_ary[14][125] , 
        \inq_ary[14][126] , \inq_ary[14][127] , \inq_ary[14][128] , 
        \inq_ary[14][129] , \inq_ary[14][130] , \inq_ary[14][131] , 
        \inq_ary[14][132] , \inq_ary[14][133] , \inq_ary[14][134] , 
        \inq_ary[14][135] , \inq_ary[14][136] , \inq_ary[14][137] , 
        \inq_ary[14][138] , \inq_ary[14][139] , \inq_ary[14][140] , 
        \inq_ary[14][141] , \inq_ary[14][142] , \inq_ary[14][143] , 
        \inq_ary[14][144] , \inq_ary[14][145] , \inq_ary[14][146] , 
        \inq_ary[14][147] , \inq_ary[14][148] , \inq_ary[14][149] , 
        \inq_ary[14][150] , \inq_ary[14][151] , \inq_ary[14][152] , 
        \inq_ary[14][153] , \inq_ary[14][154] , \inq_ary[14][155] , 
        \inq_ary[14][156] , \inq_ary[14][157] , \inq_ary[14][158] , 
        \inq_ary[14][159] }), .D15({\inq_ary[15][0] , \inq_ary[15][1] , 
        \inq_ary[15][2] , \inq_ary[15][3] , \inq_ary[15][4] , \inq_ary[15][5] , 
        \inq_ary[15][6] , \inq_ary[15][7] , \inq_ary[15][8] , \inq_ary[15][9] , 
        \inq_ary[15][10] , \inq_ary[15][11] , \inq_ary[15][12] , 
        \inq_ary[15][13] , \inq_ary[15][14] , \inq_ary[15][15] , 
        \inq_ary[15][16] , \inq_ary[15][17] , \inq_ary[15][18] , 
        \inq_ary[15][19] , \inq_ary[15][20] , \inq_ary[15][21] , 
        \inq_ary[15][22] , \inq_ary[15][23] , \inq_ary[15][24] , 
        \inq_ary[15][25] , \inq_ary[15][26] , \inq_ary[15][27] , 
        \inq_ary[15][28] , \inq_ary[15][29] , \inq_ary[15][30] , 
        \inq_ary[15][31] , \inq_ary[15][32] , \inq_ary[15][33] , 
        \inq_ary[15][34] , \inq_ary[15][35] , \inq_ary[15][36] , 
        \inq_ary[15][37] , \inq_ary[15][38] , \inq_ary[15][39] , 
        \inq_ary[15][40] , \inq_ary[15][41] , \inq_ary[15][42] , 
        \inq_ary[15][43] , \inq_ary[15][44] , \inq_ary[15][45] , 
        \inq_ary[15][46] , \inq_ary[15][47] , \inq_ary[15][48] , 
        \inq_ary[15][49] , \inq_ary[15][50] , \inq_ary[15][51] , 
        \inq_ary[15][52] , \inq_ary[15][53] , \inq_ary[15][54] , 
        \inq_ary[15][55] , \inq_ary[15][56] , \inq_ary[15][57] , 
        \inq_ary[15][58] , \inq_ary[15][59] , \inq_ary[15][60] , 
        \inq_ary[15][61] , \inq_ary[15][62] , \inq_ary[15][63] , 
        \inq_ary[15][64] , \inq_ary[15][65] , \inq_ary[15][66] , 
        \inq_ary[15][67] , \inq_ary[15][68] , \inq_ary[15][69] , 
        \inq_ary[15][70] , \inq_ary[15][71] , \inq_ary[15][72] , 
        \inq_ary[15][73] , \inq_ary[15][74] , \inq_ary[15][75] , 
        \inq_ary[15][76] , \inq_ary[15][77] , \inq_ary[15][78] , 
        \inq_ary[15][79] , \inq_ary[15][80] , \inq_ary[15][81] , 
        \inq_ary[15][82] , \inq_ary[15][83] , \inq_ary[15][84] , 
        \inq_ary[15][85] , \inq_ary[15][86] , \inq_ary[15][87] , 
        \inq_ary[15][88] , \inq_ary[15][89] , \inq_ary[15][90] , 
        \inq_ary[15][91] , \inq_ary[15][92] , \inq_ary[15][93] , 
        \inq_ary[15][94] , \inq_ary[15][95] , \inq_ary[15][96] , 
        \inq_ary[15][97] , \inq_ary[15][98] , \inq_ary[15][99] , 
        \inq_ary[15][100] , \inq_ary[15][101] , \inq_ary[15][102] , 
        \inq_ary[15][103] , \inq_ary[15][104] , \inq_ary[15][105] , 
        \inq_ary[15][106] , \inq_ary[15][107] , \inq_ary[15][108] , 
        \inq_ary[15][109] , \inq_ary[15][110] , \inq_ary[15][111] , 
        \inq_ary[15][112] , \inq_ary[15][113] , \inq_ary[15][114] , 
        \inq_ary[15][115] , \inq_ary[15][116] , \inq_ary[15][117] , 
        \inq_ary[15][118] , \inq_ary[15][119] , \inq_ary[15][120] , 
        \inq_ary[15][121] , \inq_ary[15][122] , \inq_ary[15][123] , 
        \inq_ary[15][124] , \inq_ary[15][125] , \inq_ary[15][126] , 
        \inq_ary[15][127] , \inq_ary[15][128] , \inq_ary[15][129] , 
        \inq_ary[15][130] , \inq_ary[15][131] , \inq_ary[15][132] , 
        \inq_ary[15][133] , \inq_ary[15][134] , \inq_ary[15][135] , 
        \inq_ary[15][136] , \inq_ary[15][137] , \inq_ary[15][138] , 
        \inq_ary[15][139] , \inq_ary[15][140] , \inq_ary[15][141] , 
        \inq_ary[15][142] , \inq_ary[15][143] , \inq_ary[15][144] , 
        \inq_ary[15][145] , \inq_ary[15][146] , \inq_ary[15][147] , 
        \inq_ary[15][148] , \inq_ary[15][149] , \inq_ary[15][150] , 
        \inq_ary[15][151] , \inq_ary[15][152] , \inq_ary[15][153] , 
        \inq_ary[15][154] , \inq_ary[15][155] , \inq_ary[15][156] , 
        \inq_ary[15][157] , \inq_ary[15][158] , \inq_ary[15][159] }), .S0(N91), 
        .S1(N92), .S2(N93), .S3(N94), .Z({N258, N257, N256, N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 
        N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, 
        N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, 
        N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, 
        N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, 
        N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, 
        N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99}) );
  GTECH_BUF B_83 ( .A(rdptr_d1[0]), .Z(N91) );
  GTECH_BUF B_84 ( .A(rdptr_d1[1]), .Z(N92) );
  GTECH_BUF B_85 ( .A(rdptr_d1[2]), .Z(N93) );
  GTECH_BUF B_86 ( .A(rdptr_d1[3]), .Z(N94) );
  MUX_OP C25071 ( .D0({\inq_ary[0][0] , \inq_ary[0][1] , \inq_ary[0][2] , 
        \inq_ary[0][3] , \inq_ary[0][4] , \inq_ary[0][5] , \inq_ary[0][6] , 
        \inq_ary[0][7] , \inq_ary[0][8] , \inq_ary[0][9] , \inq_ary[0][10] , 
        \inq_ary[0][11] , \inq_ary[0][12] , \inq_ary[0][13] , \inq_ary[0][14] , 
        \inq_ary[0][15] , \inq_ary[0][16] , \inq_ary[0][17] , \inq_ary[0][18] , 
        \inq_ary[0][19] , \inq_ary[0][20] , \inq_ary[0][21] , \inq_ary[0][22] , 
        \inq_ary[0][23] , \inq_ary[0][24] , \inq_ary[0][25] , \inq_ary[0][26] , 
        \inq_ary[0][27] , \inq_ary[0][28] , \inq_ary[0][29] , \inq_ary[0][30] , 
        \inq_ary[0][31] , \inq_ary[0][32] , \inq_ary[0][33] , \inq_ary[0][34] , 
        \inq_ary[0][35] , \inq_ary[0][36] , \inq_ary[0][37] , \inq_ary[0][38] , 
        \inq_ary[0][39] , \inq_ary[0][40] , \inq_ary[0][41] , \inq_ary[0][42] , 
        \inq_ary[0][43] , \inq_ary[0][44] , \inq_ary[0][45] , \inq_ary[0][46] , 
        \inq_ary[0][47] , \inq_ary[0][48] , \inq_ary[0][49] , \inq_ary[0][50] , 
        \inq_ary[0][51] , \inq_ary[0][52] , \inq_ary[0][53] , \inq_ary[0][54] , 
        \inq_ary[0][55] , \inq_ary[0][56] , \inq_ary[0][57] , \inq_ary[0][58] , 
        \inq_ary[0][59] , \inq_ary[0][60] , \inq_ary[0][61] , \inq_ary[0][62] , 
        \inq_ary[0][63] , \inq_ary[0][64] , \inq_ary[0][65] , \inq_ary[0][66] , 
        \inq_ary[0][67] , \inq_ary[0][68] , \inq_ary[0][69] , \inq_ary[0][70] , 
        \inq_ary[0][71] , \inq_ary[0][72] , \inq_ary[0][73] , \inq_ary[0][74] , 
        \inq_ary[0][75] , \inq_ary[0][76] , \inq_ary[0][77] , \inq_ary[0][78] , 
        \inq_ary[0][79] , \inq_ary[0][80] , \inq_ary[0][81] , \inq_ary[0][82] , 
        \inq_ary[0][83] , \inq_ary[0][84] , \inq_ary[0][85] , \inq_ary[0][86] , 
        \inq_ary[0][87] , \inq_ary[0][88] , \inq_ary[0][89] , \inq_ary[0][90] , 
        \inq_ary[0][91] , \inq_ary[0][92] , \inq_ary[0][93] , \inq_ary[0][94] , 
        \inq_ary[0][95] , \inq_ary[0][96] , \inq_ary[0][97] , \inq_ary[0][98] , 
        \inq_ary[0][99] , \inq_ary[0][100] , \inq_ary[0][101] , 
        \inq_ary[0][102] , \inq_ary[0][103] , \inq_ary[0][104] , 
        \inq_ary[0][105] , \inq_ary[0][106] , \inq_ary[0][107] , 
        \inq_ary[0][108] , \inq_ary[0][109] , \inq_ary[0][110] , 
        \inq_ary[0][111] , \inq_ary[0][112] , \inq_ary[0][113] , 
        \inq_ary[0][114] , \inq_ary[0][115] , \inq_ary[0][116] , 
        \inq_ary[0][117] , \inq_ary[0][118] , \inq_ary[0][119] , 
        \inq_ary[0][120] , \inq_ary[0][121] , \inq_ary[0][122] , 
        \inq_ary[0][123] , \inq_ary[0][124] , \inq_ary[0][125] , 
        \inq_ary[0][126] , \inq_ary[0][127] , \inq_ary[0][128] , 
        \inq_ary[0][129] , \inq_ary[0][130] , \inq_ary[0][131] , 
        \inq_ary[0][132] , \inq_ary[0][133] , \inq_ary[0][134] , 
        \inq_ary[0][135] , \inq_ary[0][136] , \inq_ary[0][137] , 
        \inq_ary[0][138] , \inq_ary[0][139] , \inq_ary[0][140] , 
        \inq_ary[0][141] , \inq_ary[0][142] , \inq_ary[0][143] , 
        \inq_ary[0][144] , \inq_ary[0][145] , \inq_ary[0][146] , 
        \inq_ary[0][147] , \inq_ary[0][148] , \inq_ary[0][149] , 
        \inq_ary[0][150] , \inq_ary[0][151] , \inq_ary[0][152] , 
        \inq_ary[0][153] , \inq_ary[0][154] , \inq_ary[0][155] , 
        \inq_ary[0][156] , \inq_ary[0][157] , \inq_ary[0][158] , 
        \inq_ary[0][159] }), .D1({\inq_ary[1][0] , \inq_ary[1][1] , 
        \inq_ary[1][2] , \inq_ary[1][3] , \inq_ary[1][4] , \inq_ary[1][5] , 
        \inq_ary[1][6] , \inq_ary[1][7] , \inq_ary[1][8] , \inq_ary[1][9] , 
        \inq_ary[1][10] , \inq_ary[1][11] , \inq_ary[1][12] , \inq_ary[1][13] , 
        \inq_ary[1][14] , \inq_ary[1][15] , \inq_ary[1][16] , \inq_ary[1][17] , 
        \inq_ary[1][18] , \inq_ary[1][19] , \inq_ary[1][20] , \inq_ary[1][21] , 
        \inq_ary[1][22] , \inq_ary[1][23] , \inq_ary[1][24] , \inq_ary[1][25] , 
        \inq_ary[1][26] , \inq_ary[1][27] , \inq_ary[1][28] , \inq_ary[1][29] , 
        \inq_ary[1][30] , \inq_ary[1][31] , \inq_ary[1][32] , \inq_ary[1][33] , 
        \inq_ary[1][34] , \inq_ary[1][35] , \inq_ary[1][36] , \inq_ary[1][37] , 
        \inq_ary[1][38] , \inq_ary[1][39] , \inq_ary[1][40] , \inq_ary[1][41] , 
        \inq_ary[1][42] , \inq_ary[1][43] , \inq_ary[1][44] , \inq_ary[1][45] , 
        \inq_ary[1][46] , \inq_ary[1][47] , \inq_ary[1][48] , \inq_ary[1][49] , 
        \inq_ary[1][50] , \inq_ary[1][51] , \inq_ary[1][52] , \inq_ary[1][53] , 
        \inq_ary[1][54] , \inq_ary[1][55] , \inq_ary[1][56] , \inq_ary[1][57] , 
        \inq_ary[1][58] , \inq_ary[1][59] , \inq_ary[1][60] , \inq_ary[1][61] , 
        \inq_ary[1][62] , \inq_ary[1][63] , \inq_ary[1][64] , \inq_ary[1][65] , 
        \inq_ary[1][66] , \inq_ary[1][67] , \inq_ary[1][68] , \inq_ary[1][69] , 
        \inq_ary[1][70] , \inq_ary[1][71] , \inq_ary[1][72] , \inq_ary[1][73] , 
        \inq_ary[1][74] , \inq_ary[1][75] , \inq_ary[1][76] , \inq_ary[1][77] , 
        \inq_ary[1][78] , \inq_ary[1][79] , \inq_ary[1][80] , \inq_ary[1][81] , 
        \inq_ary[1][82] , \inq_ary[1][83] , \inq_ary[1][84] , \inq_ary[1][85] , 
        \inq_ary[1][86] , \inq_ary[1][87] , \inq_ary[1][88] , \inq_ary[1][89] , 
        \inq_ary[1][90] , \inq_ary[1][91] , \inq_ary[1][92] , \inq_ary[1][93] , 
        \inq_ary[1][94] , \inq_ary[1][95] , \inq_ary[1][96] , \inq_ary[1][97] , 
        \inq_ary[1][98] , \inq_ary[1][99] , \inq_ary[1][100] , 
        \inq_ary[1][101] , \inq_ary[1][102] , \inq_ary[1][103] , 
        \inq_ary[1][104] , \inq_ary[1][105] , \inq_ary[1][106] , 
        \inq_ary[1][107] , \inq_ary[1][108] , \inq_ary[1][109] , 
        \inq_ary[1][110] , \inq_ary[1][111] , \inq_ary[1][112] , 
        \inq_ary[1][113] , \inq_ary[1][114] , \inq_ary[1][115] , 
        \inq_ary[1][116] , \inq_ary[1][117] , \inq_ary[1][118] , 
        \inq_ary[1][119] , \inq_ary[1][120] , \inq_ary[1][121] , 
        \inq_ary[1][122] , \inq_ary[1][123] , \inq_ary[1][124] , 
        \inq_ary[1][125] , \inq_ary[1][126] , \inq_ary[1][127] , 
        \inq_ary[1][128] , \inq_ary[1][129] , \inq_ary[1][130] , 
        \inq_ary[1][131] , \inq_ary[1][132] , \inq_ary[1][133] , 
        \inq_ary[1][134] , \inq_ary[1][135] , \inq_ary[1][136] , 
        \inq_ary[1][137] , \inq_ary[1][138] , \inq_ary[1][139] , 
        \inq_ary[1][140] , \inq_ary[1][141] , \inq_ary[1][142] , 
        \inq_ary[1][143] , \inq_ary[1][144] , \inq_ary[1][145] , 
        \inq_ary[1][146] , \inq_ary[1][147] , \inq_ary[1][148] , 
        \inq_ary[1][149] , \inq_ary[1][150] , \inq_ary[1][151] , 
        \inq_ary[1][152] , \inq_ary[1][153] , \inq_ary[1][154] , 
        \inq_ary[1][155] , \inq_ary[1][156] , \inq_ary[1][157] , 
        \inq_ary[1][158] , \inq_ary[1][159] }), .D2({\inq_ary[2][0] , 
        \inq_ary[2][1] , \inq_ary[2][2] , \inq_ary[2][3] , \inq_ary[2][4] , 
        \inq_ary[2][5] , \inq_ary[2][6] , \inq_ary[2][7] , \inq_ary[2][8] , 
        \inq_ary[2][9] , \inq_ary[2][10] , \inq_ary[2][11] , \inq_ary[2][12] , 
        \inq_ary[2][13] , \inq_ary[2][14] , \inq_ary[2][15] , \inq_ary[2][16] , 
        \inq_ary[2][17] , \inq_ary[2][18] , \inq_ary[2][19] , \inq_ary[2][20] , 
        \inq_ary[2][21] , \inq_ary[2][22] , \inq_ary[2][23] , \inq_ary[2][24] , 
        \inq_ary[2][25] , \inq_ary[2][26] , \inq_ary[2][27] , \inq_ary[2][28] , 
        \inq_ary[2][29] , \inq_ary[2][30] , \inq_ary[2][31] , \inq_ary[2][32] , 
        \inq_ary[2][33] , \inq_ary[2][34] , \inq_ary[2][35] , \inq_ary[2][36] , 
        \inq_ary[2][37] , \inq_ary[2][38] , \inq_ary[2][39] , \inq_ary[2][40] , 
        \inq_ary[2][41] , \inq_ary[2][42] , \inq_ary[2][43] , \inq_ary[2][44] , 
        \inq_ary[2][45] , \inq_ary[2][46] , \inq_ary[2][47] , \inq_ary[2][48] , 
        \inq_ary[2][49] , \inq_ary[2][50] , \inq_ary[2][51] , \inq_ary[2][52] , 
        \inq_ary[2][53] , \inq_ary[2][54] , \inq_ary[2][55] , \inq_ary[2][56] , 
        \inq_ary[2][57] , \inq_ary[2][58] , \inq_ary[2][59] , \inq_ary[2][60] , 
        \inq_ary[2][61] , \inq_ary[2][62] , \inq_ary[2][63] , \inq_ary[2][64] , 
        \inq_ary[2][65] , \inq_ary[2][66] , \inq_ary[2][67] , \inq_ary[2][68] , 
        \inq_ary[2][69] , \inq_ary[2][70] , \inq_ary[2][71] , \inq_ary[2][72] , 
        \inq_ary[2][73] , \inq_ary[2][74] , \inq_ary[2][75] , \inq_ary[2][76] , 
        \inq_ary[2][77] , \inq_ary[2][78] , \inq_ary[2][79] , \inq_ary[2][80] , 
        \inq_ary[2][81] , \inq_ary[2][82] , \inq_ary[2][83] , \inq_ary[2][84] , 
        \inq_ary[2][85] , \inq_ary[2][86] , \inq_ary[2][87] , \inq_ary[2][88] , 
        \inq_ary[2][89] , \inq_ary[2][90] , \inq_ary[2][91] , \inq_ary[2][92] , 
        \inq_ary[2][93] , \inq_ary[2][94] , \inq_ary[2][95] , \inq_ary[2][96] , 
        \inq_ary[2][97] , \inq_ary[2][98] , \inq_ary[2][99] , 
        \inq_ary[2][100] , \inq_ary[2][101] , \inq_ary[2][102] , 
        \inq_ary[2][103] , \inq_ary[2][104] , \inq_ary[2][105] , 
        \inq_ary[2][106] , \inq_ary[2][107] , \inq_ary[2][108] , 
        \inq_ary[2][109] , \inq_ary[2][110] , \inq_ary[2][111] , 
        \inq_ary[2][112] , \inq_ary[2][113] , \inq_ary[2][114] , 
        \inq_ary[2][115] , \inq_ary[2][116] , \inq_ary[2][117] , 
        \inq_ary[2][118] , \inq_ary[2][119] , \inq_ary[2][120] , 
        \inq_ary[2][121] , \inq_ary[2][122] , \inq_ary[2][123] , 
        \inq_ary[2][124] , \inq_ary[2][125] , \inq_ary[2][126] , 
        \inq_ary[2][127] , \inq_ary[2][128] , \inq_ary[2][129] , 
        \inq_ary[2][130] , \inq_ary[2][131] , \inq_ary[2][132] , 
        \inq_ary[2][133] , \inq_ary[2][134] , \inq_ary[2][135] , 
        \inq_ary[2][136] , \inq_ary[2][137] , \inq_ary[2][138] , 
        \inq_ary[2][139] , \inq_ary[2][140] , \inq_ary[2][141] , 
        \inq_ary[2][142] , \inq_ary[2][143] , \inq_ary[2][144] , 
        \inq_ary[2][145] , \inq_ary[2][146] , \inq_ary[2][147] , 
        \inq_ary[2][148] , \inq_ary[2][149] , \inq_ary[2][150] , 
        \inq_ary[2][151] , \inq_ary[2][152] , \inq_ary[2][153] , 
        \inq_ary[2][154] , \inq_ary[2][155] , \inq_ary[2][156] , 
        \inq_ary[2][157] , \inq_ary[2][158] , \inq_ary[2][159] }), .D3({
        \inq_ary[3][0] , \inq_ary[3][1] , \inq_ary[3][2] , \inq_ary[3][3] , 
        \inq_ary[3][4] , \inq_ary[3][5] , \inq_ary[3][6] , \inq_ary[3][7] , 
        \inq_ary[3][8] , \inq_ary[3][9] , \inq_ary[3][10] , \inq_ary[3][11] , 
        \inq_ary[3][12] , \inq_ary[3][13] , \inq_ary[3][14] , \inq_ary[3][15] , 
        \inq_ary[3][16] , \inq_ary[3][17] , \inq_ary[3][18] , \inq_ary[3][19] , 
        \inq_ary[3][20] , \inq_ary[3][21] , \inq_ary[3][22] , \inq_ary[3][23] , 
        \inq_ary[3][24] , \inq_ary[3][25] , \inq_ary[3][26] , \inq_ary[3][27] , 
        \inq_ary[3][28] , \inq_ary[3][29] , \inq_ary[3][30] , \inq_ary[3][31] , 
        \inq_ary[3][32] , \inq_ary[3][33] , \inq_ary[3][34] , \inq_ary[3][35] , 
        \inq_ary[3][36] , \inq_ary[3][37] , \inq_ary[3][38] , \inq_ary[3][39] , 
        \inq_ary[3][40] , \inq_ary[3][41] , \inq_ary[3][42] , \inq_ary[3][43] , 
        \inq_ary[3][44] , \inq_ary[3][45] , \inq_ary[3][46] , \inq_ary[3][47] , 
        \inq_ary[3][48] , \inq_ary[3][49] , \inq_ary[3][50] , \inq_ary[3][51] , 
        \inq_ary[3][52] , \inq_ary[3][53] , \inq_ary[3][54] , \inq_ary[3][55] , 
        \inq_ary[3][56] , \inq_ary[3][57] , \inq_ary[3][58] , \inq_ary[3][59] , 
        \inq_ary[3][60] , \inq_ary[3][61] , \inq_ary[3][62] , \inq_ary[3][63] , 
        \inq_ary[3][64] , \inq_ary[3][65] , \inq_ary[3][66] , \inq_ary[3][67] , 
        \inq_ary[3][68] , \inq_ary[3][69] , \inq_ary[3][70] , \inq_ary[3][71] , 
        \inq_ary[3][72] , \inq_ary[3][73] , \inq_ary[3][74] , \inq_ary[3][75] , 
        \inq_ary[3][76] , \inq_ary[3][77] , \inq_ary[3][78] , \inq_ary[3][79] , 
        \inq_ary[3][80] , \inq_ary[3][81] , \inq_ary[3][82] , \inq_ary[3][83] , 
        \inq_ary[3][84] , \inq_ary[3][85] , \inq_ary[3][86] , \inq_ary[3][87] , 
        \inq_ary[3][88] , \inq_ary[3][89] , \inq_ary[3][90] , \inq_ary[3][91] , 
        \inq_ary[3][92] , \inq_ary[3][93] , \inq_ary[3][94] , \inq_ary[3][95] , 
        \inq_ary[3][96] , \inq_ary[3][97] , \inq_ary[3][98] , \inq_ary[3][99] , 
        \inq_ary[3][100] , \inq_ary[3][101] , \inq_ary[3][102] , 
        \inq_ary[3][103] , \inq_ary[3][104] , \inq_ary[3][105] , 
        \inq_ary[3][106] , \inq_ary[3][107] , \inq_ary[3][108] , 
        \inq_ary[3][109] , \inq_ary[3][110] , \inq_ary[3][111] , 
        \inq_ary[3][112] , \inq_ary[3][113] , \inq_ary[3][114] , 
        \inq_ary[3][115] , \inq_ary[3][116] , \inq_ary[3][117] , 
        \inq_ary[3][118] , \inq_ary[3][119] , \inq_ary[3][120] , 
        \inq_ary[3][121] , \inq_ary[3][122] , \inq_ary[3][123] , 
        \inq_ary[3][124] , \inq_ary[3][125] , \inq_ary[3][126] , 
        \inq_ary[3][127] , \inq_ary[3][128] , \inq_ary[3][129] , 
        \inq_ary[3][130] , \inq_ary[3][131] , \inq_ary[3][132] , 
        \inq_ary[3][133] , \inq_ary[3][134] , \inq_ary[3][135] , 
        \inq_ary[3][136] , \inq_ary[3][137] , \inq_ary[3][138] , 
        \inq_ary[3][139] , \inq_ary[3][140] , \inq_ary[3][141] , 
        \inq_ary[3][142] , \inq_ary[3][143] , \inq_ary[3][144] , 
        \inq_ary[3][145] , \inq_ary[3][146] , \inq_ary[3][147] , 
        \inq_ary[3][148] , \inq_ary[3][149] , \inq_ary[3][150] , 
        \inq_ary[3][151] , \inq_ary[3][152] , \inq_ary[3][153] , 
        \inq_ary[3][154] , \inq_ary[3][155] , \inq_ary[3][156] , 
        \inq_ary[3][157] , \inq_ary[3][158] , \inq_ary[3][159] }), .D4({
        \inq_ary[4][0] , \inq_ary[4][1] , \inq_ary[4][2] , \inq_ary[4][3] , 
        \inq_ary[4][4] , \inq_ary[4][5] , \inq_ary[4][6] , \inq_ary[4][7] , 
        \inq_ary[4][8] , \inq_ary[4][9] , \inq_ary[4][10] , \inq_ary[4][11] , 
        \inq_ary[4][12] , \inq_ary[4][13] , \inq_ary[4][14] , \inq_ary[4][15] , 
        \inq_ary[4][16] , \inq_ary[4][17] , \inq_ary[4][18] , \inq_ary[4][19] , 
        \inq_ary[4][20] , \inq_ary[4][21] , \inq_ary[4][22] , \inq_ary[4][23] , 
        \inq_ary[4][24] , \inq_ary[4][25] , \inq_ary[4][26] , \inq_ary[4][27] , 
        \inq_ary[4][28] , \inq_ary[4][29] , \inq_ary[4][30] , \inq_ary[4][31] , 
        \inq_ary[4][32] , \inq_ary[4][33] , \inq_ary[4][34] , \inq_ary[4][35] , 
        \inq_ary[4][36] , \inq_ary[4][37] , \inq_ary[4][38] , \inq_ary[4][39] , 
        \inq_ary[4][40] , \inq_ary[4][41] , \inq_ary[4][42] , \inq_ary[4][43] , 
        \inq_ary[4][44] , \inq_ary[4][45] , \inq_ary[4][46] , \inq_ary[4][47] , 
        \inq_ary[4][48] , \inq_ary[4][49] , \inq_ary[4][50] , \inq_ary[4][51] , 
        \inq_ary[4][52] , \inq_ary[4][53] , \inq_ary[4][54] , \inq_ary[4][55] , 
        \inq_ary[4][56] , \inq_ary[4][57] , \inq_ary[4][58] , \inq_ary[4][59] , 
        \inq_ary[4][60] , \inq_ary[4][61] , \inq_ary[4][62] , \inq_ary[4][63] , 
        \inq_ary[4][64] , \inq_ary[4][65] , \inq_ary[4][66] , \inq_ary[4][67] , 
        \inq_ary[4][68] , \inq_ary[4][69] , \inq_ary[4][70] , \inq_ary[4][71] , 
        \inq_ary[4][72] , \inq_ary[4][73] , \inq_ary[4][74] , \inq_ary[4][75] , 
        \inq_ary[4][76] , \inq_ary[4][77] , \inq_ary[4][78] , \inq_ary[4][79] , 
        \inq_ary[4][80] , \inq_ary[4][81] , \inq_ary[4][82] , \inq_ary[4][83] , 
        \inq_ary[4][84] , \inq_ary[4][85] , \inq_ary[4][86] , \inq_ary[4][87] , 
        \inq_ary[4][88] , \inq_ary[4][89] , \inq_ary[4][90] , \inq_ary[4][91] , 
        \inq_ary[4][92] , \inq_ary[4][93] , \inq_ary[4][94] , \inq_ary[4][95] , 
        \inq_ary[4][96] , \inq_ary[4][97] , \inq_ary[4][98] , \inq_ary[4][99] , 
        \inq_ary[4][100] , \inq_ary[4][101] , \inq_ary[4][102] , 
        \inq_ary[4][103] , \inq_ary[4][104] , \inq_ary[4][105] , 
        \inq_ary[4][106] , \inq_ary[4][107] , \inq_ary[4][108] , 
        \inq_ary[4][109] , \inq_ary[4][110] , \inq_ary[4][111] , 
        \inq_ary[4][112] , \inq_ary[4][113] , \inq_ary[4][114] , 
        \inq_ary[4][115] , \inq_ary[4][116] , \inq_ary[4][117] , 
        \inq_ary[4][118] , \inq_ary[4][119] , \inq_ary[4][120] , 
        \inq_ary[4][121] , \inq_ary[4][122] , \inq_ary[4][123] , 
        \inq_ary[4][124] , \inq_ary[4][125] , \inq_ary[4][126] , 
        \inq_ary[4][127] , \inq_ary[4][128] , \inq_ary[4][129] , 
        \inq_ary[4][130] , \inq_ary[4][131] , \inq_ary[4][132] , 
        \inq_ary[4][133] , \inq_ary[4][134] , \inq_ary[4][135] , 
        \inq_ary[4][136] , \inq_ary[4][137] , \inq_ary[4][138] , 
        \inq_ary[4][139] , \inq_ary[4][140] , \inq_ary[4][141] , 
        \inq_ary[4][142] , \inq_ary[4][143] , \inq_ary[4][144] , 
        \inq_ary[4][145] , \inq_ary[4][146] , \inq_ary[4][147] , 
        \inq_ary[4][148] , \inq_ary[4][149] , \inq_ary[4][150] , 
        \inq_ary[4][151] , \inq_ary[4][152] , \inq_ary[4][153] , 
        \inq_ary[4][154] , \inq_ary[4][155] , \inq_ary[4][156] , 
        \inq_ary[4][157] , \inq_ary[4][158] , \inq_ary[4][159] }), .D5({
        \inq_ary[5][0] , \inq_ary[5][1] , \inq_ary[5][2] , \inq_ary[5][3] , 
        \inq_ary[5][4] , \inq_ary[5][5] , \inq_ary[5][6] , \inq_ary[5][7] , 
        \inq_ary[5][8] , \inq_ary[5][9] , \inq_ary[5][10] , \inq_ary[5][11] , 
        \inq_ary[5][12] , \inq_ary[5][13] , \inq_ary[5][14] , \inq_ary[5][15] , 
        \inq_ary[5][16] , \inq_ary[5][17] , \inq_ary[5][18] , \inq_ary[5][19] , 
        \inq_ary[5][20] , \inq_ary[5][21] , \inq_ary[5][22] , \inq_ary[5][23] , 
        \inq_ary[5][24] , \inq_ary[5][25] , \inq_ary[5][26] , \inq_ary[5][27] , 
        \inq_ary[5][28] , \inq_ary[5][29] , \inq_ary[5][30] , \inq_ary[5][31] , 
        \inq_ary[5][32] , \inq_ary[5][33] , \inq_ary[5][34] , \inq_ary[5][35] , 
        \inq_ary[5][36] , \inq_ary[5][37] , \inq_ary[5][38] , \inq_ary[5][39] , 
        \inq_ary[5][40] , \inq_ary[5][41] , \inq_ary[5][42] , \inq_ary[5][43] , 
        \inq_ary[5][44] , \inq_ary[5][45] , \inq_ary[5][46] , \inq_ary[5][47] , 
        \inq_ary[5][48] , \inq_ary[5][49] , \inq_ary[5][50] , \inq_ary[5][51] , 
        \inq_ary[5][52] , \inq_ary[5][53] , \inq_ary[5][54] , \inq_ary[5][55] , 
        \inq_ary[5][56] , \inq_ary[5][57] , \inq_ary[5][58] , \inq_ary[5][59] , 
        \inq_ary[5][60] , \inq_ary[5][61] , \inq_ary[5][62] , \inq_ary[5][63] , 
        \inq_ary[5][64] , \inq_ary[5][65] , \inq_ary[5][66] , \inq_ary[5][67] , 
        \inq_ary[5][68] , \inq_ary[5][69] , \inq_ary[5][70] , \inq_ary[5][71] , 
        \inq_ary[5][72] , \inq_ary[5][73] , \inq_ary[5][74] , \inq_ary[5][75] , 
        \inq_ary[5][76] , \inq_ary[5][77] , \inq_ary[5][78] , \inq_ary[5][79] , 
        \inq_ary[5][80] , \inq_ary[5][81] , \inq_ary[5][82] , \inq_ary[5][83] , 
        \inq_ary[5][84] , \inq_ary[5][85] , \inq_ary[5][86] , \inq_ary[5][87] , 
        \inq_ary[5][88] , \inq_ary[5][89] , \inq_ary[5][90] , \inq_ary[5][91] , 
        \inq_ary[5][92] , \inq_ary[5][93] , \inq_ary[5][94] , \inq_ary[5][95] , 
        \inq_ary[5][96] , \inq_ary[5][97] , \inq_ary[5][98] , \inq_ary[5][99] , 
        \inq_ary[5][100] , \inq_ary[5][101] , \inq_ary[5][102] , 
        \inq_ary[5][103] , \inq_ary[5][104] , \inq_ary[5][105] , 
        \inq_ary[5][106] , \inq_ary[5][107] , \inq_ary[5][108] , 
        \inq_ary[5][109] , \inq_ary[5][110] , \inq_ary[5][111] , 
        \inq_ary[5][112] , \inq_ary[5][113] , \inq_ary[5][114] , 
        \inq_ary[5][115] , \inq_ary[5][116] , \inq_ary[5][117] , 
        \inq_ary[5][118] , \inq_ary[5][119] , \inq_ary[5][120] , 
        \inq_ary[5][121] , \inq_ary[5][122] , \inq_ary[5][123] , 
        \inq_ary[5][124] , \inq_ary[5][125] , \inq_ary[5][126] , 
        \inq_ary[5][127] , \inq_ary[5][128] , \inq_ary[5][129] , 
        \inq_ary[5][130] , \inq_ary[5][131] , \inq_ary[5][132] , 
        \inq_ary[5][133] , \inq_ary[5][134] , \inq_ary[5][135] , 
        \inq_ary[5][136] , \inq_ary[5][137] , \inq_ary[5][138] , 
        \inq_ary[5][139] , \inq_ary[5][140] , \inq_ary[5][141] , 
        \inq_ary[5][142] , \inq_ary[5][143] , \inq_ary[5][144] , 
        \inq_ary[5][145] , \inq_ary[5][146] , \inq_ary[5][147] , 
        \inq_ary[5][148] , \inq_ary[5][149] , \inq_ary[5][150] , 
        \inq_ary[5][151] , \inq_ary[5][152] , \inq_ary[5][153] , 
        \inq_ary[5][154] , \inq_ary[5][155] , \inq_ary[5][156] , 
        \inq_ary[5][157] , \inq_ary[5][158] , \inq_ary[5][159] }), .D6({
        \inq_ary[6][0] , \inq_ary[6][1] , \inq_ary[6][2] , \inq_ary[6][3] , 
        \inq_ary[6][4] , \inq_ary[6][5] , \inq_ary[6][6] , \inq_ary[6][7] , 
        \inq_ary[6][8] , \inq_ary[6][9] , \inq_ary[6][10] , \inq_ary[6][11] , 
        \inq_ary[6][12] , \inq_ary[6][13] , \inq_ary[6][14] , \inq_ary[6][15] , 
        \inq_ary[6][16] , \inq_ary[6][17] , \inq_ary[6][18] , \inq_ary[6][19] , 
        \inq_ary[6][20] , \inq_ary[6][21] , \inq_ary[6][22] , \inq_ary[6][23] , 
        \inq_ary[6][24] , \inq_ary[6][25] , \inq_ary[6][26] , \inq_ary[6][27] , 
        \inq_ary[6][28] , \inq_ary[6][29] , \inq_ary[6][30] , \inq_ary[6][31] , 
        \inq_ary[6][32] , \inq_ary[6][33] , \inq_ary[6][34] , \inq_ary[6][35] , 
        \inq_ary[6][36] , \inq_ary[6][37] , \inq_ary[6][38] , \inq_ary[6][39] , 
        \inq_ary[6][40] , \inq_ary[6][41] , \inq_ary[6][42] , \inq_ary[6][43] , 
        \inq_ary[6][44] , \inq_ary[6][45] , \inq_ary[6][46] , \inq_ary[6][47] , 
        \inq_ary[6][48] , \inq_ary[6][49] , \inq_ary[6][50] , \inq_ary[6][51] , 
        \inq_ary[6][52] , \inq_ary[6][53] , \inq_ary[6][54] , \inq_ary[6][55] , 
        \inq_ary[6][56] , \inq_ary[6][57] , \inq_ary[6][58] , \inq_ary[6][59] , 
        \inq_ary[6][60] , \inq_ary[6][61] , \inq_ary[6][62] , \inq_ary[6][63] , 
        \inq_ary[6][64] , \inq_ary[6][65] , \inq_ary[6][66] , \inq_ary[6][67] , 
        \inq_ary[6][68] , \inq_ary[6][69] , \inq_ary[6][70] , \inq_ary[6][71] , 
        \inq_ary[6][72] , \inq_ary[6][73] , \inq_ary[6][74] , \inq_ary[6][75] , 
        \inq_ary[6][76] , \inq_ary[6][77] , \inq_ary[6][78] , \inq_ary[6][79] , 
        \inq_ary[6][80] , \inq_ary[6][81] , \inq_ary[6][82] , \inq_ary[6][83] , 
        \inq_ary[6][84] , \inq_ary[6][85] , \inq_ary[6][86] , \inq_ary[6][87] , 
        \inq_ary[6][88] , \inq_ary[6][89] , \inq_ary[6][90] , \inq_ary[6][91] , 
        \inq_ary[6][92] , \inq_ary[6][93] , \inq_ary[6][94] , \inq_ary[6][95] , 
        \inq_ary[6][96] , \inq_ary[6][97] , \inq_ary[6][98] , \inq_ary[6][99] , 
        \inq_ary[6][100] , \inq_ary[6][101] , \inq_ary[6][102] , 
        \inq_ary[6][103] , \inq_ary[6][104] , \inq_ary[6][105] , 
        \inq_ary[6][106] , \inq_ary[6][107] , \inq_ary[6][108] , 
        \inq_ary[6][109] , \inq_ary[6][110] , \inq_ary[6][111] , 
        \inq_ary[6][112] , \inq_ary[6][113] , \inq_ary[6][114] , 
        \inq_ary[6][115] , \inq_ary[6][116] , \inq_ary[6][117] , 
        \inq_ary[6][118] , \inq_ary[6][119] , \inq_ary[6][120] , 
        \inq_ary[6][121] , \inq_ary[6][122] , \inq_ary[6][123] , 
        \inq_ary[6][124] , \inq_ary[6][125] , \inq_ary[6][126] , 
        \inq_ary[6][127] , \inq_ary[6][128] , \inq_ary[6][129] , 
        \inq_ary[6][130] , \inq_ary[6][131] , \inq_ary[6][132] , 
        \inq_ary[6][133] , \inq_ary[6][134] , \inq_ary[6][135] , 
        \inq_ary[6][136] , \inq_ary[6][137] , \inq_ary[6][138] , 
        \inq_ary[6][139] , \inq_ary[6][140] , \inq_ary[6][141] , 
        \inq_ary[6][142] , \inq_ary[6][143] , \inq_ary[6][144] , 
        \inq_ary[6][145] , \inq_ary[6][146] , \inq_ary[6][147] , 
        \inq_ary[6][148] , \inq_ary[6][149] , \inq_ary[6][150] , 
        \inq_ary[6][151] , \inq_ary[6][152] , \inq_ary[6][153] , 
        \inq_ary[6][154] , \inq_ary[6][155] , \inq_ary[6][156] , 
        \inq_ary[6][157] , \inq_ary[6][158] , \inq_ary[6][159] }), .D7({
        \inq_ary[7][0] , \inq_ary[7][1] , \inq_ary[7][2] , \inq_ary[7][3] , 
        \inq_ary[7][4] , \inq_ary[7][5] , \inq_ary[7][6] , \inq_ary[7][7] , 
        \inq_ary[7][8] , \inq_ary[7][9] , \inq_ary[7][10] , \inq_ary[7][11] , 
        \inq_ary[7][12] , \inq_ary[7][13] , \inq_ary[7][14] , \inq_ary[7][15] , 
        \inq_ary[7][16] , \inq_ary[7][17] , \inq_ary[7][18] , \inq_ary[7][19] , 
        \inq_ary[7][20] , \inq_ary[7][21] , \inq_ary[7][22] , \inq_ary[7][23] , 
        \inq_ary[7][24] , \inq_ary[7][25] , \inq_ary[7][26] , \inq_ary[7][27] , 
        \inq_ary[7][28] , \inq_ary[7][29] , \inq_ary[7][30] , \inq_ary[7][31] , 
        \inq_ary[7][32] , \inq_ary[7][33] , \inq_ary[7][34] , \inq_ary[7][35] , 
        \inq_ary[7][36] , \inq_ary[7][37] , \inq_ary[7][38] , \inq_ary[7][39] , 
        \inq_ary[7][40] , \inq_ary[7][41] , \inq_ary[7][42] , \inq_ary[7][43] , 
        \inq_ary[7][44] , \inq_ary[7][45] , \inq_ary[7][46] , \inq_ary[7][47] , 
        \inq_ary[7][48] , \inq_ary[7][49] , \inq_ary[7][50] , \inq_ary[7][51] , 
        \inq_ary[7][52] , \inq_ary[7][53] , \inq_ary[7][54] , \inq_ary[7][55] , 
        \inq_ary[7][56] , \inq_ary[7][57] , \inq_ary[7][58] , \inq_ary[7][59] , 
        \inq_ary[7][60] , \inq_ary[7][61] , \inq_ary[7][62] , \inq_ary[7][63] , 
        \inq_ary[7][64] , \inq_ary[7][65] , \inq_ary[7][66] , \inq_ary[7][67] , 
        \inq_ary[7][68] , \inq_ary[7][69] , \inq_ary[7][70] , \inq_ary[7][71] , 
        \inq_ary[7][72] , \inq_ary[7][73] , \inq_ary[7][74] , \inq_ary[7][75] , 
        \inq_ary[7][76] , \inq_ary[7][77] , \inq_ary[7][78] , \inq_ary[7][79] , 
        \inq_ary[7][80] , \inq_ary[7][81] , \inq_ary[7][82] , \inq_ary[7][83] , 
        \inq_ary[7][84] , \inq_ary[7][85] , \inq_ary[7][86] , \inq_ary[7][87] , 
        \inq_ary[7][88] , \inq_ary[7][89] , \inq_ary[7][90] , \inq_ary[7][91] , 
        \inq_ary[7][92] , \inq_ary[7][93] , \inq_ary[7][94] , \inq_ary[7][95] , 
        \inq_ary[7][96] , \inq_ary[7][97] , \inq_ary[7][98] , \inq_ary[7][99] , 
        \inq_ary[7][100] , \inq_ary[7][101] , \inq_ary[7][102] , 
        \inq_ary[7][103] , \inq_ary[7][104] , \inq_ary[7][105] , 
        \inq_ary[7][106] , \inq_ary[7][107] , \inq_ary[7][108] , 
        \inq_ary[7][109] , \inq_ary[7][110] , \inq_ary[7][111] , 
        \inq_ary[7][112] , \inq_ary[7][113] , \inq_ary[7][114] , 
        \inq_ary[7][115] , \inq_ary[7][116] , \inq_ary[7][117] , 
        \inq_ary[7][118] , \inq_ary[7][119] , \inq_ary[7][120] , 
        \inq_ary[7][121] , \inq_ary[7][122] , \inq_ary[7][123] , 
        \inq_ary[7][124] , \inq_ary[7][125] , \inq_ary[7][126] , 
        \inq_ary[7][127] , \inq_ary[7][128] , \inq_ary[7][129] , 
        \inq_ary[7][130] , \inq_ary[7][131] , \inq_ary[7][132] , 
        \inq_ary[7][133] , \inq_ary[7][134] , \inq_ary[7][135] , 
        \inq_ary[7][136] , \inq_ary[7][137] , \inq_ary[7][138] , 
        \inq_ary[7][139] , \inq_ary[7][140] , \inq_ary[7][141] , 
        \inq_ary[7][142] , \inq_ary[7][143] , \inq_ary[7][144] , 
        \inq_ary[7][145] , \inq_ary[7][146] , \inq_ary[7][147] , 
        \inq_ary[7][148] , \inq_ary[7][149] , \inq_ary[7][150] , 
        \inq_ary[7][151] , \inq_ary[7][152] , \inq_ary[7][153] , 
        \inq_ary[7][154] , \inq_ary[7][155] , \inq_ary[7][156] , 
        \inq_ary[7][157] , \inq_ary[7][158] , \inq_ary[7][159] }), .D8({
        \inq_ary[8][0] , \inq_ary[8][1] , \inq_ary[8][2] , \inq_ary[8][3] , 
        \inq_ary[8][4] , \inq_ary[8][5] , \inq_ary[8][6] , \inq_ary[8][7] , 
        \inq_ary[8][8] , \inq_ary[8][9] , \inq_ary[8][10] , \inq_ary[8][11] , 
        \inq_ary[8][12] , \inq_ary[8][13] , \inq_ary[8][14] , \inq_ary[8][15] , 
        \inq_ary[8][16] , \inq_ary[8][17] , \inq_ary[8][18] , \inq_ary[8][19] , 
        \inq_ary[8][20] , \inq_ary[8][21] , \inq_ary[8][22] , \inq_ary[8][23] , 
        \inq_ary[8][24] , \inq_ary[8][25] , \inq_ary[8][26] , \inq_ary[8][27] , 
        \inq_ary[8][28] , \inq_ary[8][29] , \inq_ary[8][30] , \inq_ary[8][31] , 
        \inq_ary[8][32] , \inq_ary[8][33] , \inq_ary[8][34] , \inq_ary[8][35] , 
        \inq_ary[8][36] , \inq_ary[8][37] , \inq_ary[8][38] , \inq_ary[8][39] , 
        \inq_ary[8][40] , \inq_ary[8][41] , \inq_ary[8][42] , \inq_ary[8][43] , 
        \inq_ary[8][44] , \inq_ary[8][45] , \inq_ary[8][46] , \inq_ary[8][47] , 
        \inq_ary[8][48] , \inq_ary[8][49] , \inq_ary[8][50] , \inq_ary[8][51] , 
        \inq_ary[8][52] , \inq_ary[8][53] , \inq_ary[8][54] , \inq_ary[8][55] , 
        \inq_ary[8][56] , \inq_ary[8][57] , \inq_ary[8][58] , \inq_ary[8][59] , 
        \inq_ary[8][60] , \inq_ary[8][61] , \inq_ary[8][62] , \inq_ary[8][63] , 
        \inq_ary[8][64] , \inq_ary[8][65] , \inq_ary[8][66] , \inq_ary[8][67] , 
        \inq_ary[8][68] , \inq_ary[8][69] , \inq_ary[8][70] , \inq_ary[8][71] , 
        \inq_ary[8][72] , \inq_ary[8][73] , \inq_ary[8][74] , \inq_ary[8][75] , 
        \inq_ary[8][76] , \inq_ary[8][77] , \inq_ary[8][78] , \inq_ary[8][79] , 
        \inq_ary[8][80] , \inq_ary[8][81] , \inq_ary[8][82] , \inq_ary[8][83] , 
        \inq_ary[8][84] , \inq_ary[8][85] , \inq_ary[8][86] , \inq_ary[8][87] , 
        \inq_ary[8][88] , \inq_ary[8][89] , \inq_ary[8][90] , \inq_ary[8][91] , 
        \inq_ary[8][92] , \inq_ary[8][93] , \inq_ary[8][94] , \inq_ary[8][95] , 
        \inq_ary[8][96] , \inq_ary[8][97] , \inq_ary[8][98] , \inq_ary[8][99] , 
        \inq_ary[8][100] , \inq_ary[8][101] , \inq_ary[8][102] , 
        \inq_ary[8][103] , \inq_ary[8][104] , \inq_ary[8][105] , 
        \inq_ary[8][106] , \inq_ary[8][107] , \inq_ary[8][108] , 
        \inq_ary[8][109] , \inq_ary[8][110] , \inq_ary[8][111] , 
        \inq_ary[8][112] , \inq_ary[8][113] , \inq_ary[8][114] , 
        \inq_ary[8][115] , \inq_ary[8][116] , \inq_ary[8][117] , 
        \inq_ary[8][118] , \inq_ary[8][119] , \inq_ary[8][120] , 
        \inq_ary[8][121] , \inq_ary[8][122] , \inq_ary[8][123] , 
        \inq_ary[8][124] , \inq_ary[8][125] , \inq_ary[8][126] , 
        \inq_ary[8][127] , \inq_ary[8][128] , \inq_ary[8][129] , 
        \inq_ary[8][130] , \inq_ary[8][131] , \inq_ary[8][132] , 
        \inq_ary[8][133] , \inq_ary[8][134] , \inq_ary[8][135] , 
        \inq_ary[8][136] , \inq_ary[8][137] , \inq_ary[8][138] , 
        \inq_ary[8][139] , \inq_ary[8][140] , \inq_ary[8][141] , 
        \inq_ary[8][142] , \inq_ary[8][143] , \inq_ary[8][144] , 
        \inq_ary[8][145] , \inq_ary[8][146] , \inq_ary[8][147] , 
        \inq_ary[8][148] , \inq_ary[8][149] , \inq_ary[8][150] , 
        \inq_ary[8][151] , \inq_ary[8][152] , \inq_ary[8][153] , 
        \inq_ary[8][154] , \inq_ary[8][155] , \inq_ary[8][156] , 
        \inq_ary[8][157] , \inq_ary[8][158] , \inq_ary[8][159] }), .D9({
        \inq_ary[9][0] , \inq_ary[9][1] , \inq_ary[9][2] , \inq_ary[9][3] , 
        \inq_ary[9][4] , \inq_ary[9][5] , \inq_ary[9][6] , \inq_ary[9][7] , 
        \inq_ary[9][8] , \inq_ary[9][9] , \inq_ary[9][10] , \inq_ary[9][11] , 
        \inq_ary[9][12] , \inq_ary[9][13] , \inq_ary[9][14] , \inq_ary[9][15] , 
        \inq_ary[9][16] , \inq_ary[9][17] , \inq_ary[9][18] , \inq_ary[9][19] , 
        \inq_ary[9][20] , \inq_ary[9][21] , \inq_ary[9][22] , \inq_ary[9][23] , 
        \inq_ary[9][24] , \inq_ary[9][25] , \inq_ary[9][26] , \inq_ary[9][27] , 
        \inq_ary[9][28] , \inq_ary[9][29] , \inq_ary[9][30] , \inq_ary[9][31] , 
        \inq_ary[9][32] , \inq_ary[9][33] , \inq_ary[9][34] , \inq_ary[9][35] , 
        \inq_ary[9][36] , \inq_ary[9][37] , \inq_ary[9][38] , \inq_ary[9][39] , 
        \inq_ary[9][40] , \inq_ary[9][41] , \inq_ary[9][42] , \inq_ary[9][43] , 
        \inq_ary[9][44] , \inq_ary[9][45] , \inq_ary[9][46] , \inq_ary[9][47] , 
        \inq_ary[9][48] , \inq_ary[9][49] , \inq_ary[9][50] , \inq_ary[9][51] , 
        \inq_ary[9][52] , \inq_ary[9][53] , \inq_ary[9][54] , \inq_ary[9][55] , 
        \inq_ary[9][56] , \inq_ary[9][57] , \inq_ary[9][58] , \inq_ary[9][59] , 
        \inq_ary[9][60] , \inq_ary[9][61] , \inq_ary[9][62] , \inq_ary[9][63] , 
        \inq_ary[9][64] , \inq_ary[9][65] , \inq_ary[9][66] , \inq_ary[9][67] , 
        \inq_ary[9][68] , \inq_ary[9][69] , \inq_ary[9][70] , \inq_ary[9][71] , 
        \inq_ary[9][72] , \inq_ary[9][73] , \inq_ary[9][74] , \inq_ary[9][75] , 
        \inq_ary[9][76] , \inq_ary[9][77] , \inq_ary[9][78] , \inq_ary[9][79] , 
        \inq_ary[9][80] , \inq_ary[9][81] , \inq_ary[9][82] , \inq_ary[9][83] , 
        \inq_ary[9][84] , \inq_ary[9][85] , \inq_ary[9][86] , \inq_ary[9][87] , 
        \inq_ary[9][88] , \inq_ary[9][89] , \inq_ary[9][90] , \inq_ary[9][91] , 
        \inq_ary[9][92] , \inq_ary[9][93] , \inq_ary[9][94] , \inq_ary[9][95] , 
        \inq_ary[9][96] , \inq_ary[9][97] , \inq_ary[9][98] , \inq_ary[9][99] , 
        \inq_ary[9][100] , \inq_ary[9][101] , \inq_ary[9][102] , 
        \inq_ary[9][103] , \inq_ary[9][104] , \inq_ary[9][105] , 
        \inq_ary[9][106] , \inq_ary[9][107] , \inq_ary[9][108] , 
        \inq_ary[9][109] , \inq_ary[9][110] , \inq_ary[9][111] , 
        \inq_ary[9][112] , \inq_ary[9][113] , \inq_ary[9][114] , 
        \inq_ary[9][115] , \inq_ary[9][116] , \inq_ary[9][117] , 
        \inq_ary[9][118] , \inq_ary[9][119] , \inq_ary[9][120] , 
        \inq_ary[9][121] , \inq_ary[9][122] , \inq_ary[9][123] , 
        \inq_ary[9][124] , \inq_ary[9][125] , \inq_ary[9][126] , 
        \inq_ary[9][127] , \inq_ary[9][128] , \inq_ary[9][129] , 
        \inq_ary[9][130] , \inq_ary[9][131] , \inq_ary[9][132] , 
        \inq_ary[9][133] , \inq_ary[9][134] , \inq_ary[9][135] , 
        \inq_ary[9][136] , \inq_ary[9][137] , \inq_ary[9][138] , 
        \inq_ary[9][139] , \inq_ary[9][140] , \inq_ary[9][141] , 
        \inq_ary[9][142] , \inq_ary[9][143] , \inq_ary[9][144] , 
        \inq_ary[9][145] , \inq_ary[9][146] , \inq_ary[9][147] , 
        \inq_ary[9][148] , \inq_ary[9][149] , \inq_ary[9][150] , 
        \inq_ary[9][151] , \inq_ary[9][152] , \inq_ary[9][153] , 
        \inq_ary[9][154] , \inq_ary[9][155] , \inq_ary[9][156] , 
        \inq_ary[9][157] , \inq_ary[9][158] , \inq_ary[9][159] }), .D10({
        \inq_ary[10][0] , \inq_ary[10][1] , \inq_ary[10][2] , \inq_ary[10][3] , 
        \inq_ary[10][4] , \inq_ary[10][5] , \inq_ary[10][6] , \inq_ary[10][7] , 
        \inq_ary[10][8] , \inq_ary[10][9] , \inq_ary[10][10] , 
        \inq_ary[10][11] , \inq_ary[10][12] , \inq_ary[10][13] , 
        \inq_ary[10][14] , \inq_ary[10][15] , \inq_ary[10][16] , 
        \inq_ary[10][17] , \inq_ary[10][18] , \inq_ary[10][19] , 
        \inq_ary[10][20] , \inq_ary[10][21] , \inq_ary[10][22] , 
        \inq_ary[10][23] , \inq_ary[10][24] , \inq_ary[10][25] , 
        \inq_ary[10][26] , \inq_ary[10][27] , \inq_ary[10][28] , 
        \inq_ary[10][29] , \inq_ary[10][30] , \inq_ary[10][31] , 
        \inq_ary[10][32] , \inq_ary[10][33] , \inq_ary[10][34] , 
        \inq_ary[10][35] , \inq_ary[10][36] , \inq_ary[10][37] , 
        \inq_ary[10][38] , \inq_ary[10][39] , \inq_ary[10][40] , 
        \inq_ary[10][41] , \inq_ary[10][42] , \inq_ary[10][43] , 
        \inq_ary[10][44] , \inq_ary[10][45] , \inq_ary[10][46] , 
        \inq_ary[10][47] , \inq_ary[10][48] , \inq_ary[10][49] , 
        \inq_ary[10][50] , \inq_ary[10][51] , \inq_ary[10][52] , 
        \inq_ary[10][53] , \inq_ary[10][54] , \inq_ary[10][55] , 
        \inq_ary[10][56] , \inq_ary[10][57] , \inq_ary[10][58] , 
        \inq_ary[10][59] , \inq_ary[10][60] , \inq_ary[10][61] , 
        \inq_ary[10][62] , \inq_ary[10][63] , \inq_ary[10][64] , 
        \inq_ary[10][65] , \inq_ary[10][66] , \inq_ary[10][67] , 
        \inq_ary[10][68] , \inq_ary[10][69] , \inq_ary[10][70] , 
        \inq_ary[10][71] , \inq_ary[10][72] , \inq_ary[10][73] , 
        \inq_ary[10][74] , \inq_ary[10][75] , \inq_ary[10][76] , 
        \inq_ary[10][77] , \inq_ary[10][78] , \inq_ary[10][79] , 
        \inq_ary[10][80] , \inq_ary[10][81] , \inq_ary[10][82] , 
        \inq_ary[10][83] , \inq_ary[10][84] , \inq_ary[10][85] , 
        \inq_ary[10][86] , \inq_ary[10][87] , \inq_ary[10][88] , 
        \inq_ary[10][89] , \inq_ary[10][90] , \inq_ary[10][91] , 
        \inq_ary[10][92] , \inq_ary[10][93] , \inq_ary[10][94] , 
        \inq_ary[10][95] , \inq_ary[10][96] , \inq_ary[10][97] , 
        \inq_ary[10][98] , \inq_ary[10][99] , \inq_ary[10][100] , 
        \inq_ary[10][101] , \inq_ary[10][102] , \inq_ary[10][103] , 
        \inq_ary[10][104] , \inq_ary[10][105] , \inq_ary[10][106] , 
        \inq_ary[10][107] , \inq_ary[10][108] , \inq_ary[10][109] , 
        \inq_ary[10][110] , \inq_ary[10][111] , \inq_ary[10][112] , 
        \inq_ary[10][113] , \inq_ary[10][114] , \inq_ary[10][115] , 
        \inq_ary[10][116] , \inq_ary[10][117] , \inq_ary[10][118] , 
        \inq_ary[10][119] , \inq_ary[10][120] , \inq_ary[10][121] , 
        \inq_ary[10][122] , \inq_ary[10][123] , \inq_ary[10][124] , 
        \inq_ary[10][125] , \inq_ary[10][126] , \inq_ary[10][127] , 
        \inq_ary[10][128] , \inq_ary[10][129] , \inq_ary[10][130] , 
        \inq_ary[10][131] , \inq_ary[10][132] , \inq_ary[10][133] , 
        \inq_ary[10][134] , \inq_ary[10][135] , \inq_ary[10][136] , 
        \inq_ary[10][137] , \inq_ary[10][138] , \inq_ary[10][139] , 
        \inq_ary[10][140] , \inq_ary[10][141] , \inq_ary[10][142] , 
        \inq_ary[10][143] , \inq_ary[10][144] , \inq_ary[10][145] , 
        \inq_ary[10][146] , \inq_ary[10][147] , \inq_ary[10][148] , 
        \inq_ary[10][149] , \inq_ary[10][150] , \inq_ary[10][151] , 
        \inq_ary[10][152] , \inq_ary[10][153] , \inq_ary[10][154] , 
        \inq_ary[10][155] , \inq_ary[10][156] , \inq_ary[10][157] , 
        \inq_ary[10][158] , \inq_ary[10][159] }), .D11({\inq_ary[11][0] , 
        \inq_ary[11][1] , \inq_ary[11][2] , \inq_ary[11][3] , \inq_ary[11][4] , 
        \inq_ary[11][5] , \inq_ary[11][6] , \inq_ary[11][7] , \inq_ary[11][8] , 
        \inq_ary[11][9] , \inq_ary[11][10] , \inq_ary[11][11] , 
        \inq_ary[11][12] , \inq_ary[11][13] , \inq_ary[11][14] , 
        \inq_ary[11][15] , \inq_ary[11][16] , \inq_ary[11][17] , 
        \inq_ary[11][18] , \inq_ary[11][19] , \inq_ary[11][20] , 
        \inq_ary[11][21] , \inq_ary[11][22] , \inq_ary[11][23] , 
        \inq_ary[11][24] , \inq_ary[11][25] , \inq_ary[11][26] , 
        \inq_ary[11][27] , \inq_ary[11][28] , \inq_ary[11][29] , 
        \inq_ary[11][30] , \inq_ary[11][31] , \inq_ary[11][32] , 
        \inq_ary[11][33] , \inq_ary[11][34] , \inq_ary[11][35] , 
        \inq_ary[11][36] , \inq_ary[11][37] , \inq_ary[11][38] , 
        \inq_ary[11][39] , \inq_ary[11][40] , \inq_ary[11][41] , 
        \inq_ary[11][42] , \inq_ary[11][43] , \inq_ary[11][44] , 
        \inq_ary[11][45] , \inq_ary[11][46] , \inq_ary[11][47] , 
        \inq_ary[11][48] , \inq_ary[11][49] , \inq_ary[11][50] , 
        \inq_ary[11][51] , \inq_ary[11][52] , \inq_ary[11][53] , 
        \inq_ary[11][54] , \inq_ary[11][55] , \inq_ary[11][56] , 
        \inq_ary[11][57] , \inq_ary[11][58] , \inq_ary[11][59] , 
        \inq_ary[11][60] , \inq_ary[11][61] , \inq_ary[11][62] , 
        \inq_ary[11][63] , \inq_ary[11][64] , \inq_ary[11][65] , 
        \inq_ary[11][66] , \inq_ary[11][67] , \inq_ary[11][68] , 
        \inq_ary[11][69] , \inq_ary[11][70] , \inq_ary[11][71] , 
        \inq_ary[11][72] , \inq_ary[11][73] , \inq_ary[11][74] , 
        \inq_ary[11][75] , \inq_ary[11][76] , \inq_ary[11][77] , 
        \inq_ary[11][78] , \inq_ary[11][79] , \inq_ary[11][80] , 
        \inq_ary[11][81] , \inq_ary[11][82] , \inq_ary[11][83] , 
        \inq_ary[11][84] , \inq_ary[11][85] , \inq_ary[11][86] , 
        \inq_ary[11][87] , \inq_ary[11][88] , \inq_ary[11][89] , 
        \inq_ary[11][90] , \inq_ary[11][91] , \inq_ary[11][92] , 
        \inq_ary[11][93] , \inq_ary[11][94] , \inq_ary[11][95] , 
        \inq_ary[11][96] , \inq_ary[11][97] , \inq_ary[11][98] , 
        \inq_ary[11][99] , \inq_ary[11][100] , \inq_ary[11][101] , 
        \inq_ary[11][102] , \inq_ary[11][103] , \inq_ary[11][104] , 
        \inq_ary[11][105] , \inq_ary[11][106] , \inq_ary[11][107] , 
        \inq_ary[11][108] , \inq_ary[11][109] , \inq_ary[11][110] , 
        \inq_ary[11][111] , \inq_ary[11][112] , \inq_ary[11][113] , 
        \inq_ary[11][114] , \inq_ary[11][115] , \inq_ary[11][116] , 
        \inq_ary[11][117] , \inq_ary[11][118] , \inq_ary[11][119] , 
        \inq_ary[11][120] , \inq_ary[11][121] , \inq_ary[11][122] , 
        \inq_ary[11][123] , \inq_ary[11][124] , \inq_ary[11][125] , 
        \inq_ary[11][126] , \inq_ary[11][127] , \inq_ary[11][128] , 
        \inq_ary[11][129] , \inq_ary[11][130] , \inq_ary[11][131] , 
        \inq_ary[11][132] , \inq_ary[11][133] , \inq_ary[11][134] , 
        \inq_ary[11][135] , \inq_ary[11][136] , \inq_ary[11][137] , 
        \inq_ary[11][138] , \inq_ary[11][139] , \inq_ary[11][140] , 
        \inq_ary[11][141] , \inq_ary[11][142] , \inq_ary[11][143] , 
        \inq_ary[11][144] , \inq_ary[11][145] , \inq_ary[11][146] , 
        \inq_ary[11][147] , \inq_ary[11][148] , \inq_ary[11][149] , 
        \inq_ary[11][150] , \inq_ary[11][151] , \inq_ary[11][152] , 
        \inq_ary[11][153] , \inq_ary[11][154] , \inq_ary[11][155] , 
        \inq_ary[11][156] , \inq_ary[11][157] , \inq_ary[11][158] , 
        \inq_ary[11][159] }), .D12({\inq_ary[12][0] , \inq_ary[12][1] , 
        \inq_ary[12][2] , \inq_ary[12][3] , \inq_ary[12][4] , \inq_ary[12][5] , 
        \inq_ary[12][6] , \inq_ary[12][7] , \inq_ary[12][8] , \inq_ary[12][9] , 
        \inq_ary[12][10] , \inq_ary[12][11] , \inq_ary[12][12] , 
        \inq_ary[12][13] , \inq_ary[12][14] , \inq_ary[12][15] , 
        \inq_ary[12][16] , \inq_ary[12][17] , \inq_ary[12][18] , 
        \inq_ary[12][19] , \inq_ary[12][20] , \inq_ary[12][21] , 
        \inq_ary[12][22] , \inq_ary[12][23] , \inq_ary[12][24] , 
        \inq_ary[12][25] , \inq_ary[12][26] , \inq_ary[12][27] , 
        \inq_ary[12][28] , \inq_ary[12][29] , \inq_ary[12][30] , 
        \inq_ary[12][31] , \inq_ary[12][32] , \inq_ary[12][33] , 
        \inq_ary[12][34] , \inq_ary[12][35] , \inq_ary[12][36] , 
        \inq_ary[12][37] , \inq_ary[12][38] , \inq_ary[12][39] , 
        \inq_ary[12][40] , \inq_ary[12][41] , \inq_ary[12][42] , 
        \inq_ary[12][43] , \inq_ary[12][44] , \inq_ary[12][45] , 
        \inq_ary[12][46] , \inq_ary[12][47] , \inq_ary[12][48] , 
        \inq_ary[12][49] , \inq_ary[12][50] , \inq_ary[12][51] , 
        \inq_ary[12][52] , \inq_ary[12][53] , \inq_ary[12][54] , 
        \inq_ary[12][55] , \inq_ary[12][56] , \inq_ary[12][57] , 
        \inq_ary[12][58] , \inq_ary[12][59] , \inq_ary[12][60] , 
        \inq_ary[12][61] , \inq_ary[12][62] , \inq_ary[12][63] , 
        \inq_ary[12][64] , \inq_ary[12][65] , \inq_ary[12][66] , 
        \inq_ary[12][67] , \inq_ary[12][68] , \inq_ary[12][69] , 
        \inq_ary[12][70] , \inq_ary[12][71] , \inq_ary[12][72] , 
        \inq_ary[12][73] , \inq_ary[12][74] , \inq_ary[12][75] , 
        \inq_ary[12][76] , \inq_ary[12][77] , \inq_ary[12][78] , 
        \inq_ary[12][79] , \inq_ary[12][80] , \inq_ary[12][81] , 
        \inq_ary[12][82] , \inq_ary[12][83] , \inq_ary[12][84] , 
        \inq_ary[12][85] , \inq_ary[12][86] , \inq_ary[12][87] , 
        \inq_ary[12][88] , \inq_ary[12][89] , \inq_ary[12][90] , 
        \inq_ary[12][91] , \inq_ary[12][92] , \inq_ary[12][93] , 
        \inq_ary[12][94] , \inq_ary[12][95] , \inq_ary[12][96] , 
        \inq_ary[12][97] , \inq_ary[12][98] , \inq_ary[12][99] , 
        \inq_ary[12][100] , \inq_ary[12][101] , \inq_ary[12][102] , 
        \inq_ary[12][103] , \inq_ary[12][104] , \inq_ary[12][105] , 
        \inq_ary[12][106] , \inq_ary[12][107] , \inq_ary[12][108] , 
        \inq_ary[12][109] , \inq_ary[12][110] , \inq_ary[12][111] , 
        \inq_ary[12][112] , \inq_ary[12][113] , \inq_ary[12][114] , 
        \inq_ary[12][115] , \inq_ary[12][116] , \inq_ary[12][117] , 
        \inq_ary[12][118] , \inq_ary[12][119] , \inq_ary[12][120] , 
        \inq_ary[12][121] , \inq_ary[12][122] , \inq_ary[12][123] , 
        \inq_ary[12][124] , \inq_ary[12][125] , \inq_ary[12][126] , 
        \inq_ary[12][127] , \inq_ary[12][128] , \inq_ary[12][129] , 
        \inq_ary[12][130] , \inq_ary[12][131] , \inq_ary[12][132] , 
        \inq_ary[12][133] , \inq_ary[12][134] , \inq_ary[12][135] , 
        \inq_ary[12][136] , \inq_ary[12][137] , \inq_ary[12][138] , 
        \inq_ary[12][139] , \inq_ary[12][140] , \inq_ary[12][141] , 
        \inq_ary[12][142] , \inq_ary[12][143] , \inq_ary[12][144] , 
        \inq_ary[12][145] , \inq_ary[12][146] , \inq_ary[12][147] , 
        \inq_ary[12][148] , \inq_ary[12][149] , \inq_ary[12][150] , 
        \inq_ary[12][151] , \inq_ary[12][152] , \inq_ary[12][153] , 
        \inq_ary[12][154] , \inq_ary[12][155] , \inq_ary[12][156] , 
        \inq_ary[12][157] , \inq_ary[12][158] , \inq_ary[12][159] }), .D13({
        \inq_ary[13][0] , \inq_ary[13][1] , \inq_ary[13][2] , \inq_ary[13][3] , 
        \inq_ary[13][4] , \inq_ary[13][5] , \inq_ary[13][6] , \inq_ary[13][7] , 
        \inq_ary[13][8] , \inq_ary[13][9] , \inq_ary[13][10] , 
        \inq_ary[13][11] , \inq_ary[13][12] , \inq_ary[13][13] , 
        \inq_ary[13][14] , \inq_ary[13][15] , \inq_ary[13][16] , 
        \inq_ary[13][17] , \inq_ary[13][18] , \inq_ary[13][19] , 
        \inq_ary[13][20] , \inq_ary[13][21] , \inq_ary[13][22] , 
        \inq_ary[13][23] , \inq_ary[13][24] , \inq_ary[13][25] , 
        \inq_ary[13][26] , \inq_ary[13][27] , \inq_ary[13][28] , 
        \inq_ary[13][29] , \inq_ary[13][30] , \inq_ary[13][31] , 
        \inq_ary[13][32] , \inq_ary[13][33] , \inq_ary[13][34] , 
        \inq_ary[13][35] , \inq_ary[13][36] , \inq_ary[13][37] , 
        \inq_ary[13][38] , \inq_ary[13][39] , \inq_ary[13][40] , 
        \inq_ary[13][41] , \inq_ary[13][42] , \inq_ary[13][43] , 
        \inq_ary[13][44] , \inq_ary[13][45] , \inq_ary[13][46] , 
        \inq_ary[13][47] , \inq_ary[13][48] , \inq_ary[13][49] , 
        \inq_ary[13][50] , \inq_ary[13][51] , \inq_ary[13][52] , 
        \inq_ary[13][53] , \inq_ary[13][54] , \inq_ary[13][55] , 
        \inq_ary[13][56] , \inq_ary[13][57] , \inq_ary[13][58] , 
        \inq_ary[13][59] , \inq_ary[13][60] , \inq_ary[13][61] , 
        \inq_ary[13][62] , \inq_ary[13][63] , \inq_ary[13][64] , 
        \inq_ary[13][65] , \inq_ary[13][66] , \inq_ary[13][67] , 
        \inq_ary[13][68] , \inq_ary[13][69] , \inq_ary[13][70] , 
        \inq_ary[13][71] , \inq_ary[13][72] , \inq_ary[13][73] , 
        \inq_ary[13][74] , \inq_ary[13][75] , \inq_ary[13][76] , 
        \inq_ary[13][77] , \inq_ary[13][78] , \inq_ary[13][79] , 
        \inq_ary[13][80] , \inq_ary[13][81] , \inq_ary[13][82] , 
        \inq_ary[13][83] , \inq_ary[13][84] , \inq_ary[13][85] , 
        \inq_ary[13][86] , \inq_ary[13][87] , \inq_ary[13][88] , 
        \inq_ary[13][89] , \inq_ary[13][90] , \inq_ary[13][91] , 
        \inq_ary[13][92] , \inq_ary[13][93] , \inq_ary[13][94] , 
        \inq_ary[13][95] , \inq_ary[13][96] , \inq_ary[13][97] , 
        \inq_ary[13][98] , \inq_ary[13][99] , \inq_ary[13][100] , 
        \inq_ary[13][101] , \inq_ary[13][102] , \inq_ary[13][103] , 
        \inq_ary[13][104] , \inq_ary[13][105] , \inq_ary[13][106] , 
        \inq_ary[13][107] , \inq_ary[13][108] , \inq_ary[13][109] , 
        \inq_ary[13][110] , \inq_ary[13][111] , \inq_ary[13][112] , 
        \inq_ary[13][113] , \inq_ary[13][114] , \inq_ary[13][115] , 
        \inq_ary[13][116] , \inq_ary[13][117] , \inq_ary[13][118] , 
        \inq_ary[13][119] , \inq_ary[13][120] , \inq_ary[13][121] , 
        \inq_ary[13][122] , \inq_ary[13][123] , \inq_ary[13][124] , 
        \inq_ary[13][125] , \inq_ary[13][126] , \inq_ary[13][127] , 
        \inq_ary[13][128] , \inq_ary[13][129] , \inq_ary[13][130] , 
        \inq_ary[13][131] , \inq_ary[13][132] , \inq_ary[13][133] , 
        \inq_ary[13][134] , \inq_ary[13][135] , \inq_ary[13][136] , 
        \inq_ary[13][137] , \inq_ary[13][138] , \inq_ary[13][139] , 
        \inq_ary[13][140] , \inq_ary[13][141] , \inq_ary[13][142] , 
        \inq_ary[13][143] , \inq_ary[13][144] , \inq_ary[13][145] , 
        \inq_ary[13][146] , \inq_ary[13][147] , \inq_ary[13][148] , 
        \inq_ary[13][149] , \inq_ary[13][150] , \inq_ary[13][151] , 
        \inq_ary[13][152] , \inq_ary[13][153] , \inq_ary[13][154] , 
        \inq_ary[13][155] , \inq_ary[13][156] , \inq_ary[13][157] , 
        \inq_ary[13][158] , \inq_ary[13][159] }), .D14({\inq_ary[14][0] , 
        \inq_ary[14][1] , \inq_ary[14][2] , \inq_ary[14][3] , \inq_ary[14][4] , 
        \inq_ary[14][5] , \inq_ary[14][6] , \inq_ary[14][7] , \inq_ary[14][8] , 
        \inq_ary[14][9] , \inq_ary[14][10] , \inq_ary[14][11] , 
        \inq_ary[14][12] , \inq_ary[14][13] , \inq_ary[14][14] , 
        \inq_ary[14][15] , \inq_ary[14][16] , \inq_ary[14][17] , 
        \inq_ary[14][18] , \inq_ary[14][19] , \inq_ary[14][20] , 
        \inq_ary[14][21] , \inq_ary[14][22] , \inq_ary[14][23] , 
        \inq_ary[14][24] , \inq_ary[14][25] , \inq_ary[14][26] , 
        \inq_ary[14][27] , \inq_ary[14][28] , \inq_ary[14][29] , 
        \inq_ary[14][30] , \inq_ary[14][31] , \inq_ary[14][32] , 
        \inq_ary[14][33] , \inq_ary[14][34] , \inq_ary[14][35] , 
        \inq_ary[14][36] , \inq_ary[14][37] , \inq_ary[14][38] , 
        \inq_ary[14][39] , \inq_ary[14][40] , \inq_ary[14][41] , 
        \inq_ary[14][42] , \inq_ary[14][43] , \inq_ary[14][44] , 
        \inq_ary[14][45] , \inq_ary[14][46] , \inq_ary[14][47] , 
        \inq_ary[14][48] , \inq_ary[14][49] , \inq_ary[14][50] , 
        \inq_ary[14][51] , \inq_ary[14][52] , \inq_ary[14][53] , 
        \inq_ary[14][54] , \inq_ary[14][55] , \inq_ary[14][56] , 
        \inq_ary[14][57] , \inq_ary[14][58] , \inq_ary[14][59] , 
        \inq_ary[14][60] , \inq_ary[14][61] , \inq_ary[14][62] , 
        \inq_ary[14][63] , \inq_ary[14][64] , \inq_ary[14][65] , 
        \inq_ary[14][66] , \inq_ary[14][67] , \inq_ary[14][68] , 
        \inq_ary[14][69] , \inq_ary[14][70] , \inq_ary[14][71] , 
        \inq_ary[14][72] , \inq_ary[14][73] , \inq_ary[14][74] , 
        \inq_ary[14][75] , \inq_ary[14][76] , \inq_ary[14][77] , 
        \inq_ary[14][78] , \inq_ary[14][79] , \inq_ary[14][80] , 
        \inq_ary[14][81] , \inq_ary[14][82] , \inq_ary[14][83] , 
        \inq_ary[14][84] , \inq_ary[14][85] , \inq_ary[14][86] , 
        \inq_ary[14][87] , \inq_ary[14][88] , \inq_ary[14][89] , 
        \inq_ary[14][90] , \inq_ary[14][91] , \inq_ary[14][92] , 
        \inq_ary[14][93] , \inq_ary[14][94] , \inq_ary[14][95] , 
        \inq_ary[14][96] , \inq_ary[14][97] , \inq_ary[14][98] , 
        \inq_ary[14][99] , \inq_ary[14][100] , \inq_ary[14][101] , 
        \inq_ary[14][102] , \inq_ary[14][103] , \inq_ary[14][104] , 
        \inq_ary[14][105] , \inq_ary[14][106] , \inq_ary[14][107] , 
        \inq_ary[14][108] , \inq_ary[14][109] , \inq_ary[14][110] , 
        \inq_ary[14][111] , \inq_ary[14][112] , \inq_ary[14][113] , 
        \inq_ary[14][114] , \inq_ary[14][115] , \inq_ary[14][116] , 
        \inq_ary[14][117] , \inq_ary[14][118] , \inq_ary[14][119] , 
        \inq_ary[14][120] , \inq_ary[14][121] , \inq_ary[14][122] , 
        \inq_ary[14][123] , \inq_ary[14][124] , \inq_ary[14][125] , 
        \inq_ary[14][126] , \inq_ary[14][127] , \inq_ary[14][128] , 
        \inq_ary[14][129] , \inq_ary[14][130] , \inq_ary[14][131] , 
        \inq_ary[14][132] , \inq_ary[14][133] , \inq_ary[14][134] , 
        \inq_ary[14][135] , \inq_ary[14][136] , \inq_ary[14][137] , 
        \inq_ary[14][138] , \inq_ary[14][139] , \inq_ary[14][140] , 
        \inq_ary[14][141] , \inq_ary[14][142] , \inq_ary[14][143] , 
        \inq_ary[14][144] , \inq_ary[14][145] , \inq_ary[14][146] , 
        \inq_ary[14][147] , \inq_ary[14][148] , \inq_ary[14][149] , 
        \inq_ary[14][150] , \inq_ary[14][151] , \inq_ary[14][152] , 
        \inq_ary[14][153] , \inq_ary[14][154] , \inq_ary[14][155] , 
        \inq_ary[14][156] , \inq_ary[14][157] , \inq_ary[14][158] , 
        \inq_ary[14][159] }), .D15({\inq_ary[15][0] , \inq_ary[15][1] , 
        \inq_ary[15][2] , \inq_ary[15][3] , \inq_ary[15][4] , \inq_ary[15][5] , 
        \inq_ary[15][6] , \inq_ary[15][7] , \inq_ary[15][8] , \inq_ary[15][9] , 
        \inq_ary[15][10] , \inq_ary[15][11] , \inq_ary[15][12] , 
        \inq_ary[15][13] , \inq_ary[15][14] , \inq_ary[15][15] , 
        \inq_ary[15][16] , \inq_ary[15][17] , \inq_ary[15][18] , 
        \inq_ary[15][19] , \inq_ary[15][20] , \inq_ary[15][21] , 
        \inq_ary[15][22] , \inq_ary[15][23] , \inq_ary[15][24] , 
        \inq_ary[15][25] , \inq_ary[15][26] , \inq_ary[15][27] , 
        \inq_ary[15][28] , \inq_ary[15][29] , \inq_ary[15][30] , 
        \inq_ary[15][31] , \inq_ary[15][32] , \inq_ary[15][33] , 
        \inq_ary[15][34] , \inq_ary[15][35] , \inq_ary[15][36] , 
        \inq_ary[15][37] , \inq_ary[15][38] , \inq_ary[15][39] , 
        \inq_ary[15][40] , \inq_ary[15][41] , \inq_ary[15][42] , 
        \inq_ary[15][43] , \inq_ary[15][44] , \inq_ary[15][45] , 
        \inq_ary[15][46] , \inq_ary[15][47] , \inq_ary[15][48] , 
        \inq_ary[15][49] , \inq_ary[15][50] , \inq_ary[15][51] , 
        \inq_ary[15][52] , \inq_ary[15][53] , \inq_ary[15][54] , 
        \inq_ary[15][55] , \inq_ary[15][56] , \inq_ary[15][57] , 
        \inq_ary[15][58] , \inq_ary[15][59] , \inq_ary[15][60] , 
        \inq_ary[15][61] , \inq_ary[15][62] , \inq_ary[15][63] , 
        \inq_ary[15][64] , \inq_ary[15][65] , \inq_ary[15][66] , 
        \inq_ary[15][67] , \inq_ary[15][68] , \inq_ary[15][69] , 
        \inq_ary[15][70] , \inq_ary[15][71] , \inq_ary[15][72] , 
        \inq_ary[15][73] , \inq_ary[15][74] , \inq_ary[15][75] , 
        \inq_ary[15][76] , \inq_ary[15][77] , \inq_ary[15][78] , 
        \inq_ary[15][79] , \inq_ary[15][80] , \inq_ary[15][81] , 
        \inq_ary[15][82] , \inq_ary[15][83] , \inq_ary[15][84] , 
        \inq_ary[15][85] , \inq_ary[15][86] , \inq_ary[15][87] , 
        \inq_ary[15][88] , \inq_ary[15][89] , \inq_ary[15][90] , 
        \inq_ary[15][91] , \inq_ary[15][92] , \inq_ary[15][93] , 
        \inq_ary[15][94] , \inq_ary[15][95] , \inq_ary[15][96] , 
        \inq_ary[15][97] , \inq_ary[15][98] , \inq_ary[15][99] , 
        \inq_ary[15][100] , \inq_ary[15][101] , \inq_ary[15][102] , 
        \inq_ary[15][103] , \inq_ary[15][104] , \inq_ary[15][105] , 
        \inq_ary[15][106] , \inq_ary[15][107] , \inq_ary[15][108] , 
        \inq_ary[15][109] , \inq_ary[15][110] , \inq_ary[15][111] , 
        \inq_ary[15][112] , \inq_ary[15][113] , \inq_ary[15][114] , 
        \inq_ary[15][115] , \inq_ary[15][116] , \inq_ary[15][117] , 
        \inq_ary[15][118] , \inq_ary[15][119] , \inq_ary[15][120] , 
        \inq_ary[15][121] , \inq_ary[15][122] , \inq_ary[15][123] , 
        \inq_ary[15][124] , \inq_ary[15][125] , \inq_ary[15][126] , 
        \inq_ary[15][127] , \inq_ary[15][128] , \inq_ary[15][129] , 
        \inq_ary[15][130] , \inq_ary[15][131] , \inq_ary[15][132] , 
        \inq_ary[15][133] , \inq_ary[15][134] , \inq_ary[15][135] , 
        \inq_ary[15][136] , \inq_ary[15][137] , \inq_ary[15][138] , 
        \inq_ary[15][139] , \inq_ary[15][140] , \inq_ary[15][141] , 
        \inq_ary[15][142] , \inq_ary[15][143] , \inq_ary[15][144] , 
        \inq_ary[15][145] , \inq_ary[15][146] , \inq_ary[15][147] , 
        \inq_ary[15][148] , \inq_ary[15][149] , \inq_ary[15][150] , 
        \inq_ary[15][151] , \inq_ary[15][152] , \inq_ary[15][153] , 
        \inq_ary[15][154] , \inq_ary[15][155] , \inq_ary[15][156] , 
        \inq_ary[15][157] , \inq_ary[15][158] , \inq_ary[15][159] }), .S0(N95), 
        .S1(N96), .S2(N97), .S3(N98), .Z({N581, N580, N579, N578, N577, N576, 
        N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, 
        N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, 
        N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, 
        N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, 
        N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, 
        N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, 
        N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, 
        N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, 
        N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, 
        N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, 
        N431, N430, N429, N428, N427, N426, N425, N424, N423, N422}) );
  GTECH_BUF B_87 ( .A(wrptr_d1[0]), .Z(N95) );
  GTECH_BUF B_88 ( .A(wrptr_d1[1]), .Z(N96) );
  GTECH_BUF B_89 ( .A(wrptr_d1[2]), .Z(N97) );
  GTECH_BUF B_90 ( .A(wrptr_d1[3]), .Z(N98) );
  GTECH_NOT I_8 ( .A(reset_l), .Z(N259) );
  GTECH_AND2 C25083 ( .A(wr_en_d1), .B(word_wen_d1[0]), .Z(N582) );
  GTECH_NOT I_9 ( .A(rst_tri_en), .Z(N583) );
  GTECH_AND2 C25085 ( .A(wr_en_d1), .B(word_wen_d1[1]), .Z(N584) );
  GTECH_AND2 C25086 ( .A(wr_en_d1), .B(word_wen_d1[2]), .Z(N585) );
  GTECH_AND2 C25087 ( .A(wr_en_d1), .B(word_wen_d1[3]), .Z(N586) );
  GTECH_AND2 C25090 ( .A(wr_en_d1), .B(N583), .Z(N587) );
  GTECH_NOT I_10 ( .A(N587), .Z(N588) );
  GTECH_AND2 C25093 ( .A(N998), .B(N583), .Z(N589) );
  GTECH_AND2 C25094 ( .A(N582), .B(byte_wen_d1[0]), .Z(N998) );
  GTECH_NOT I_11 ( .A(N589), .Z(N590) );
  GTECH_AND2 C25097 ( .A(N999), .B(N583), .Z(N592) );
  GTECH_AND2 C25098 ( .A(N584), .B(byte_wen_d1[0]), .Z(N999) );
  GTECH_NOT I_12 ( .A(N592), .Z(N593) );
  GTECH_AND2 C25101 ( .A(N1000), .B(N583), .Z(N595) );
  GTECH_AND2 C25102 ( .A(N585), .B(byte_wen_d1[0]), .Z(N1000) );
  GTECH_NOT I_13 ( .A(N595), .Z(N596) );
  GTECH_AND2 C25105 ( .A(N1001), .B(N583), .Z(N598) );
  GTECH_AND2 C25106 ( .A(N586), .B(byte_wen_d1[0]), .Z(N1001) );
  GTECH_NOT I_14 ( .A(N598), .Z(N599) );
  GTECH_AND2 C25109 ( .A(N1002), .B(N583), .Z(N605) );
  GTECH_AND2 C25110 ( .A(N582), .B(byte_wen_d1[1]), .Z(N1002) );
  GTECH_NOT I_15 ( .A(N605), .Z(N606) );
  GTECH_AND2 C25113 ( .A(N1003), .B(N583), .Z(N608) );
  GTECH_AND2 C25114 ( .A(N584), .B(byte_wen_d1[1]), .Z(N1003) );
  GTECH_NOT I_16 ( .A(N608), .Z(N609) );
  GTECH_AND2 C25117 ( .A(N1004), .B(N583), .Z(N611) );
  GTECH_AND2 C25118 ( .A(N585), .B(byte_wen_d1[1]), .Z(N1004) );
  GTECH_NOT I_17 ( .A(N611), .Z(N612) );
  GTECH_AND2 C25121 ( .A(N1005), .B(N583), .Z(N614) );
  GTECH_AND2 C25122 ( .A(N586), .B(byte_wen_d1[1]), .Z(N1005) );
  GTECH_NOT I_18 ( .A(N614), .Z(N615) );
  GTECH_AND2 C25125 ( .A(N1006), .B(N583), .Z(N621) );
  GTECH_AND2 C25126 ( .A(N582), .B(byte_wen_d1[2]), .Z(N1006) );
  GTECH_NOT I_19 ( .A(N621), .Z(N622) );
  GTECH_AND2 C25129 ( .A(N1007), .B(N583), .Z(N624) );
  GTECH_AND2 C25130 ( .A(N584), .B(byte_wen_d1[2]), .Z(N1007) );
  GTECH_NOT I_20 ( .A(N624), .Z(N625) );
  GTECH_AND2 C25133 ( .A(N1008), .B(N583), .Z(N627) );
  GTECH_AND2 C25134 ( .A(N585), .B(byte_wen_d1[2]), .Z(N1008) );
  GTECH_NOT I_21 ( .A(N627), .Z(N628) );
  GTECH_AND2 C25137 ( .A(N1009), .B(N583), .Z(N630) );
  GTECH_AND2 C25138 ( .A(N586), .B(byte_wen_d1[2]), .Z(N1009) );
  GTECH_NOT I_22 ( .A(N630), .Z(N631) );
  GTECH_AND2 C25141 ( .A(N1010), .B(N583), .Z(N637) );
  GTECH_AND2 C25142 ( .A(N582), .B(byte_wen_d1[3]), .Z(N1010) );
  GTECH_NOT I_23 ( .A(N637), .Z(N638) );
  GTECH_AND2 C25145 ( .A(N1011), .B(N583), .Z(N640) );
  GTECH_AND2 C25146 ( .A(N584), .B(byte_wen_d1[3]), .Z(N1011) );
  GTECH_NOT I_24 ( .A(N640), .Z(N641) );
  GTECH_AND2 C25149 ( .A(N1012), .B(N583), .Z(N643) );
  GTECH_AND2 C25150 ( .A(N585), .B(byte_wen_d1[3]), .Z(N1012) );
  GTECH_NOT I_25 ( .A(N643), .Z(N644) );
  GTECH_AND2 C25153 ( .A(N1013), .B(N583), .Z(N646) );
  GTECH_AND2 C25154 ( .A(N586), .B(byte_wen_d1[3]), .Z(N1013) );
  GTECH_NOT I_26 ( .A(N646), .Z(N647) );
  GTECH_AND2 C25157 ( .A(N1014), .B(N583), .Z(N653) );
  GTECH_AND2 C25158 ( .A(N582), .B(byte_wen_d1[4]), .Z(N1014) );
  GTECH_NOT I_27 ( .A(N653), .Z(N654) );
  GTECH_AND2 C25161 ( .A(N1015), .B(N583), .Z(N656) );
  GTECH_AND2 C25162 ( .A(N584), .B(byte_wen_d1[4]), .Z(N1015) );
  GTECH_NOT I_28 ( .A(N656), .Z(N657) );
  GTECH_AND2 C25165 ( .A(N1016), .B(N583), .Z(N659) );
  GTECH_AND2 C25166 ( .A(N585), .B(byte_wen_d1[4]), .Z(N1016) );
  GTECH_NOT I_29 ( .A(N659), .Z(N660) );
  GTECH_AND2 C25169 ( .A(N1017), .B(N583), .Z(N662) );
  GTECH_AND2 C25170 ( .A(N586), .B(byte_wen_d1[4]), .Z(N1017) );
  GTECH_NOT I_30 ( .A(N662), .Z(N663) );
  GTECH_AND2 C25173 ( .A(N1018), .B(N583), .Z(N669) );
  GTECH_AND2 C25174 ( .A(N582), .B(byte_wen_d1[5]), .Z(N1018) );
  GTECH_NOT I_31 ( .A(N669), .Z(N670) );
  GTECH_AND2 C25177 ( .A(N1019), .B(N583), .Z(N672) );
  GTECH_AND2 C25178 ( .A(N584), .B(byte_wen_d1[5]), .Z(N1019) );
  GTECH_NOT I_32 ( .A(N672), .Z(N673) );
  GTECH_AND2 C25181 ( .A(N1020), .B(N583), .Z(N675) );
  GTECH_AND2 C25182 ( .A(N585), .B(byte_wen_d1[5]), .Z(N1020) );
  GTECH_NOT I_33 ( .A(N675), .Z(N676) );
  GTECH_AND2 C25185 ( .A(N1021), .B(N583), .Z(N678) );
  GTECH_AND2 C25186 ( .A(N586), .B(byte_wen_d1[5]), .Z(N1021) );
  GTECH_NOT I_34 ( .A(N678), .Z(N679) );
  GTECH_AND2 C25189 ( .A(N1022), .B(N583), .Z(N685) );
  GTECH_AND2 C25190 ( .A(N582), .B(byte_wen_d1[6]), .Z(N1022) );
  GTECH_NOT I_35 ( .A(N685), .Z(N686) );
  GTECH_AND2 C25193 ( .A(N1023), .B(N583), .Z(N688) );
  GTECH_AND2 C25194 ( .A(N584), .B(byte_wen_d1[6]), .Z(N1023) );
  GTECH_NOT I_36 ( .A(N688), .Z(N689) );
  GTECH_AND2 C25197 ( .A(N1024), .B(N583), .Z(N691) );
  GTECH_AND2 C25198 ( .A(N585), .B(byte_wen_d1[6]), .Z(N1024) );
  GTECH_NOT I_37 ( .A(N691), .Z(N692) );
  GTECH_AND2 C25201 ( .A(N1025), .B(N583), .Z(N694) );
  GTECH_AND2 C25202 ( .A(N586), .B(byte_wen_d1[6]), .Z(N1025) );
  GTECH_NOT I_38 ( .A(N694), .Z(N695) );
  GTECH_AND2 C25205 ( .A(N1026), .B(N583), .Z(N701) );
  GTECH_AND2 C25206 ( .A(N582), .B(byte_wen_d1[7]), .Z(N1026) );
  GTECH_NOT I_39 ( .A(N701), .Z(N702) );
  GTECH_AND2 C25209 ( .A(N1027), .B(N583), .Z(N704) );
  GTECH_AND2 C25210 ( .A(N584), .B(byte_wen_d1[7]), .Z(N1027) );
  GTECH_NOT I_40 ( .A(N704), .Z(N705) );
  GTECH_AND2 C25213 ( .A(N1028), .B(N583), .Z(N707) );
  GTECH_AND2 C25214 ( .A(N585), .B(byte_wen_d1[7]), .Z(N1028) );
  GTECH_NOT I_41 ( .A(N707), .Z(N708) );
  GTECH_AND2 C25217 ( .A(N1029), .B(N583), .Z(N710) );
  GTECH_AND2 C25218 ( .A(N586), .B(byte_wen_d1[7]), .Z(N1029) );
  GTECH_NOT I_42 ( .A(N710), .Z(N711) );
  GTECH_AND2 C25221 ( .A(N1030), .B(N583), .Z(N717) );
  GTECH_AND2 C25222 ( .A(N582), .B(byte_wen_d1[8]), .Z(N1030) );
  GTECH_NOT I_43 ( .A(N717), .Z(N718) );
  GTECH_AND2 C25225 ( .A(N1031), .B(N583), .Z(N720) );
  GTECH_AND2 C25226 ( .A(N584), .B(byte_wen_d1[8]), .Z(N1031) );
  GTECH_NOT I_44 ( .A(N720), .Z(N721) );
  GTECH_AND2 C25229 ( .A(N1032), .B(N583), .Z(N723) );
  GTECH_AND2 C25230 ( .A(N585), .B(byte_wen_d1[8]), .Z(N1032) );
  GTECH_NOT I_45 ( .A(N723), .Z(N724) );
  GTECH_AND2 C25233 ( .A(N1033), .B(N583), .Z(N726) );
  GTECH_AND2 C25234 ( .A(N586), .B(byte_wen_d1[8]), .Z(N1033) );
  GTECH_NOT I_46 ( .A(N726), .Z(N727) );
  GTECH_AND2 C25237 ( .A(N1034), .B(N583), .Z(N733) );
  GTECH_AND2 C25238 ( .A(N582), .B(byte_wen_d1[9]), .Z(N1034) );
  GTECH_NOT I_47 ( .A(N733), .Z(N734) );
  GTECH_AND2 C25241 ( .A(N1035), .B(N583), .Z(N736) );
  GTECH_AND2 C25242 ( .A(N584), .B(byte_wen_d1[9]), .Z(N1035) );
  GTECH_NOT I_48 ( .A(N736), .Z(N737) );
  GTECH_AND2 C25245 ( .A(N1036), .B(N583), .Z(N739) );
  GTECH_AND2 C25246 ( .A(N585), .B(byte_wen_d1[9]), .Z(N1036) );
  GTECH_NOT I_49 ( .A(N739), .Z(N740) );
  GTECH_AND2 C25249 ( .A(N1037), .B(N583), .Z(N742) );
  GTECH_AND2 C25250 ( .A(N586), .B(byte_wen_d1[9]), .Z(N1037) );
  GTECH_NOT I_50 ( .A(N742), .Z(N743) );
  GTECH_AND2 C25253 ( .A(N1038), .B(N583), .Z(N749) );
  GTECH_AND2 C25254 ( .A(N582), .B(byte_wen_d1[10]), .Z(N1038) );
  GTECH_NOT I_51 ( .A(N749), .Z(N750) );
  GTECH_AND2 C25257 ( .A(N1039), .B(N583), .Z(N752) );
  GTECH_AND2 C25258 ( .A(N584), .B(byte_wen_d1[10]), .Z(N1039) );
  GTECH_NOT I_52 ( .A(N752), .Z(N753) );
  GTECH_AND2 C25261 ( .A(N1040), .B(N583), .Z(N755) );
  GTECH_AND2 C25262 ( .A(N585), .B(byte_wen_d1[10]), .Z(N1040) );
  GTECH_NOT I_53 ( .A(N755), .Z(N756) );
  GTECH_AND2 C25265 ( .A(N1041), .B(N583), .Z(N758) );
  GTECH_AND2 C25266 ( .A(N586), .B(byte_wen_d1[10]), .Z(N1041) );
  GTECH_NOT I_54 ( .A(N758), .Z(N759) );
  GTECH_AND2 C25269 ( .A(N1042), .B(N583), .Z(N765) );
  GTECH_AND2 C25270 ( .A(N582), .B(byte_wen_d1[11]), .Z(N1042) );
  GTECH_NOT I_55 ( .A(N765), .Z(N766) );
  GTECH_AND2 C25273 ( .A(N1043), .B(N583), .Z(N768) );
  GTECH_AND2 C25274 ( .A(N584), .B(byte_wen_d1[11]), .Z(N1043) );
  GTECH_NOT I_56 ( .A(N768), .Z(N769) );
  GTECH_AND2 C25277 ( .A(N1044), .B(N583), .Z(N771) );
  GTECH_AND2 C25278 ( .A(N585), .B(byte_wen_d1[11]), .Z(N1044) );
  GTECH_NOT I_57 ( .A(N771), .Z(N772) );
  GTECH_AND2 C25281 ( .A(N1045), .B(N583), .Z(N774) );
  GTECH_AND2 C25282 ( .A(N586), .B(byte_wen_d1[11]), .Z(N1045) );
  GTECH_NOT I_58 ( .A(N774), .Z(N775) );
  GTECH_AND2 C25285 ( .A(N1046), .B(N583), .Z(N781) );
  GTECH_AND2 C25286 ( .A(N582), .B(byte_wen_d1[12]), .Z(N1046) );
  GTECH_NOT I_59 ( .A(N781), .Z(N782) );
  GTECH_AND2 C25289 ( .A(N1047), .B(N583), .Z(N784) );
  GTECH_AND2 C25290 ( .A(N584), .B(byte_wen_d1[12]), .Z(N1047) );
  GTECH_NOT I_60 ( .A(N784), .Z(N785) );
  GTECH_AND2 C25293 ( .A(N1048), .B(N583), .Z(N787) );
  GTECH_AND2 C25294 ( .A(N585), .B(byte_wen_d1[12]), .Z(N1048) );
  GTECH_NOT I_61 ( .A(N787), .Z(N788) );
  GTECH_AND2 C25297 ( .A(N1049), .B(N583), .Z(N790) );
  GTECH_AND2 C25298 ( .A(N586), .B(byte_wen_d1[12]), .Z(N1049) );
  GTECH_NOT I_62 ( .A(N790), .Z(N791) );
  GTECH_AND2 C25301 ( .A(N1050), .B(N583), .Z(N797) );
  GTECH_AND2 C25302 ( .A(N582), .B(byte_wen_d1[13]), .Z(N1050) );
  GTECH_NOT I_63 ( .A(N797), .Z(N798) );
  GTECH_AND2 C25305 ( .A(N1051), .B(N583), .Z(N800) );
  GTECH_AND2 C25306 ( .A(N584), .B(byte_wen_d1[13]), .Z(N1051) );
  GTECH_NOT I_64 ( .A(N800), .Z(N801) );
  GTECH_AND2 C25309 ( .A(N1052), .B(N583), .Z(N803) );
  GTECH_AND2 C25310 ( .A(N585), .B(byte_wen_d1[13]), .Z(N1052) );
  GTECH_NOT I_65 ( .A(N803), .Z(N804) );
  GTECH_AND2 C25313 ( .A(N1053), .B(N583), .Z(N806) );
  GTECH_AND2 C25314 ( .A(N586), .B(byte_wen_d1[13]), .Z(N1053) );
  GTECH_NOT I_66 ( .A(N806), .Z(N807) );
  GTECH_AND2 C25317 ( .A(N1054), .B(N583), .Z(N813) );
  GTECH_AND2 C25318 ( .A(N582), .B(byte_wen_d1[14]), .Z(N1054) );
  GTECH_NOT I_67 ( .A(N813), .Z(N814) );
  GTECH_AND2 C25321 ( .A(N1055), .B(N583), .Z(N816) );
  GTECH_AND2 C25322 ( .A(N584), .B(byte_wen_d1[14]), .Z(N1055) );
  GTECH_NOT I_68 ( .A(N816), .Z(N817) );
  GTECH_AND2 C25325 ( .A(N1056), .B(N583), .Z(N819) );
  GTECH_AND2 C25326 ( .A(N585), .B(byte_wen_d1[14]), .Z(N1056) );
  GTECH_NOT I_69 ( .A(N819), .Z(N820) );
  GTECH_AND2 C25329 ( .A(N1057), .B(N583), .Z(N822) );
  GTECH_AND2 C25330 ( .A(N586), .B(byte_wen_d1[14]), .Z(N1057) );
  GTECH_NOT I_70 ( .A(N822), .Z(N823) );
  GTECH_AND2 C25333 ( .A(N1058), .B(N583), .Z(N829) );
  GTECH_AND2 C25334 ( .A(N582), .B(byte_wen_d1[15]), .Z(N1058) );
  GTECH_NOT I_71 ( .A(N829), .Z(N830) );
  GTECH_AND2 C25337 ( .A(N1059), .B(N583), .Z(N832) );
  GTECH_AND2 C25338 ( .A(N584), .B(byte_wen_d1[15]), .Z(N1059) );
  GTECH_NOT I_72 ( .A(N832), .Z(N833) );
  GTECH_AND2 C25341 ( .A(N1060), .B(N583), .Z(N835) );
  GTECH_AND2 C25342 ( .A(N585), .B(byte_wen_d1[15]), .Z(N1060) );
  GTECH_NOT I_73 ( .A(N835), .Z(N836) );
  GTECH_AND2 C25345 ( .A(N1061), .B(N583), .Z(N838) );
  GTECH_AND2 C25346 ( .A(N586), .B(byte_wen_d1[15]), .Z(N1061) );
  GTECH_NOT I_74 ( .A(N838), .Z(N839) );
  GTECH_AND2 C25349 ( .A(N1062), .B(N583), .Z(N845) );
  GTECH_AND2 C25350 ( .A(N582), .B(byte_wen_d1[16]), .Z(N1062) );
  GTECH_NOT I_75 ( .A(N845), .Z(N846) );
  GTECH_AND2 C25353 ( .A(N1063), .B(N583), .Z(N848) );
  GTECH_AND2 C25354 ( .A(N584), .B(byte_wen_d1[16]), .Z(N1063) );
  GTECH_NOT I_76 ( .A(N848), .Z(N849) );
  GTECH_AND2 C25357 ( .A(N1064), .B(N583), .Z(N851) );
  GTECH_AND2 C25358 ( .A(N585), .B(byte_wen_d1[16]), .Z(N1064) );
  GTECH_NOT I_77 ( .A(N851), .Z(N852) );
  GTECH_AND2 C25361 ( .A(N1065), .B(N583), .Z(N854) );
  GTECH_AND2 C25362 ( .A(N586), .B(byte_wen_d1[16]), .Z(N1065) );
  GTECH_NOT I_78 ( .A(N854), .Z(N855) );
  GTECH_AND2 C25365 ( .A(N1066), .B(N583), .Z(N861) );
  GTECH_AND2 C25366 ( .A(N582), .B(byte_wen_d1[17]), .Z(N1066) );
  GTECH_NOT I_79 ( .A(N861), .Z(N862) );
  GTECH_AND2 C25369 ( .A(N1067), .B(N583), .Z(N864) );
  GTECH_AND2 C25370 ( .A(N584), .B(byte_wen_d1[17]), .Z(N1067) );
  GTECH_NOT I_80 ( .A(N864), .Z(N865) );
  GTECH_AND2 C25373 ( .A(N1068), .B(N583), .Z(N867) );
  GTECH_AND2 C25374 ( .A(N585), .B(byte_wen_d1[17]), .Z(N1068) );
  GTECH_NOT I_81 ( .A(N867), .Z(N868) );
  GTECH_AND2 C25377 ( .A(N1069), .B(N583), .Z(N870) );
  GTECH_AND2 C25378 ( .A(N586), .B(byte_wen_d1[17]), .Z(N1069) );
  GTECH_NOT I_82 ( .A(N870), .Z(N871) );
  GTECH_AND2 C25381 ( .A(N1070), .B(N583), .Z(N877) );
  GTECH_AND2 C25382 ( .A(N582), .B(byte_wen_d1[18]), .Z(N1070) );
  GTECH_NOT I_83 ( .A(N877), .Z(N878) );
  GTECH_AND2 C25385 ( .A(N1071), .B(N583), .Z(N880) );
  GTECH_AND2 C25386 ( .A(N584), .B(byte_wen_d1[18]), .Z(N1071) );
  GTECH_NOT I_84 ( .A(N880), .Z(N881) );
  GTECH_AND2 C25389 ( .A(N1072), .B(N583), .Z(N883) );
  GTECH_AND2 C25390 ( .A(N585), .B(byte_wen_d1[18]), .Z(N1072) );
  GTECH_NOT I_85 ( .A(N883), .Z(N884) );
  GTECH_AND2 C25393 ( .A(N1073), .B(N583), .Z(N886) );
  GTECH_AND2 C25394 ( .A(N586), .B(byte_wen_d1[18]), .Z(N1073) );
  GTECH_NOT I_86 ( .A(N886), .Z(N887) );
  GTECH_AND2 C25397 ( .A(N1074), .B(N583), .Z(N893) );
  GTECH_AND2 C25398 ( .A(N582), .B(byte_wen_d1[19]), .Z(N1074) );
  GTECH_NOT I_87 ( .A(N893), .Z(N894) );
  GTECH_AND2 C25401 ( .A(N1075), .B(N583), .Z(N896) );
  GTECH_AND2 C25402 ( .A(N584), .B(byte_wen_d1[19]), .Z(N1075) );
  GTECH_NOT I_88 ( .A(N896), .Z(N897) );
  GTECH_AND2 C25405 ( .A(N1076), .B(N583), .Z(N899) );
  GTECH_AND2 C25406 ( .A(N585), .B(byte_wen_d1[19]), .Z(N1076) );
  GTECH_NOT I_89 ( .A(N899), .Z(N900) );
  GTECH_AND2 C25409 ( .A(N1077), .B(N583), .Z(N902) );
  GTECH_AND2 C25410 ( .A(N586), .B(byte_wen_d1[19]), .Z(N1077) );
  GTECH_NOT I_90 ( .A(N902), .Z(N903) );
  GTECH_NOT I_91 ( .A(sehold), .Z(N989) );
endmodule


module dffe_SIZE1 ( din, en, clk, q, se, si, so );
  input [0:0] din;
  output [0:0] q;
  input [0:0] si;
  output [0:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6;
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N6) );
  SELECT_OP C19 ( .DATA1(si[0]), .DATA2(din[0]), .CONTROL1(N0), .CONTROL2(N1), 
        .Z(N4) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C27 ( .A(N3), .B(N2), .Z(N5) );
  GTECH_NOT I_2 ( .A(N5), .Z(N6) );
endmodule


module dffre_SIZE8 ( din, rst, en, clk, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25;
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N25) );
  SELECT_OP C62 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(din), .CONTROL1(N0), .CONTROL2(N23), .Z({N13, N12, N11, N10, N9, 
        N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C63 ( .DATA1(si), .DATA2({N13, N12, N11, N10, N9, N8, N7, N6}), 
        .CONTROL1(N1), .CONTROL2(N2), .Z({N21, N20, N19, N18, N17, N16, N15, 
        N14}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C71 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N22) );
  GTECH_AND2 C74 ( .A(en), .B(N22), .Z(N23) );
  GTECH_AND2 C75 ( .A(N5), .B(N3), .Z(N24) );
  GTECH_NOT I_3 ( .A(N24), .Z(N25) );
endmodule


module dffe_SIZE4 ( din, en, clk, q, se, si, so );
  input [3:0] din;
  output [3:0] q;
  input [3:0] si;
  output [3:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N9) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N9) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N9) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N9) );
  SELECT_OP C31 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C39 ( .A(N3), .B(N2), .Z(N8) );
  GTECH_NOT I_2 ( .A(N8), .Z(N9) );
endmodule


module dffe_SIZE2 ( din, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7;
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N7) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N7) );
  SELECT_OP C23 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C31 ( .A(N3), .B(N2), .Z(N6) );
  GTECH_NOT I_2 ( .A(N6), .Z(N7) );
endmodule


module dffe_SIZE5 ( din, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10;
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N10) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N10) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N10) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N10) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N10) );
  SELECT_OP C35 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C43 ( .A(N3), .B(N2), .Z(N9) );
  GTECH_NOT I_2 ( .A(N9), .Z(N10) );
endmodule


module dffre_SIZE31 ( din, rst, en, clk, q, se, si, so );
  input [30:0] din;
  output [30:0] q;
  input [30:0] si;
  output [30:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71;
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N71) );
  SELECT_OP C177 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(din), .CONTROL1(N0), .CONTROL2(N69), .Z({N36, N35, N34, N33, 
        N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C178 ( .DATA1(si), .DATA2({N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6}), .CONTROL1(N1), .CONTROL2(N2), .Z({N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C186 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N68) );
  GTECH_AND2 C189 ( .A(en), .B(N68), .Z(N69) );
  GTECH_AND2 C190 ( .A(N5), .B(N3), .Z(N70) );
  GTECH_NOT I_3 ( .A(N70), .Z(N71) );
endmodule


module dffre_SIZE19 ( din, rst, en, clk, q, se, si, so );
  input [18:0] din;
  output [18:0] q;
  input [18:0] si;
  output [18:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47;
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N47) );
  SELECT_OP C117 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(din), .CONTROL1(N0), .CONTROL2(N45), .Z({N24, N23, N22, N21, 
        N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C118 ( .DATA1(si), .DATA2({N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}), .CONTROL1(N1), 
        .CONTROL2(N2), .Z({N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C126 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N44) );
  GTECH_AND2 C129 ( .A(en), .B(N44), .Z(N45) );
  GTECH_AND2 C130 ( .A(N5), .B(N3), .Z(N46) );
  GTECH_NOT I_3 ( .A(N46), .Z(N47) );
endmodule


module dffre_SIZE2 ( din, rst, en, clk, q, se, si, so );
  input [1:0] din;
  output [1:0] q;
  input [1:0] si;
  output [1:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13;
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N13) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N13) );
  SELECT_OP C32 ( .DATA1({1'b0, 1'b0}), .DATA2(din), .CONTROL1(N0), .CONTROL2(
        N11), .Z({N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C33 ( .DATA1(si), .DATA2({N7, N6}), .CONTROL1(N1), .CONTROL2(N2), 
        .Z({N9, N8}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C41 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N10) );
  GTECH_AND2 C44 ( .A(en), .B(N10), .Z(N11) );
  GTECH_AND2 C45 ( .A(N5), .B(N3), .Z(N12) );
  GTECH_NOT I_3 ( .A(N12), .Z(N13) );
endmodule


module dffre_SIZE18 ( din, rst, en, clk, q, se, si, so );
  input [17:0] din;
  output [17:0] q;
  input [17:0] si;
  output [17:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45;
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N45) );
  SELECT_OP C112 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(
        din), .CONTROL1(N0), .CONTROL2(N43), .Z({N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C113 ( .DATA1(si), .DATA2({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}), .CONTROL1(N1), 
        .CONTROL2(N2), .Z({N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C121 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N42) );
  GTECH_AND2 C124 ( .A(en), .B(N42), .Z(N43) );
  GTECH_AND2 C125 ( .A(N5), .B(N3), .Z(N44) );
  GTECH_NOT I_3 ( .A(N44), .Z(N45) );
endmodule


module dffe_SIZE10 ( din, en, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15;
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N15) );
  SELECT_OP C55 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C63 ( .A(N3), .B(N2), .Z(N14) );
  GTECH_NOT I_2 ( .A(N14), .Z(N15) );
endmodule


module dffre_SIZE9 ( din, rst, en, clk, q, se, si, so );
  input [8:0] din;
  output [8:0] q;
  input [8:0] si;
  output [8:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27;
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N27) );
  SELECT_OP C67 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(din), .CONTROL1(N0), .CONTROL2(N25), .Z({N14, N13, N12, N11, N10, N9, 
        N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C68 ( .DATA1(si), .DATA2({N14, N13, N12, N11, N10, N9, N8, N7, N6}), .CONTROL1(N1), .CONTROL2(N2), .Z({N23, N22, N21, N20, N19, N18, N17, N16, 
        N15}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C76 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N24) );
  GTECH_AND2 C79 ( .A(en), .B(N24), .Z(N25) );
  GTECH_AND2 C80 ( .A(N5), .B(N3), .Z(N26) );
  GTECH_NOT I_3 ( .A(N26), .Z(N27) );
endmodule


module dffre_SIZE6 ( din, rst, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21;
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N21) );
  SELECT_OP C52 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(din), 
        .CONTROL1(N0), .CONTROL2(N19), .Z({N11, N10, N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C53 ( .DATA1(si), .DATA2({N11, N10, N9, N8, N7, N6}), .CONTROL1(N1), .CONTROL2(N2), .Z({N17, N16, N15, N14, N13, N12}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C61 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N18) );
  GTECH_AND2 C64 ( .A(en), .B(N18), .Z(N19) );
  GTECH_AND2 C65 ( .A(N5), .B(N3), .Z(N20) );
  GTECH_NOT I_3 ( .A(N20), .Z(N21) );
endmodule


module dff_SIZE10 ( din, clk, q, se, si, so );
  input [9:0] din;
  output [9:0] q;
  input [9:0] si;
  output [9:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12;
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C20 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module fpu_add_ctl ( inq_in1_51, inq_in1_54, inq_in1_63, inq_in1_50_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_51, 
        inq_in2_54, inq_in2_63, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_op, inq_rnd_mode, inq_id, 
        inq_fcc, inq_add, add_dest_rdy, a1stg_in2_neq_in1_frac, 
        a1stg_in2_gt_in1_frac, a1stg_in2_eq_in1_exp, a1stg_expadd1, 
        a2stg_expadd, a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0, a2stg_exp, 
        a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a2stg_frac2_63, a4stg_exp, 
        add_of_out_cout, a4stg_frac_neq_0, a4stg_shl_data_neq_0, 
        a4stg_frac_dbl_nx, a4stg_frac_sng_nx, a1stg_expadd2, a1stg_expadd4_inv, 
        a3stg_denorm, a3stg_denorm_inv, a4stg_denorm_inv, a3stg_exp, 
        a4stg_round, a3stg_lead0, a4stg_rnd_frac_40, a4stg_rnd_frac_39, 
        a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_frac_38_0_nx, 
        a4stg_frac_9_0_nx, arst_l, grst_l, rclk, add_pipe_active, 
        a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1, a1stg_denorm_sng_in2, 
        a1stg_denorm_dbl_in2, a1stg_norm_sng_in1, a1stg_norm_dbl_in1, 
        a1stg_norm_sng_in2, a1stg_norm_dbl_in2, a1stg_step, a1stg_stepa, 
        a1stg_sngop, a1stg_intlngop, a1stg_fsdtoix, a1stg_fstod, a1stg_fstoi, 
        a1stg_fstox, a1stg_fdtoi, a1stg_fdtox, a1stg_faddsubs, a1stg_faddsubd, 
        a1stg_fdtos, a2stg_faddsubop, a2stg_fsdtoix_fdtos, a2stg_fitos, 
        a2stg_fitod, a2stg_fxtos, a2stg_fxtod, a3stg_faddsubop, 
        a3stg_faddsubopa, a4stg_dblop, a6stg_fadd_in, add_id_out_in, 
        add_fcc_out, a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, 
        a6stg_int_dst, a6stg_fcmpop, a6stg_step, a3stg_sub_in, add_sign_out, 
        add_cc_out, a4stg_in_of, add_exc_out, a2stg_frac1_in_frac1, 
        a2stg_frac1_in_frac2, a1stg_2nan_in_inv, a1stg_faddsubop_inv, 
        a2stg_frac1_in_qnan, a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, 
        a2stg_frac2_in_frac1, a2stg_frac2_in_qnan, a2stg_shr_cnt_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int, 
        a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max, 
        a2stg_sub_step, a2stg_fracadd_frac2_inv_in, 
        a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2, 
        a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add, 
        a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, 
        a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv, 
        a4stg_shl_cnt_in, a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0, 
        add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1, 
        add_exp_out_expadd, a4stg_to_0_inv, se, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [1:0] inq_fcc;
  input [11:0] a1stg_expadd1;
  input [11:0] a2stg_expadd;
  input [11:0] a2stg_exp;
  input [11:0] a4stg_exp;
  input [5:0] a1stg_expadd2;
  input [10:0] a1stg_expadd4_inv;
  input [10:0] a3stg_exp;
  input [5:0] a3stg_lead0;
  output [1:0] a3stg_faddsubopa;
  output [9:0] add_id_out_in;
  output [1:0] add_fcc_out;
  output [1:0] add_cc_out;
  output [4:0] add_exc_out;
  output [5:0] a2stg_shr_cnt_in;
  output [9:0] a4stg_shl_cnt_in;
  input inq_in1_51, inq_in1_54, inq_in1_63, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_63, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add,
         add_dest_rdy, a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac,
         a1stg_in2_eq_in1_exp, a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0,
         a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a2stg_frac2_63, add_of_out_cout,
         a4stg_frac_neq_0, a4stg_shl_data_neq_0, a4stg_frac_dbl_nx,
         a4stg_frac_sng_nx, a3stg_denorm, a3stg_denorm_inv, a4stg_denorm_inv,
         a4stg_round, a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac_11,
         a4stg_rnd_frac_10, a4stg_frac_38_0_nx, a4stg_frac_9_0_nx, arst_l,
         grst_l, rclk, se, si;
  output add_pipe_active, a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1,
         a1stg_denorm_sng_in2, a1stg_denorm_dbl_in2, a1stg_norm_sng_in1,
         a1stg_norm_dbl_in1, a1stg_norm_sng_in2, a1stg_norm_dbl_in2,
         a1stg_step, a1stg_stepa, a1stg_sngop, a1stg_intlngop, a1stg_fsdtoix,
         a1stg_fstod, a1stg_fstoi, a1stg_fstox, a1stg_fdtoi, a1stg_fdtox,
         a1stg_faddsubs, a1stg_faddsubd, a1stg_fdtos, a2stg_faddsubop,
         a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod, a2stg_fxtos,
         a2stg_fxtod, a3stg_faddsubop, a4stg_dblop, a6stg_fadd_in,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         a6stg_fcmpop, a6stg_step, a3stg_sub_in, add_sign_out, a4stg_in_of,
         a2stg_frac1_in_frac1, a2stg_frac1_in_frac2, a1stg_2nan_in_inv,
         a1stg_faddsubop_inv, a2stg_frac1_in_qnan, a2stg_frac1_in_nv,
         a2stg_frac1_in_nv_dbl, a2stg_frac2_in_frac1, a2stg_frac2_in_qnan,
         a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add,
         a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0,
         a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1,
         add_exp_out_expadd, a4stg_to_0_inv, so;
  wire   a1stg_step, add_exc_out_0, add_ctl_rst_l, reset, a1stg_in1_51,
         a1stg_in1_54, a1stg_in1_63, a1stg_in1_50_0_neq_0,
         a1stg_in1_53_32_neq_0, a1stg_in1_exp_eq_0, a1stg_in1_exp_neq_ffs,
         a1stg_in2_51, a1stg_in2_54, a1stg_in2_63, a1stg_in2_50_0_neq_0,
         a1stg_in2_53_32_neq_0, a1stg_in2_exp_eq_0, a1stg_in2_exp_neq_ffs,
         a1stg_snan_sng_in1, a1stg_snan_dbl_in1, a1stg_snan_sng_in2,
         a1stg_snan_dbl_in2, a1stg_qnan_sng_in1, a1stg_qnan_dbl_in1,
         a1stg_qnan_sng_in2, a1stg_qnan_dbl_in2, a1stg_snan_in1,
         a1stg_snan_in2, a1stg_qnan_in1, a1stg_qnan_in2, a1stg_nan_sng_in1,
         a1stg_nan_dbl_in1, a1stg_nan_sng_in2, a1stg_nan_dbl_in2,
         a1stg_nan_in1, a1stg_nan_in2, a1stg_nan_in, a1stg_2nan_in,
         a1stg_inf_sng_in1, a1stg_inf_dbl_in1, a1stg_inf_sng_in2,
         a1stg_inf_dbl_in2, a1stg_inf_in1, a1stg_inf_in2, a1stg_2inf_in,
         a1stg_infnan_sng_in1, a1stg_infnan_dbl_in1, a1stg_infnan_sng_in2,
         a1stg_infnan_dbl_in2, a1stg_infnan_in1, a1stg_infnan_in2,
         a1stg_infnan_in, a1stg_2zero_in, fixtosd_hold, a6stg_hold,
         a1stg_dblop, a1stg_fsdtox, a1stg_fcmpesd, a1stg_fcmpsd, a1stg_fixtosd,
         a1stg_opdec_9_0_2, a1stg_opdec_9_0_1, a2stg_opdec_36, a2stg_opdec_28,
         a3stg_opdec_36, a3stg_opdec_24, a3stg_fsdtoix, a4stg_faddsub_dtosop,
         a4stg_fsdtoix, a4stg_fcmpop, a5stg_opdec_9, a5stg_fixtos_fxtod,
         a5stg_fixtos, a5stg_fxtod, a6stg_opdec_in_9, N0, add_pipe_active_in,
         a1stg_sub, a2stg_sign1, a2stg_sign2, a2stg_sub,
         a2stg_in2_neq_in1_frac, a2stg_in2_gt_in1_frac, a2stg_in2_eq_in1_exp,
         a2stg_in2_gt_in1_exp, a2stg_nan_in, a2stg_nan_in2, a2stg_snan_in2,
         a2stg_qnan_in2, a2stg_snan_in1, a2stg_qnan_in1, a2stg_2zero_in,
         a2stg_2inf_in, a2stg_in2_eq_in1, a2stg_in2_gt_in1, N1, N2, N3, N4,
         a2stg_faddsub_sign, a3stg_sign_in, a3stg_sign, a4stg_sign2,
         a4stg_sign_in, a4stg_sign, a1stg_nv, a2stg_nv, a1stg_of_mask,
         a2stg_of_mask, a3stg_nv_in, a3stg_nv, a3stg_of_mask, a2stg_nx_tmp1,
         a2stg_nx_tmp2, a2stg_nx_tmp3, a3stg_a2_expadd_11, a3stg_nx_tmp1,
         a3stg_nx_tmp2, a3stg_nx_tmp3, a3stg_nx, N5, a4stg_nv2, a4stg_nv_in,
         a4stg_nv, N6, a4stg_of_mask2, a4stg_of_mask_in, a4stg_of_mask, N7,
         a4stg_nx2, a4stg_nx_in, a4stg_nx, a4stg_rndup, add_of_out_tmp1_in,
         add_of_out_tmp1, add_of_out_tmp2, N8, a4stg_uf, add_nx_out_in,
         add_nx_out, a1stg_exp_diff_add1, a1stg_exp_diff_add2,
         a1stg_exp_diff_5, a1stg_faddsub_clamp63_0, a2stg_fracadd_frac2_in, N9,
         a4stg_rndup_sng, a4stg_rndup_dbl, a5stg_rndup, N10, N11, N12, N13,
         N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285,
         N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296,
         N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307,
         N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318,
         N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329,
         N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340,
         N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351,
         N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362,
         N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384,
         N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417,
         N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450,
         N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483,
         N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516,
         N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
         N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538,
         N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604,
         N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648,
         N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714,
         N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725,
         N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901,
         N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020,
         N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030,
         N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040,
         N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050,
         N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060,
         N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070,
         N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080,
         N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090,
         N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100,
         N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110,
         N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120,
         N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130,
         N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140,
         N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150,
         N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160,
         N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170,
         N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180,
         N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190,
         N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200,
         N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210,
         N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220,
         N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230,
         N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240,
         N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250,
         N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260,
         N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270,
         N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280,
         N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290,
         N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300,
         N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310,
         N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320,
         N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330,
         N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340,
         N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350,
         N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370,
         N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380,
         N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390,
         N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400,
         N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410,
         N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420,
         N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430,
         N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440,
         N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470,
         N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480,
         N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490,
         N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500,
         N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510,
         N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, N1519, N1520,
         N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530,
         N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540,
         N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550,
         N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560,
         N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570,
         N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580,
         N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590,
         N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600,
         N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610,
         N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620,
         N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630,
         N1631, N1632, N1633, N1634, N1635, N1636, N1637, net16106, net16107,
         net16108, net16109, net16110, net16111, net16112, net16113, net16114,
         net16115, net16116, net16117, net16118, net16119, net16120, net16121,
         net16122, net16123, net16124, net16125, net16126, net16127, net16128,
         net16129, net16130, net16131, net16132, net16133, net16134, net16135,
         net16136, net16137, net16138, net16139, net16140, net16141, net16142,
         net16143, net16144, net16145, net16146, net16147, net16148, net16149,
         net16150, net16151, net16152, net16153, net16154, net16155, net16156,
         net16157, net16158, net16159, net16160, net16161, net16162, net16163,
         net16164, net16165, net16166, net16167, net16168, net16169, net16170,
         net16171, net16172, net16173, net16174, net16175, net16176, net16177,
         net16178, net16179, net16180, net16181, net16182, net16183, net16184,
         net16185, net16186, net16187, net16188, net16189, net16190, net16191,
         net16192, net16193, net16194, net16195, net16196, net16197, net16198,
         net16199, net16200, net16201, net16202, net16203, net16204, net16205,
         net16206, net16207, net16208, net16209, net16210, net16211, net16212,
         net16213, net16214, net16215, net16216, net16217, net16218, net16219,
         net16220, net16221, net16222, net16223, net16224, net16225, net16226,
         net16227, net16228, net16229, net16230, net16231, net16232, net16233,
         net16234, net16235, net16236, net16237, net16238, net16239, net16240,
         net16241, net16242, net16243, net16244, net16245, net16246, net16247,
         net16248, net16249, net16250, net16251, net16252, net16253, net16254,
         net16255, net16256, net16257, net16258, net16259, net16260, net16261,
         net16262, net16263, net16264, net16265, net16266, net16267, net16268,
         net16269, net16270, net16271, net16272, net16273, net16274, net16275,
         net16276, net16277, net16278, net16279, net16280, net16281, net16282,
         net16283, net16284, net16285, net16286, net16287, net16288, net16289,
         net16290, net16291, net16292, net16293, net16294, net16295, net16296,
         net16297, net16298, net16299, net16300, net16301, net16302, net16303,
         net16304, net16305, net16306, net16307, net16308, net16309, net16310,
         net16311, net16312, net16313, net16314, net16315, net16316, net16317,
         net16318, net16319, net16320, net16321, net16322, net16323, net16324,
         net16325, net16326, net16327, net16328, net16329, net16330, net16331,
         net16332, net16333, net16334, net16335;
  wire   [3:0] a1stg_sngopa;
  wire   [3:0] a1stg_dblopa;
  wire   [7:0] a1stg_op_in;
  wire   [7:0] a1stg_op;
  wire   [1:0] a1stg_rnd_mode;
  wire   [4:0] a1stg_id;
  wire   [1:0] a1stg_fcc;
  wire   [34:28] a1stg_opdec;
  wire   [3:1] a1stg_opdec_24_21;
  wire   [3:3] a1stg_opdec_19_11;
  wire   [9:6] a1stg_opdec_9_0;
  wire   [30:0] a2stg_opdec_in;
  wire   [34:30] a2stg_opdec;
  wire   [3:0] a2stg_opdec_24_21;
  wire   [8:4] a2stg_opdec_19_11;
  wire   [9:1] a2stg_opdec_9_0;
  wire   [1:0] a2stg_rnd_mode;
  wire   [4:0] a2stg_id;
  wire   [1:0] a2stg_fcc;
  wire   [34:30] a3stg_opdec;
  wire   [9:0] a3stg_opdec_9_0;
  wire   [1:0] a3stg_rnd_mode;
  wire   [4:0] a3stg_id;
  wire   [1:0] a3stg_fcc;
  wire   [34:29] a4stg_opdec;
  wire   [7:0] a4stg_opdec_7_0;
  wire   [1:0] a4stg_rnd_mode2;
  wire   [1:0] a4stg_rnd_mode_in;
  wire   [1:0] a4stg_rnd_mode;
  wire   [9:0] a4stg_id;
  wire   [1:0] a4stg_fcc;
  wire   [34:30] a5stg_opdec;
  wire   [9:0] a5stg_id;
  wire   [34:30] a6stg_opdec_in;
  wire   [34:34] a6stg_opdec;
  wire   [9:0] add_id_out;
  wire   [1:0] add_fcc_out_in;
  wire   [1:0] a2stg_cc;
  wire   [1:0] a3stg_cc;
  wire   [1:0] a4stg_cc;
  wire   [1:0] add_cc_out_in;
  wire   [10:0] a1stg_exp_diff;
  assign add_exc_out[1] = 1'b0;
  assign a1stg_stepa = a1stg_step;
  assign add_exc_out[0] = add_exc_out_0;
  assign a3stg_exp10_1_eq0 = N25;
  assign a3stg_exp10_0_eq0 = N53;
  assign a1stg_fstoi = N83;
  assign a1stg_fstox = N91;
  assign a1stg_fdtoi = N100;
  assign a1stg_fdtox = N108;
  assign a1stg_fstod = N168;
  assign a1stg_fdtos = N775;

  dffrl_async_SIZE1 dffrl_add_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(add_ctl_rst_l), .se(se), .si(net16335) );
  dffe_SIZE1 i_a1stg_in1_51 ( .din(inq_in1_51), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in1_51), .se(se), .si(net16334) );
  dffe_SIZE1 i_a1stg_in1_54 ( .din(inq_in1_54), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in1_54), .se(se), .si(net16333) );
  dffe_SIZE1 i_a1stg_in1_63 ( .din(inq_in1_63), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in1_63), .se(se), .si(net16332) );
  dffe_SIZE1 i_a1stg_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(a1stg_step), .clk(rclk), .q(a1stg_in1_50_0_neq_0), .se(se), .si(net16331) );
  dffe_SIZE1 i_a1stg_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        a1stg_step), .clk(rclk), .q(a1stg_in1_53_32_neq_0), .se(se), .si(
        net16330) );
  dffe_SIZE1 i_a1stg_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(a1stg_step), 
        .clk(rclk), .q(a1stg_in1_exp_eq_0), .se(se), .si(net16329) );
  dffe_SIZE1 i_a1stg_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        a1stg_step), .clk(rclk), .q(a1stg_in1_exp_neq_ffs), .se(se), .si(
        net16328) );
  dffe_SIZE1 i_a1stg_in2_51 ( .din(inq_in2_51), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in2_51), .se(se), .si(net16327) );
  dffe_SIZE1 i_a1stg_in2_54 ( .din(inq_in2_54), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in2_54), .se(se), .si(net16326) );
  dffe_SIZE1 i_a1stg_in2_63 ( .din(inq_in2_63), .en(a1stg_step), .clk(rclk), 
        .q(a1stg_in2_63), .se(se), .si(net16325) );
  dffe_SIZE1 i_a1stg_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(a1stg_step), .clk(rclk), .q(a1stg_in2_50_0_neq_0), .se(se), .si(net16324) );
  dffe_SIZE1 i_a1stg_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        a1stg_step), .clk(rclk), .q(a1stg_in2_53_32_neq_0), .se(se), .si(
        net16323) );
  dffe_SIZE1 i_a1stg_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(a1stg_step), 
        .clk(rclk), .q(a1stg_in2_exp_eq_0), .se(se), .si(net16322) );
  dffe_SIZE1 i_a1stg_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        a1stg_step), .clk(rclk), .q(a1stg_in2_exp_neq_ffs), .se(se), .si(
        net16321) );
  dffre_SIZE8 i_a1stg_op ( .din(a1stg_op_in), .rst(reset), .en(a1stg_step), 
        .clk(rclk), .q(a1stg_op), .se(se), .si({net16313, net16314, net16315, 
        net16316, net16317, net16318, net16319, net16320}) );
  dffe_SIZE1 i_a1stg_sngop ( .din(inq_op[0]), .en(a1stg_step), .clk(rclk), .q(
        a1stg_sngop), .se(se), .si(net16312) );
  dffe_SIZE4 i_a1stg_sngopa ( .din({inq_op[0], inq_op[0], inq_op[0], inq_op[0]}), .en(a1stg_step), .clk(rclk), .q(a1stg_sngopa), .se(se), .si({net16308, 
        net16309, net16310, net16311}) );
  dffe_SIZE1 i_a1stg_dblop ( .din(inq_op[1]), .en(a1stg_step), .clk(rclk), .q(
        a1stg_dblop), .se(se), .si(net16307) );
  dffe_SIZE4 i_a1stg_dblopa ( .din({inq_op[1], inq_op[1], inq_op[1], inq_op[1]}), .en(a1stg_step), .clk(rclk), .q(a1stg_dblopa), .se(se), .si({net16303, 
        net16304, net16305, net16306}) );
  dffe_SIZE2 i_a1stg_rnd_mode ( .din(inq_rnd_mode), .en(a1stg_step), .clk(rclk), .q(a1stg_rnd_mode), .se(se), .si({net16301, net16302}) );
  dffe_SIZE5 i_a1stg_id ( .din(inq_id), .en(a1stg_step), .clk(rclk), .q(
        a1stg_id), .se(se), .si({net16296, net16297, net16298, net16299, 
        net16300}) );
  dffe_SIZE2 i_a1stg_fcc ( .din(inq_fcc), .en(a1stg_step), .clk(rclk), .q(
        a1stg_fcc), .se(se), .si({net16294, net16295}) );
  dffre_SIZE31 i_a2stg_opdec ( .din(a2stg_opdec_in), .rst(reset), .en(
        a6stg_step), .clk(rclk), .q({a2stg_opdec_36, a2stg_opdec, 
        a2stg_faddsubop, a2stg_opdec_28, a2stg_opdec_24_21, a2stg_opdec_19_11, 
        a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod, a2stg_fxtos, 
        a2stg_opdec_9_0, a2stg_fxtod}), .se(se), .si({net16263, net16264, 
        net16265, net16266, net16267, net16268, net16269, net16270, net16271, 
        net16272, net16273, net16274, net16275, net16276, net16277, net16278, 
        net16279, net16280, net16281, net16282, net16283, net16284, net16285, 
        net16286, net16287, net16288, net16289, net16290, net16291, net16292, 
        net16293}) );
  dffe_SIZE2 i_a2stg_rnd_mode ( .din(a1stg_rnd_mode), .en(a6stg_step), .clk(
        rclk), .q(a2stg_rnd_mode), .se(se), .si({net16261, net16262}) );
  dffe_SIZE5 i_a2stg_id ( .din(a1stg_id), .en(a6stg_step), .clk(rclk), .q(
        a2stg_id), .se(se), .si({net16256, net16257, net16258, net16259, 
        net16260}) );
  dffe_SIZE2 i_a2stg_fcc ( .din(a1stg_fcc), .en(a6stg_step), .clk(rclk), .q(
        a2stg_fcc), .se(se), .si({net16254, net16255}) );
  dffre_SIZE19 i_a3stg_opdec ( .din({a2stg_opdec_36, a2stg_opdec, 
        a2stg_faddsubop, a2stg_opdec_24_21[3], a2stg_opdec_24_21[0], 
        a2stg_opdec_9_0, a2stg_fxtod}), .rst(reset), .en(a6stg_step), .clk(
        rclk), .q({a3stg_opdec_36, a3stg_opdec, a3stg_faddsubop, 
        a3stg_opdec_24, a3stg_fsdtoix, a3stg_opdec_9_0}), .se(se), .si({
        net16235, net16236, net16237, net16238, net16239, net16240, net16241, 
        net16242, net16243, net16244, net16245, net16246, net16247, net16248, 
        net16249, net16250, net16251, net16252, net16253}) );
  dffre_SIZE2 i_a3stg_faddsubopa ( .din({a2stg_faddsubop, a2stg_faddsubop}), 
        .rst(reset), .en(a6stg_step), .clk(rclk), .q(a3stg_faddsubopa), .se(se), .si({net16233, net16234}) );
  dffe_SIZE2 i_a3stg_rnd_mode ( .din(a2stg_rnd_mode), .en(a6stg_step), .clk(
        rclk), .q(a3stg_rnd_mode), .se(se), .si({net16231, net16232}) );
  dffe_SIZE5 i_a3stg_id ( .din(a2stg_id), .en(a6stg_step), .clk(rclk), .q(
        a3stg_id), .se(se), .si({net16226, net16227, net16228, net16229, 
        net16230}) );
  dffe_SIZE2 i_a3stg_fcc ( .din(a2stg_fcc), .en(a6stg_step), .clk(rclk), .q(
        a3stg_fcc), .se(se), .si({net16224, net16225}) );
  dffre_SIZE18 i_a4stg_opdec ( .din({a3stg_opdec_36, a3stg_opdec, 
        a3stg_faddsubop, a3stg_opdec_24, a3stg_fsdtoix, a3stg_opdec_9_0[9], 
        a3stg_opdec_9_0[7:0]}), .rst(reset), .en(a6stg_step), .clk(rclk), .q({
        a4stg_dblop, a4stg_opdec, a4stg_faddsub_dtosop, a4stg_fsdtoix, 
        a4stg_fcmpop, a4stg_opdec_7_0}), .se(se), .si({net16206, net16207, 
        net16208, net16209, net16210, net16211, net16212, net16213, net16214, 
        net16215, net16216, net16217, net16218, net16219, net16220, net16221, 
        net16222, net16223}) );
  dffe_SIZE2 i_a4stg_rnd_mode ( .din(a4stg_rnd_mode_in), .en(a6stg_step), 
        .clk(rclk), .q(a4stg_rnd_mode), .se(se), .si({net16204, net16205}) );
  dffe_SIZE2 i_a4stg_rnd_mode2 ( .din(a3stg_rnd_mode), .en(a6stg_step), .clk(
        rclk), .q(a4stg_rnd_mode2), .se(se), .si({net16202, net16203}) );
  dffe_SIZE10 i_a4stg_id ( .din({N27, N32, N36, N39, N42, N45, N48, N51, 
        a3stg_id[1:0]}), .en(a6stg_step), .clk(rclk), .q(a4stg_id), .se(se), 
        .si({net16192, net16193, net16194, net16195, net16196, net16197, 
        net16198, net16199, net16200, net16201}) );
  dffe_SIZE2 i_a4stg_fcc ( .din(a3stg_fcc), .en(a6stg_step), .clk(rclk), .q(
        a4stg_fcc), .se(se), .si({net16190, net16191}) );
  dffre_SIZE9 i_a5stg_opdec ( .din({a4stg_opdec[34:30], a4stg_fcmpop, 
        a4stg_opdec_7_0[7], a4stg_opdec_7_0[1:0]}), .rst(reset), .en(
        a6stg_step), .clk(rclk), .q({a5stg_opdec, a5stg_opdec_9, 
        a5stg_fixtos_fxtod, a5stg_fixtos, a5stg_fxtod}), .se(se), .si({
        net16181, net16182, net16183, net16184, net16185, net16186, net16187, 
        net16188, net16189}) );
  dffe_SIZE10 i_a5stg_id ( .din(a4stg_id), .en(a6stg_step), .clk(rclk), .q(
        a5stg_id), .se(se), .si({net16171, net16172, net16173, net16174, 
        net16175, net16176, net16177, net16178, net16179, net16180}) );
  dffre_SIZE6 i_a6stg_opdec ( .din({a6stg_opdec_in, a6stg_opdec_in_9}), .rst(
        reset), .en(a6stg_step), .clk(rclk), .q({a6stg_opdec[34], 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        a6stg_fcmpop}), .se(se), .si({net16165, net16166, net16167, net16168, 
        net16169, net16170}) );
  dff_SIZE10 i_add_id_out ( .din(add_id_out_in), .clk(rclk), .q(add_id_out), 
        .se(se), .si({net16155, net16156, net16157, net16158, net16159, 
        net16160, net16161, net16162, net16163, net16164}) );
  dffe_SIZE2 i_add_fcc_out ( .din(add_fcc_out_in), .en(a6stg_step), .clk(rclk), 
        .q(add_fcc_out), .se(se), .si({net16153, net16154}) );
  dffre_SIZE1 i_add_pipe_active ( .din(add_pipe_active_in), .rst(reset), .en(
        1'b1), .clk(rclk), .q(add_pipe_active), .se(se), .si(net16152) );
  dffe_SIZE1 i_a2stg_sign1 ( .din(a1stg_in1_63), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_sign1), .se(se), .si(net16151) );
  dffe_SIZE1 i_a2stg_sign2 ( .din(a1stg_in2_63), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_sign2), .se(se), .si(net16150) );
  dffe_SIZE1 i_a2stg_sub ( .din(a1stg_sub), .en(a6stg_step), .clk(rclk), .q(
        a2stg_sub), .se(se), .si(net16149) );
  dffe_SIZE1 i_a2stg_in2_neq_in1_frac ( .din(a1stg_in2_neq_in1_frac), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_neq_in1_frac), .se(se), .si(
        net16148) );
  dffe_SIZE1 i_a2stg_in2_gt_in1_frac ( .din(a1stg_in2_gt_in1_frac), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_gt_in1_frac), .se(se), .si(
        net16147) );
  dffe_SIZE1 i_a2stg_in2_eq_in1_exp ( .din(a1stg_in2_eq_in1_exp), .en(
        a6stg_step), .clk(rclk), .q(a2stg_in2_eq_in1_exp), .se(se), .si(
        net16146) );
  dffe_SIZE1 i_a2stg_in2_gt_in1_exp ( .din(a1stg_expadd1[11]), .en(a6stg_step), 
        .clk(rclk), .q(a2stg_in2_gt_in1_exp), .se(se), .si(net16145) );
  dffe_SIZE1 i_a2stg_nan_in ( .din(a1stg_nan_in), .en(a6stg_step), .clk(rclk), 
        .q(a2stg_nan_in), .se(se), .si(net16144) );
  dffe_SIZE1 i_a2stg_nan_in2 ( .din(a1stg_nan_in2), .en(a6stg_step), .clk(rclk), .q(a2stg_nan_in2), .se(se), .si(net16143) );
  dffe_SIZE1 i_a2stg_snan_in2 ( .din(a1stg_snan_in2), .en(a6stg_step), .clk(
        rclk), .q(a2stg_snan_in2), .se(se), .si(net16142) );
  dffe_SIZE1 i_a2stg_qnan_in2 ( .din(a1stg_qnan_in2), .en(a6stg_step), .clk(
        rclk), .q(a2stg_qnan_in2), .se(se), .si(net16141) );
  dffe_SIZE1 i_a2stg_snan_in1 ( .din(a1stg_snan_in1), .en(a6stg_step), .clk(
        rclk), .q(a2stg_snan_in1), .se(se), .si(net16140) );
  dffe_SIZE1 i_a2stg_qnan_in1 ( .din(a1stg_qnan_in1), .en(a6stg_step), .clk(
        rclk), .q(a2stg_qnan_in1), .se(se), .si(net16139) );
  dffe_SIZE1 i_a2stg_2zero_in ( .din(a1stg_2zero_in), .en(a6stg_step), .clk(
        rclk), .q(a2stg_2zero_in), .se(se), .si(net16138) );
  dffe_SIZE1 i_a2stg_2inf_in ( .din(a1stg_2inf_in), .en(a6stg_step), .clk(rclk), .q(a2stg_2inf_in), .se(se), .si(net16137) );
  dffe_SIZE1 i_a3stg_sign ( .din(a3stg_sign_in), .en(a6stg_step), .clk(rclk), 
        .q(a3stg_sign), .se(se), .si(net16136) );
  dffe_SIZE2 i_a3stg_cc ( .din(a2stg_cc), .en(a6stg_step), .clk(rclk), .q(
        a3stg_cc), .se(se), .si({net16134, net16135}) );
  dffe_SIZE1 i_a4stg_sign ( .din(a4stg_sign_in), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_sign), .se(se), .si(net16133) );
  dffe_SIZE1 i_a4stg_sign2 ( .din(a3stg_sign), .en(a6stg_step), .clk(rclk), 
        .q(a4stg_sign2), .se(se), .si(net16132) );
  dffe_SIZE2 i_a4stg_cc ( .din(a3stg_cc), .en(a6stg_step), .clk(rclk), .q(
        a4stg_cc), .se(se), .si({net16130, net16131}) );
  dffe_SIZE1 i_add_sign_out ( .din(a4stg_sign), .en(a6stg_step), .clk(rclk), 
        .q(add_sign_out), .se(se), .si(net16129) );
  dffe_SIZE2 i_add_cc_out ( .din(add_cc_out_in), .en(a6stg_step), .clk(rclk), 
        .q(add_cc_out), .se(se), .si({net16127, net16128}) );
  dffe_SIZE1 i_a2stg_nv ( .din(a1stg_nv), .en(a6stg_step), .clk(rclk), .q(
        a2stg_nv), .se(se), .si(net16126) );
  dffe_SIZE1 i_a2stg_of_mask ( .din(a1stg_of_mask), .en(a6stg_step), .clk(rclk), .q(a2stg_of_mask), .se(se), .si(net16125) );
  dffe_SIZE1 i_a3stg_nv ( .din(a3stg_nv_in), .en(a6stg_step), .clk(rclk), .q(
        a3stg_nv), .se(se), .si(net16124) );
  dffe_SIZE1 i_a3stg_of_mask ( .din(a2stg_of_mask), .en(a6stg_step), .clk(rclk), .q(a3stg_of_mask), .se(se), .si(net16123) );
  dffe_SIZE1 i_a3stg_a2_expadd_11 ( .din(a2stg_expadd[11]), .en(a6stg_step), 
        .clk(rclk), .q(a3stg_a2_expadd_11), .se(se), .si(net16122) );
  dffe_SIZE1 i_a3stg_nx_tmp1 ( .din(a2stg_nx_tmp1), .en(a6stg_step), .clk(rclk), .q(a3stg_nx_tmp1), .se(se), .si(net16121) );
  dffe_SIZE1 i_a3stg_nx_tmp2 ( .din(a2stg_nx_tmp2), .en(a6stg_step), .clk(rclk), .q(a3stg_nx_tmp2), .se(se), .si(net16120) );
  dffe_SIZE1 i_a3stg_nx_tmp3 ( .din(a2stg_nx_tmp3), .en(a6stg_step), .clk(rclk), .q(a3stg_nx_tmp3), .se(se), .si(net16119) );
  dffe_SIZE1 i_a4stg_nv ( .din(a4stg_nv_in), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nv), .se(se), .si(net16118) );
  dffe_SIZE1 i_a4stg_nv2 ( .din(a3stg_nv), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nv2), .se(se), .si(net16117) );
  dffe_SIZE1 i_a4stg_of_mask ( .din(a4stg_of_mask_in), .en(a6stg_step), .clk(
        rclk), .q(a4stg_of_mask), .se(se), .si(net16116) );
  dffe_SIZE1 i_a4stg_of_mask2 ( .din(a3stg_of_mask), .en(a6stg_step), .clk(
        rclk), .q(a4stg_of_mask2), .se(se), .si(net16115) );
  dffe_SIZE1 i_a4stg_nx ( .din(a4stg_nx_in), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nx), .se(se), .si(net16114) );
  dffe_SIZE1 i_a4stg_nx2 ( .din(a3stg_nx), .en(a6stg_step), .clk(rclk), .q(
        a4stg_nx2), .se(se), .si(net16113) );
  dffe_SIZE1 i_add_nv_out ( .din(a4stg_nv), .en(a6stg_step), .clk(rclk), .q(
        add_exc_out[4]), .se(se), .si(net16112) );
  dffe_SIZE1 i_add_of_out_tmp1 ( .din(add_of_out_tmp1_in), .en(a6stg_step), 
        .clk(rclk), .q(add_of_out_tmp1), .se(se), .si(net16111) );
  dffe_SIZE1 i_add_of_out_tmp2 ( .din(a4stg_in_of), .en(a6stg_step), .clk(rclk), .q(add_of_out_tmp2), .se(se), .si(net16110) );
  dffe_SIZE1 i_add_uf_out ( .din(a4stg_uf), .en(a6stg_step), .clk(rclk), .q(
        add_exc_out[2]), .se(se), .si(net16109) );
  dffe_SIZE1 i_add_nx_out ( .din(add_nx_out_in), .en(a6stg_step), .clk(rclk), 
        .q(add_nx_out), .se(se), .si(net16108) );
  dffe_SIZE1 i_a2stg_fracadd_frac2 ( .din(a2stg_fracadd_frac2_in), .en(
        a6stg_step), .clk(rclk), .q(a2stg_fracadd_frac2), .se(se), .si(
        net16107) );
  LT_UNS_OP lt_2599 ( .A(a2stg_exp[10:0]), .B({1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 
        1'b0}), .Z(N9) );
  GTECH_OR2 C255 ( .A(a3stg_exp[9]), .B(a3stg_exp[10]), .Z(N16) );
  GTECH_OR2 C256 ( .A(a3stg_exp[8]), .B(N16), .Z(N17) );
  GTECH_OR2 C257 ( .A(a3stg_exp[7]), .B(N17), .Z(N18) );
  GTECH_OR2 C258 ( .A(a3stg_exp[6]), .B(N18), .Z(N19) );
  GTECH_OR2 C259 ( .A(a3stg_exp[5]), .B(N19), .Z(N20) );
  GTECH_OR2 C260 ( .A(a3stg_exp[4]), .B(N20), .Z(N21) );
  GTECH_OR2 C261 ( .A(a3stg_exp[3]), .B(N21), .Z(N22) );
  GTECH_OR2 C262 ( .A(a3stg_exp[2]), .B(N22), .Z(N23) );
  GTECH_OR2 C263 ( .A(a3stg_exp[1]), .B(N23), .Z(N24) );
  GTECH_NOT I_0 ( .A(N24), .Z(N25) );
  GTECH_AND2 C265 ( .A(a3stg_id[3]), .B(a3stg_id[4]), .Z(N26) );
  GTECH_AND2 C266 ( .A(a3stg_id[2]), .B(N26), .Z(N27) );
  GTECH_NOT I_1 ( .A(a3stg_id[4]), .Z(N28) );
  GTECH_NOT I_2 ( .A(a3stg_id[3]), .Z(N29) );
  GTECH_OR2 C269 ( .A(N29), .B(N28), .Z(N30) );
  GTECH_OR2 C270 ( .A(a3stg_id[2]), .B(N30), .Z(N31) );
  GTECH_NOT I_3 ( .A(N31), .Z(N32) );
  GTECH_NOT I_4 ( .A(a3stg_id[2]), .Z(N33) );
  GTECH_OR2 C274 ( .A(a3stg_id[3]), .B(N28), .Z(N34) );
  GTECH_OR2 C275 ( .A(N33), .B(N34), .Z(N35) );
  GTECH_NOT I_5 ( .A(N35), .Z(N36) );
  GTECH_OR2 C278 ( .A(a3stg_id[3]), .B(N28), .Z(N37) );
  GTECH_OR2 C279 ( .A(a3stg_id[2]), .B(N37), .Z(N38) );
  GTECH_NOT I_6 ( .A(N38), .Z(N39) );
  GTECH_OR2 C283 ( .A(N29), .B(a3stg_id[4]), .Z(N40) );
  GTECH_OR2 C284 ( .A(N33), .B(N40), .Z(N41) );
  GTECH_NOT I_7 ( .A(N41), .Z(N42) );
  GTECH_OR2 C287 ( .A(N29), .B(a3stg_id[4]), .Z(N43) );
  GTECH_OR2 C288 ( .A(a3stg_id[2]), .B(N43), .Z(N44) );
  GTECH_NOT I_8 ( .A(N44), .Z(N45) );
  GTECH_OR2 C291 ( .A(a3stg_id[3]), .B(a3stg_id[4]), .Z(N46) );
  GTECH_OR2 C292 ( .A(N33), .B(N46), .Z(N47) );
  GTECH_NOT I_9 ( .A(N47), .Z(N48) );
  GTECH_OR2 C294 ( .A(a3stg_id[3]), .B(a3stg_id[4]), .Z(N49) );
  GTECH_OR2 C295 ( .A(a3stg_id[2]), .B(N49), .Z(N50) );
  GTECH_NOT I_10 ( .A(N50), .Z(N51) );
  GTECH_OR2 C306 ( .A(a3stg_exp[0]), .B(N24), .Z(N52) );
  GTECH_NOT I_11 ( .A(N52), .Z(N53) );
  GTECH_AND2 C308 ( .A(a3stg_exp[4]), .B(a3stg_exp[5]), .Z(N54) );
  GTECH_AND2 C309 ( .A(a3stg_lead0[4]), .B(a3stg_lead0[5]), .Z(N55) );
  GTECH_NOT I_12 ( .A(a3stg_exp[5]), .Z(N56) );
  GTECH_OR2 C311 ( .A(a3stg_exp[4]), .B(N56), .Z(N57) );
  GTECH_NOT I_13 ( .A(N57), .Z(N58) );
  GTECH_NOT I_14 ( .A(a3stg_lead0[5]), .Z(N59) );
  GTECH_OR2 C314 ( .A(a3stg_lead0[4]), .B(N59), .Z(N60) );
  GTECH_NOT I_15 ( .A(N60), .Z(N61) );
  GTECH_NOT I_16 ( .A(a3stg_exp[4]), .Z(N62) );
  GTECH_OR2 C317 ( .A(N62), .B(a3stg_exp[5]), .Z(N63) );
  GTECH_NOT I_17 ( .A(N63), .Z(N64) );
  GTECH_NOT I_18 ( .A(a3stg_lead0[4]), .Z(N65) );
  GTECH_OR2 C320 ( .A(N65), .B(a3stg_lead0[5]), .Z(N66) );
  GTECH_NOT I_19 ( .A(N66), .Z(N67) );
  GTECH_OR2 C322 ( .A(a3stg_exp[4]), .B(a3stg_exp[5]), .Z(N68) );
  GTECH_NOT I_20 ( .A(N68), .Z(N69) );
  GTECH_OR2 C324 ( .A(a3stg_lead0[4]), .B(a3stg_lead0[5]), .Z(N70) );
  GTECH_NOT I_21 ( .A(N70), .Z(N71) );
  GTECH_NOT I_22 ( .A(a1stg_op[7]), .Z(N72) );
  GTECH_NOT I_23 ( .A(a1stg_op[6]), .Z(N73) );
  GTECH_NOT I_24 ( .A(a1stg_op[4]), .Z(N74) );
  GTECH_NOT I_25 ( .A(a1stg_op[0]), .Z(N75) );
  GTECH_OR2 C330 ( .A(N73), .B(N72), .Z(N76) );
  GTECH_OR2 C331 ( .A(a1stg_op[5]), .B(N76), .Z(N77) );
  GTECH_OR2 C332 ( .A(N74), .B(N77), .Z(N78) );
  GTECH_OR2 C333 ( .A(a1stg_op[3]), .B(N78), .Z(N79) );
  GTECH_OR2 C334 ( .A(a1stg_op[2]), .B(N79), .Z(N80) );
  GTECH_OR2 C335 ( .A(a1stg_op[1]), .B(N80), .Z(N81) );
  GTECH_OR2 C336 ( .A(N75), .B(N81), .Z(N82) );
  GTECH_NOT I_26 ( .A(N82), .Z(N83) );
  GTECH_OR2 C340 ( .A(a1stg_op[6]), .B(N72), .Z(N84) );
  GTECH_OR2 C341 ( .A(a1stg_op[5]), .B(N84), .Z(N85) );
  GTECH_OR2 C342 ( .A(a1stg_op[4]), .B(N85), .Z(N86) );
  GTECH_OR2 C343 ( .A(a1stg_op[3]), .B(N86), .Z(N87) );
  GTECH_OR2 C344 ( .A(a1stg_op[2]), .B(N87), .Z(N88) );
  GTECH_OR2 C345 ( .A(a1stg_op[1]), .B(N88), .Z(N89) );
  GTECH_OR2 C346 ( .A(N75), .B(N89), .Z(N90) );
  GTECH_NOT I_27 ( .A(N90), .Z(N91) );
  GTECH_NOT I_28 ( .A(a1stg_op[1]), .Z(N92) );
  GTECH_OR2 C352 ( .A(N73), .B(N72), .Z(N93) );
  GTECH_OR2 C353 ( .A(a1stg_op[5]), .B(N93), .Z(N94) );
  GTECH_OR2 C354 ( .A(N74), .B(N94), .Z(N95) );
  GTECH_OR2 C355 ( .A(a1stg_op[3]), .B(N95), .Z(N96) );
  GTECH_OR2 C356 ( .A(a1stg_op[2]), .B(N96), .Z(N97) );
  GTECH_OR2 C357 ( .A(N92), .B(N97), .Z(N98) );
  GTECH_OR2 C358 ( .A(a1stg_op[0]), .B(N98), .Z(N99) );
  GTECH_NOT I_29 ( .A(N99), .Z(N100) );
  GTECH_OR2 C362 ( .A(a1stg_op[6]), .B(N72), .Z(N101) );
  GTECH_OR2 C363 ( .A(a1stg_op[5]), .B(N101), .Z(N102) );
  GTECH_OR2 C364 ( .A(a1stg_op[4]), .B(N102), .Z(N103) );
  GTECH_OR2 C365 ( .A(a1stg_op[3]), .B(N103), .Z(N104) );
  GTECH_OR2 C366 ( .A(a1stg_op[2]), .B(N104), .Z(N105) );
  GTECH_OR2 C367 ( .A(N92), .B(N105), .Z(N106) );
  GTECH_OR2 C368 ( .A(a1stg_op[0]), .B(N106), .Z(N107) );
  GTECH_NOT I_30 ( .A(N107), .Z(N108) );
  GTECH_NOT I_31 ( .A(a1stg_op[2]), .Z(N109) );
  GTECH_OR2 C373 ( .A(N73), .B(N72), .Z(N110) );
  GTECH_OR2 C374 ( .A(a1stg_op[5]), .B(N110), .Z(N111) );
  GTECH_OR2 C375 ( .A(a1stg_op[4]), .B(N111), .Z(N112) );
  GTECH_OR2 C376 ( .A(a1stg_op[3]), .B(N112), .Z(N113) );
  GTECH_OR2 C377 ( .A(N109), .B(N113), .Z(N114) );
  GTECH_OR2 C378 ( .A(a1stg_op[1]), .B(N114), .Z(N115) );
  GTECH_OR2 C379 ( .A(a1stg_op[0]), .B(N115), .Z(N116) );
  GTECH_NOT I_32 ( .A(N116), .Z(N117) );
  GTECH_NOT I_33 ( .A(a1stg_op[3]), .Z(N118) );
  GTECH_OR2 C384 ( .A(N73), .B(N72), .Z(N119) );
  GTECH_OR2 C385 ( .A(a1stg_op[5]), .B(N119), .Z(N120) );
  GTECH_OR2 C386 ( .A(a1stg_op[4]), .B(N120), .Z(N121) );
  GTECH_OR2 C387 ( .A(N118), .B(N121), .Z(N122) );
  GTECH_OR2 C388 ( .A(a1stg_op[2]), .B(N122), .Z(N123) );
  GTECH_OR2 C389 ( .A(a1stg_op[1]), .B(N123), .Z(N124) );
  GTECH_OR2 C390 ( .A(a1stg_op[0]), .B(N124), .Z(N125) );
  GTECH_NOT I_34 ( .A(N125), .Z(N126) );
  GTECH_OR2 C394 ( .A(a1stg_op[6]), .B(N72), .Z(N127) );
  GTECH_OR2 C395 ( .A(a1stg_op[5]), .B(N127), .Z(N128) );
  GTECH_OR2 C396 ( .A(a1stg_op[4]), .B(N128), .Z(N129) );
  GTECH_OR2 C397 ( .A(a1stg_op[3]), .B(N129), .Z(N130) );
  GTECH_OR2 C398 ( .A(N109), .B(N130), .Z(N131) );
  GTECH_OR2 C399 ( .A(a1stg_op[1]), .B(N131), .Z(N132) );
  GTECH_OR2 C400 ( .A(a1stg_op[0]), .B(N132), .Z(N133) );
  GTECH_NOT I_35 ( .A(N133), .Z(N134) );
  GTECH_OR2 C404 ( .A(a1stg_op[6]), .B(N72), .Z(N135) );
  GTECH_OR2 C405 ( .A(a1stg_op[5]), .B(N135), .Z(N136) );
  GTECH_OR2 C406 ( .A(a1stg_op[4]), .B(N136), .Z(N137) );
  GTECH_OR2 C407 ( .A(N118), .B(N137), .Z(N138) );
  GTECH_OR2 C408 ( .A(a1stg_op[2]), .B(N138), .Z(N139) );
  GTECH_OR2 C409 ( .A(a1stg_op[1]), .B(N139), .Z(N140) );
  GTECH_OR2 C410 ( .A(a1stg_op[0]), .B(N140), .Z(N141) );
  GTECH_NOT I_36 ( .A(N141), .Z(N142) );
  GTECH_NOT I_37 ( .A(a2stg_exp[10]), .Z(N143) );
  GTECH_NOT I_38 ( .A(a2stg_exp[4]), .Z(N144) );
  GTECH_NOT I_39 ( .A(a2stg_exp[3]), .Z(N145) );
  GTECH_NOT I_40 ( .A(a2stg_exp[2]), .Z(N146) );
  GTECH_NOT I_41 ( .A(a2stg_exp[1]), .Z(N147) );
  GTECH_NOT I_42 ( .A(a2stg_exp[0]), .Z(N148) );
  GTECH_OR2 C418 ( .A(N143), .B(a2stg_exp[11]), .Z(N149) );
  GTECH_OR2 C419 ( .A(a2stg_exp[9]), .B(N149), .Z(N150) );
  GTECH_OR2 C420 ( .A(a2stg_exp[8]), .B(N150), .Z(N151) );
  GTECH_OR2 C421 ( .A(a2stg_exp[7]), .B(N151), .Z(N152) );
  GTECH_OR2 C422 ( .A(a2stg_exp[6]), .B(N152), .Z(N153) );
  GTECH_OR2 C423 ( .A(a2stg_exp[5]), .B(N153), .Z(N154) );
  GTECH_OR2 C424 ( .A(N144), .B(N154), .Z(N155) );
  GTECH_OR2 C425 ( .A(N145), .B(N155), .Z(N156) );
  GTECH_OR2 C426 ( .A(N146), .B(N156), .Z(N157) );
  GTECH_OR2 C427 ( .A(N147), .B(N157), .Z(N158) );
  GTECH_OR2 C428 ( .A(N148), .B(N158), .Z(N159) );
  GTECH_NOT I_43 ( .A(N159), .Z(N160) );
  GTECH_OR2 C434 ( .A(N73), .B(N72), .Z(N161) );
  GTECH_OR2 C435 ( .A(a1stg_op[5]), .B(N161), .Z(N162) );
  GTECH_OR2 C436 ( .A(a1stg_op[4]), .B(N162), .Z(N163) );
  GTECH_OR2 C437 ( .A(N118), .B(N163), .Z(N164) );
  GTECH_OR2 C438 ( .A(a1stg_op[2]), .B(N164), .Z(N165) );
  GTECH_OR2 C439 ( .A(a1stg_op[1]), .B(N165), .Z(N166) );
  GTECH_OR2 C440 ( .A(N75), .B(N166), .Z(N167) );
  GTECH_NOT I_44 ( .A(N167), .Z(N168) );
  GTECH_OR2 C442 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N169) );
  GTECH_NOT I_45 ( .A(N169), .Z(N170) );
  GTECH_NOT I_46 ( .A(a4stg_rnd_mode[1]), .Z(N171) );
  GTECH_OR2 C445 ( .A(a4stg_rnd_mode[0]), .B(N171), .Z(N172) );
  GTECH_NOT I_47 ( .A(N172), .Z(N173) );
  GTECH_AND2 C447 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N174) );
  GTECH_OR2 C450 ( .A(N73), .B(a1stg_op[7]), .Z(N175) );
  GTECH_OR2 C451 ( .A(a1stg_op[5]), .B(N175), .Z(N176) );
  GTECH_OR2 C452 ( .A(a1stg_op[4]), .B(N176), .Z(N177) );
  GTECH_OR2 C453 ( .A(a1stg_op[3]), .B(N177), .Z(N178) );
  GTECH_OR2 C454 ( .A(a1stg_op[2]), .B(N178), .Z(N179) );
  GTECH_OR2 C455 ( .A(N92), .B(N179), .Z(N180) );
  GTECH_OR2 C456 ( .A(a1stg_op[0]), .B(N180), .Z(N181) );
  GTECH_NOT I_48 ( .A(N181), .Z(N182) );
  GTECH_OR2 C461 ( .A(N73), .B(a1stg_op[7]), .Z(N183) );
  GTECH_OR2 C462 ( .A(a1stg_op[5]), .B(N183), .Z(N184) );
  GTECH_OR2 C463 ( .A(a1stg_op[4]), .B(N184), .Z(N185) );
  GTECH_OR2 C464 ( .A(a1stg_op[3]), .B(N185), .Z(N186) );
  GTECH_OR2 C465 ( .A(N109), .B(N186), .Z(N187) );
  GTECH_OR2 C466 ( .A(N92), .B(N187), .Z(N188) );
  GTECH_OR2 C467 ( .A(a1stg_op[0]), .B(N188), .Z(N189) );
  GTECH_NOT I_49 ( .A(N189), .Z(N190) );
  GTECH_OR2 C472 ( .A(N73), .B(N72), .Z(N191) );
  GTECH_OR2 C473 ( .A(a1stg_op[5]), .B(N191), .Z(N192) );
  GTECH_OR2 C474 ( .A(a1stg_op[4]), .B(N192), .Z(N193) );
  GTECH_OR2 C475 ( .A(N118), .B(N193), .Z(N194) );
  GTECH_OR2 C476 ( .A(a1stg_op[2]), .B(N194), .Z(N195) );
  GTECH_OR2 C477 ( .A(a1stg_op[1]), .B(N195), .Z(N196) );
  GTECH_OR2 C478 ( .A(a1stg_op[0]), .B(N196), .Z(N197) );
  GTECH_NOT I_50 ( .A(N197), .Z(N198) );
  GTECH_OR2 C482 ( .A(a1stg_op[6]), .B(N72), .Z(N199) );
  GTECH_OR2 C483 ( .A(a1stg_op[5]), .B(N199), .Z(N200) );
  GTECH_OR2 C484 ( .A(a1stg_op[4]), .B(N200), .Z(N201) );
  GTECH_OR2 C485 ( .A(N118), .B(N201), .Z(N202) );
  GTECH_OR2 C486 ( .A(a1stg_op[2]), .B(N202), .Z(N203) );
  GTECH_OR2 C487 ( .A(a1stg_op[1]), .B(N203), .Z(N204) );
  GTECH_OR2 C488 ( .A(a1stg_op[0]), .B(N204), .Z(N205) );
  GTECH_NOT I_51 ( .A(N205), .Z(N206) );
  GTECH_OR2 C494 ( .A(N73), .B(N72), .Z(N207) );
  GTECH_OR2 C495 ( .A(a1stg_op[5]), .B(N207), .Z(N208) );
  GTECH_OR2 C496 ( .A(a1stg_op[4]), .B(N208), .Z(N209) );
  GTECH_OR2 C497 ( .A(N118), .B(N209), .Z(N210) );
  GTECH_OR2 C498 ( .A(a1stg_op[2]), .B(N210), .Z(N211) );
  GTECH_OR2 C499 ( .A(a1stg_op[1]), .B(N211), .Z(N212) );
  GTECH_OR2 C500 ( .A(N75), .B(N212), .Z(N213) );
  GTECH_NOT I_52 ( .A(N213), .Z(N214) );
  GTECH_OR2 C504 ( .A(N73), .B(a1stg_op[7]), .Z(N215) );
  GTECH_OR2 C505 ( .A(a1stg_op[5]), .B(N215), .Z(N216) );
  GTECH_OR2 C506 ( .A(a1stg_op[4]), .B(N216), .Z(N217) );
  GTECH_OR2 C507 ( .A(a1stg_op[3]), .B(N217), .Z(N218) );
  GTECH_OR2 C508 ( .A(a1stg_op[2]), .B(N218), .Z(N219) );
  GTECH_OR2 C509 ( .A(a1stg_op[1]), .B(N219), .Z(N220) );
  GTECH_OR2 C510 ( .A(N75), .B(N220), .Z(N221) );
  GTECH_NOT I_53 ( .A(N221), .Z(N222) );
  GTECH_OR2 C515 ( .A(N73), .B(a1stg_op[7]), .Z(N223) );
  GTECH_OR2 C516 ( .A(a1stg_op[5]), .B(N223), .Z(N224) );
  GTECH_OR2 C517 ( .A(a1stg_op[4]), .B(N224), .Z(N225) );
  GTECH_OR2 C518 ( .A(a1stg_op[3]), .B(N225), .Z(N226) );
  GTECH_OR2 C519 ( .A(N109), .B(N226), .Z(N227) );
  GTECH_OR2 C520 ( .A(a1stg_op[1]), .B(N227), .Z(N228) );
  GTECH_OR2 C521 ( .A(N75), .B(N228), .Z(N229) );
  GTECH_NOT I_54 ( .A(N229), .Z(N230) );
  GTECH_OR2 C526 ( .A(N73), .B(N72), .Z(N231) );
  GTECH_OR2 C527 ( .A(a1stg_op[5]), .B(N231), .Z(N232) );
  GTECH_OR2 C528 ( .A(a1stg_op[4]), .B(N232), .Z(N233) );
  GTECH_OR2 C529 ( .A(a1stg_op[3]), .B(N233), .Z(N234) );
  GTECH_OR2 C530 ( .A(N109), .B(N234), .Z(N235) );
  GTECH_OR2 C531 ( .A(a1stg_op[1]), .B(N235), .Z(N236) );
  GTECH_OR2 C532 ( .A(a1stg_op[0]), .B(N236), .Z(N237) );
  GTECH_NOT I_55 ( .A(N237), .Z(N238) );
  GTECH_OR2 C536 ( .A(a1stg_op[6]), .B(N72), .Z(N239) );
  GTECH_OR2 C537 ( .A(a1stg_op[5]), .B(N239), .Z(N240) );
  GTECH_OR2 C538 ( .A(a1stg_op[4]), .B(N240), .Z(N241) );
  GTECH_OR2 C539 ( .A(a1stg_op[3]), .B(N241), .Z(N242) );
  GTECH_OR2 C540 ( .A(N109), .B(N242), .Z(N243) );
  GTECH_OR2 C541 ( .A(a1stg_op[1]), .B(N243), .Z(N244) );
  GTECH_OR2 C542 ( .A(a1stg_op[0]), .B(N244), .Z(N245) );
  GTECH_NOT I_56 ( .A(N245), .Z(N246) );
  GTECH_OR2 C548 ( .A(N73), .B(N72), .Z(N247) );
  GTECH_OR2 C549 ( .A(a1stg_op[5]), .B(N247), .Z(N248) );
  GTECH_OR2 C550 ( .A(a1stg_op[4]), .B(N248), .Z(N249) );
  GTECH_OR2 C551 ( .A(a1stg_op[3]), .B(N249), .Z(N250) );
  GTECH_OR2 C552 ( .A(N109), .B(N250), .Z(N251) );
  GTECH_OR2 C553 ( .A(N92), .B(N251), .Z(N252) );
  GTECH_OR2 C554 ( .A(a1stg_op[0]), .B(N252), .Z(N253) );
  GTECH_NOT I_57 ( .A(N253), .Z(N254) );
  GTECH_OR2 C558 ( .A(a1stg_op[6]), .B(N72), .Z(N255) );
  GTECH_OR2 C559 ( .A(a1stg_op[5]), .B(N255), .Z(N256) );
  GTECH_OR2 C560 ( .A(a1stg_op[4]), .B(N256), .Z(N257) );
  GTECH_OR2 C561 ( .A(a1stg_op[3]), .B(N257), .Z(N258) );
  GTECH_OR2 C562 ( .A(a1stg_op[2]), .B(N258), .Z(N259) );
  GTECH_OR2 C563 ( .A(a1stg_op[1]), .B(N259), .Z(N260) );
  GTECH_OR2 C564 ( .A(N75), .B(N260), .Z(N261) );
  GTECH_NOT I_58 ( .A(N261), .Z(N262) );
  GTECH_OR2 C568 ( .A(a1stg_op[6]), .B(N72), .Z(N263) );
  GTECH_OR2 C569 ( .A(a1stg_op[5]), .B(N263), .Z(N264) );
  GTECH_OR2 C570 ( .A(a1stg_op[4]), .B(N264), .Z(N265) );
  GTECH_OR2 C571 ( .A(a1stg_op[3]), .B(N265), .Z(N266) );
  GTECH_OR2 C572 ( .A(a1stg_op[2]), .B(N266), .Z(N267) );
  GTECH_OR2 C573 ( .A(N92), .B(N267), .Z(N268) );
  GTECH_OR2 C574 ( .A(a1stg_op[0]), .B(N268), .Z(N269) );
  GTECH_NOT I_59 ( .A(N269), .Z(N270) );
  GTECH_OR2 C580 ( .A(N73), .B(N72), .Z(N271) );
  GTECH_OR2 C581 ( .A(a1stg_op[5]), .B(N271), .Z(N272) );
  GTECH_OR2 C582 ( .A(N74), .B(N272), .Z(N273) );
  GTECH_OR2 C583 ( .A(a1stg_op[3]), .B(N273), .Z(N274) );
  GTECH_OR2 C584 ( .A(a1stg_op[2]), .B(N274), .Z(N275) );
  GTECH_OR2 C585 ( .A(a1stg_op[1]), .B(N275), .Z(N276) );
  GTECH_OR2 C586 ( .A(N75), .B(N276), .Z(N277) );
  GTECH_NOT I_60 ( .A(N277), .Z(N278) );
  GTECH_OR2 C592 ( .A(N73), .B(N72), .Z(N279) );
  GTECH_OR2 C593 ( .A(a1stg_op[5]), .B(N279), .Z(N280) );
  GTECH_OR2 C594 ( .A(N74), .B(N280), .Z(N281) );
  GTECH_OR2 C595 ( .A(a1stg_op[3]), .B(N281), .Z(N282) );
  GTECH_OR2 C596 ( .A(a1stg_op[2]), .B(N282), .Z(N283) );
  GTECH_OR2 C597 ( .A(N92), .B(N283), .Z(N284) );
  GTECH_OR2 C598 ( .A(a1stg_op[0]), .B(N284), .Z(N285) );
  GTECH_NOT I_61 ( .A(N285), .Z(N286) );
  GTECH_OR2 C604 ( .A(N73), .B(N72), .Z(N287) );
  GTECH_OR2 C605 ( .A(a1stg_op[5]), .B(N287), .Z(N288) );
  GTECH_OR2 C606 ( .A(N74), .B(N288), .Z(N289) );
  GTECH_OR2 C607 ( .A(a1stg_op[3]), .B(N289), .Z(N290) );
  GTECH_OR2 C608 ( .A(a1stg_op[2]), .B(N290), .Z(N291) );
  GTECH_OR2 C609 ( .A(N92), .B(N291), .Z(N292) );
  GTECH_OR2 C610 ( .A(a1stg_op[0]), .B(N292), .Z(N293) );
  GTECH_NOT I_62 ( .A(N293), .Z(N294) );
  GTECH_OR2 C614 ( .A(a1stg_op[6]), .B(N72), .Z(N295) );
  GTECH_OR2 C615 ( .A(a1stg_op[5]), .B(N295), .Z(N296) );
  GTECH_OR2 C616 ( .A(a1stg_op[4]), .B(N296), .Z(N297) );
  GTECH_OR2 C617 ( .A(a1stg_op[3]), .B(N297), .Z(N298) );
  GTECH_OR2 C618 ( .A(a1stg_op[2]), .B(N298), .Z(N299) );
  GTECH_OR2 C619 ( .A(N92), .B(N299), .Z(N300) );
  GTECH_OR2 C620 ( .A(a1stg_op[0]), .B(N300), .Z(N301) );
  GTECH_NOT I_63 ( .A(N301), .Z(N302) );
  GTECH_OR2 C626 ( .A(N73), .B(N72), .Z(N303) );
  GTECH_OR2 C627 ( .A(a1stg_op[5]), .B(N303), .Z(N304) );
  GTECH_OR2 C628 ( .A(N74), .B(N304), .Z(N305) );
  GTECH_OR2 C629 ( .A(a1stg_op[3]), .B(N305), .Z(N306) );
  GTECH_OR2 C630 ( .A(a1stg_op[2]), .B(N306), .Z(N307) );
  GTECH_OR2 C631 ( .A(a1stg_op[1]), .B(N307), .Z(N308) );
  GTECH_OR2 C632 ( .A(N75), .B(N308), .Z(N309) );
  GTECH_NOT I_64 ( .A(N309), .Z(N310) );
  GTECH_OR2 C636 ( .A(a1stg_op[6]), .B(N72), .Z(N311) );
  GTECH_OR2 C637 ( .A(a1stg_op[5]), .B(N311), .Z(N312) );
  GTECH_OR2 C638 ( .A(a1stg_op[4]), .B(N312), .Z(N313) );
  GTECH_OR2 C639 ( .A(a1stg_op[3]), .B(N313), .Z(N314) );
  GTECH_OR2 C640 ( .A(a1stg_op[2]), .B(N314), .Z(N315) );
  GTECH_OR2 C641 ( .A(a1stg_op[1]), .B(N315), .Z(N316) );
  GTECH_OR2 C642 ( .A(N75), .B(N316), .Z(N317) );
  GTECH_NOT I_65 ( .A(N317), .Z(N318) );
  GTECH_OR2 C648 ( .A(N73), .B(N72), .Z(N319) );
  GTECH_OR2 C649 ( .A(a1stg_op[5]), .B(N319), .Z(N320) );
  GTECH_OR2 C650 ( .A(N74), .B(N320), .Z(N321) );
  GTECH_OR2 C651 ( .A(a1stg_op[3]), .B(N321), .Z(N322) );
  GTECH_OR2 C652 ( .A(a1stg_op[2]), .B(N322), .Z(N323) );
  GTECH_OR2 C653 ( .A(a1stg_op[1]), .B(N323), .Z(N324) );
  GTECH_OR2 C654 ( .A(N75), .B(N324), .Z(N325) );
  GTECH_NOT I_66 ( .A(N325), .Z(N326) );
  GTECH_OR2 C658 ( .A(a1stg_op[6]), .B(N72), .Z(N327) );
  GTECH_OR2 C659 ( .A(a1stg_op[5]), .B(N327), .Z(N328) );
  GTECH_OR2 C660 ( .A(a1stg_op[4]), .B(N328), .Z(N329) );
  GTECH_OR2 C661 ( .A(a1stg_op[3]), .B(N329), .Z(N330) );
  GTECH_OR2 C662 ( .A(a1stg_op[2]), .B(N330), .Z(N331) );
  GTECH_OR2 C663 ( .A(a1stg_op[1]), .B(N331), .Z(N332) );
  GTECH_OR2 C664 ( .A(N75), .B(N332), .Z(N333) );
  GTECH_NOT I_67 ( .A(N333), .Z(N334) );
  GTECH_OR2 C670 ( .A(N73), .B(N72), .Z(N335) );
  GTECH_OR2 C671 ( .A(a1stg_op[5]), .B(N335), .Z(N336) );
  GTECH_OR2 C672 ( .A(N74), .B(N336), .Z(N337) );
  GTECH_OR2 C673 ( .A(a1stg_op[3]), .B(N337), .Z(N338) );
  GTECH_OR2 C674 ( .A(a1stg_op[2]), .B(N338), .Z(N339) );
  GTECH_OR2 C675 ( .A(N92), .B(N339), .Z(N340) );
  GTECH_OR2 C676 ( .A(a1stg_op[0]), .B(N340), .Z(N341) );
  GTECH_NOT I_68 ( .A(N341), .Z(N342) );
  GTECH_OR2 C680 ( .A(a1stg_op[6]), .B(N72), .Z(N343) );
  GTECH_OR2 C681 ( .A(a1stg_op[5]), .B(N343), .Z(N344) );
  GTECH_OR2 C682 ( .A(a1stg_op[4]), .B(N344), .Z(N345) );
  GTECH_OR2 C683 ( .A(a1stg_op[3]), .B(N345), .Z(N346) );
  GTECH_OR2 C684 ( .A(a1stg_op[2]), .B(N346), .Z(N347) );
  GTECH_OR2 C685 ( .A(N92), .B(N347), .Z(N348) );
  GTECH_OR2 C686 ( .A(a1stg_op[0]), .B(N348), .Z(N349) );
  GTECH_NOT I_69 ( .A(N349), .Z(N350) );
  GTECH_OR2 C692 ( .A(N73), .B(N72), .Z(N351) );
  GTECH_OR2 C693 ( .A(a1stg_op[5]), .B(N351), .Z(N352) );
  GTECH_OR2 C694 ( .A(a1stg_op[4]), .B(N352), .Z(N353) );
  GTECH_OR2 C695 ( .A(a1stg_op[3]), .B(N353), .Z(N354) );
  GTECH_OR2 C696 ( .A(N109), .B(N354), .Z(N355) );
  GTECH_OR2 C697 ( .A(N92), .B(N355), .Z(N356) );
  GTECH_OR2 C698 ( .A(a1stg_op[0]), .B(N356), .Z(N357) );
  GTECH_NOT I_70 ( .A(N357), .Z(N358) );
  GTECH_OR2 C703 ( .A(N73), .B(a1stg_op[7]), .Z(N359) );
  GTECH_OR2 C704 ( .A(a1stg_op[5]), .B(N359), .Z(N360) );
  GTECH_OR2 C705 ( .A(N74), .B(N360), .Z(N361) );
  GTECH_OR2 C706 ( .A(a1stg_op[3]), .B(N361), .Z(N362) );
  GTECH_OR2 C707 ( .A(a1stg_op[2]), .B(N362), .Z(N363) );
  GTECH_OR2 C708 ( .A(a1stg_op[1]), .B(N363), .Z(N364) );
  GTECH_OR2 C709 ( .A(N75), .B(N364), .Z(N365) );
  GTECH_NOT I_71 ( .A(N365), .Z(N366) );
  GTECH_OR2 C714 ( .A(N73), .B(a1stg_op[7]), .Z(N367) );
  GTECH_OR2 C715 ( .A(a1stg_op[5]), .B(N367), .Z(N368) );
  GTECH_OR2 C716 ( .A(N74), .B(N368), .Z(N369) );
  GTECH_OR2 C717 ( .A(a1stg_op[3]), .B(N369), .Z(N370) );
  GTECH_OR2 C718 ( .A(a1stg_op[2]), .B(N370), .Z(N371) );
  GTECH_OR2 C719 ( .A(N92), .B(N371), .Z(N372) );
  GTECH_OR2 C720 ( .A(a1stg_op[0]), .B(N372), .Z(N373) );
  GTECH_NOT I_72 ( .A(N373), .Z(N374) );
  GTECH_OR2 C726 ( .A(N73), .B(a1stg_op[7]), .Z(N375) );
  GTECH_OR2 C727 ( .A(a1stg_op[5]), .B(N375), .Z(N376) );
  GTECH_OR2 C728 ( .A(N74), .B(N376), .Z(N377) );
  GTECH_OR2 C729 ( .A(a1stg_op[3]), .B(N377), .Z(N378) );
  GTECH_OR2 C730 ( .A(N109), .B(N378), .Z(N379) );
  GTECH_OR2 C731 ( .A(a1stg_op[1]), .B(N379), .Z(N380) );
  GTECH_OR2 C732 ( .A(N75), .B(N380), .Z(N381) );
  GTECH_NOT I_73 ( .A(N381), .Z(N382) );
  GTECH_OR2 C738 ( .A(N73), .B(a1stg_op[7]), .Z(N383) );
  GTECH_OR2 C739 ( .A(a1stg_op[5]), .B(N383), .Z(N384) );
  GTECH_OR2 C740 ( .A(N74), .B(N384), .Z(N385) );
  GTECH_OR2 C741 ( .A(a1stg_op[3]), .B(N385), .Z(N386) );
  GTECH_OR2 C742 ( .A(N109), .B(N386), .Z(N387) );
  GTECH_OR2 C743 ( .A(N92), .B(N387), .Z(N388) );
  GTECH_OR2 C744 ( .A(a1stg_op[0]), .B(N388), .Z(N389) );
  GTECH_NOT I_74 ( .A(N389), .Z(N390) );
  GTECH_OR2 C748 ( .A(N73), .B(a1stg_op[7]), .Z(N391) );
  GTECH_OR2 C749 ( .A(a1stg_op[5]), .B(N391), .Z(N392) );
  GTECH_OR2 C750 ( .A(a1stg_op[4]), .B(N392), .Z(N393) );
  GTECH_OR2 C751 ( .A(a1stg_op[3]), .B(N393), .Z(N394) );
  GTECH_OR2 C752 ( .A(a1stg_op[2]), .B(N394), .Z(N395) );
  GTECH_OR2 C753 ( .A(a1stg_op[1]), .B(N395), .Z(N396) );
  GTECH_OR2 C754 ( .A(N75), .B(N396), .Z(N397) );
  GTECH_NOT I_75 ( .A(N397), .Z(N398) );
  GTECH_OR2 C758 ( .A(N73), .B(a1stg_op[7]), .Z(N399) );
  GTECH_OR2 C759 ( .A(a1stg_op[5]), .B(N399), .Z(N400) );
  GTECH_OR2 C760 ( .A(a1stg_op[4]), .B(N400), .Z(N401) );
  GTECH_OR2 C761 ( .A(a1stg_op[3]), .B(N401), .Z(N402) );
  GTECH_OR2 C762 ( .A(a1stg_op[2]), .B(N402), .Z(N403) );
  GTECH_OR2 C763 ( .A(N92), .B(N403), .Z(N404) );
  GTECH_OR2 C764 ( .A(a1stg_op[0]), .B(N404), .Z(N405) );
  GTECH_NOT I_76 ( .A(N405), .Z(N406) );
  GTECH_OR2 C769 ( .A(N73), .B(a1stg_op[7]), .Z(N407) );
  GTECH_OR2 C770 ( .A(a1stg_op[5]), .B(N407), .Z(N408) );
  GTECH_OR2 C771 ( .A(a1stg_op[4]), .B(N408), .Z(N409) );
  GTECH_OR2 C772 ( .A(a1stg_op[3]), .B(N409), .Z(N410) );
  GTECH_OR2 C773 ( .A(N109), .B(N410), .Z(N411) );
  GTECH_OR2 C774 ( .A(a1stg_op[1]), .B(N411), .Z(N412) );
  GTECH_OR2 C775 ( .A(N75), .B(N412), .Z(N413) );
  GTECH_NOT I_77 ( .A(N413), .Z(N414) );
  GTECH_OR2 C780 ( .A(N73), .B(a1stg_op[7]), .Z(N415) );
  GTECH_OR2 C781 ( .A(a1stg_op[5]), .B(N415), .Z(N416) );
  GTECH_OR2 C782 ( .A(a1stg_op[4]), .B(N416), .Z(N417) );
  GTECH_OR2 C783 ( .A(a1stg_op[3]), .B(N417), .Z(N418) );
  GTECH_OR2 C784 ( .A(N109), .B(N418), .Z(N419) );
  GTECH_OR2 C785 ( .A(N92), .B(N419), .Z(N420) );
  GTECH_OR2 C786 ( .A(a1stg_op[0]), .B(N420), .Z(N421) );
  GTECH_NOT I_78 ( .A(N421), .Z(N422) );
  GTECH_OR2 C792 ( .A(N73), .B(N72), .Z(N423) );
  GTECH_OR2 C793 ( .A(a1stg_op[5]), .B(N423), .Z(N424) );
  GTECH_OR2 C794 ( .A(a1stg_op[4]), .B(N424), .Z(N425) );
  GTECH_OR2 C795 ( .A(a1stg_op[3]), .B(N425), .Z(N426) );
  GTECH_OR2 C796 ( .A(N109), .B(N426), .Z(N427) );
  GTECH_OR2 C797 ( .A(N92), .B(N427), .Z(N428) );
  GTECH_OR2 C798 ( .A(a1stg_op[0]), .B(N428), .Z(N429) );
  GTECH_NOT I_79 ( .A(N429), .Z(N430) );
  GTECH_OR2 C804 ( .A(N73), .B(N72), .Z(N431) );
  GTECH_OR2 C805 ( .A(a1stg_op[5]), .B(N431), .Z(N432) );
  GTECH_OR2 C806 ( .A(a1stg_op[4]), .B(N432), .Z(N433) );
  GTECH_OR2 C807 ( .A(N118), .B(N433), .Z(N434) );
  GTECH_OR2 C808 ( .A(a1stg_op[2]), .B(N434), .Z(N435) );
  GTECH_OR2 C809 ( .A(a1stg_op[1]), .B(N435), .Z(N436) );
  GTECH_OR2 C810 ( .A(N75), .B(N436), .Z(N437) );
  GTECH_NOT I_80 ( .A(N437), .Z(N438) );
  GTECH_OR2 C815 ( .A(N73), .B(N72), .Z(N439) );
  GTECH_OR2 C816 ( .A(a1stg_op[5]), .B(N439), .Z(N440) );
  GTECH_OR2 C817 ( .A(a1stg_op[4]), .B(N440), .Z(N441) );
  GTECH_OR2 C818 ( .A(N118), .B(N441), .Z(N442) );
  GTECH_OR2 C819 ( .A(a1stg_op[2]), .B(N442), .Z(N443) );
  GTECH_OR2 C820 ( .A(a1stg_op[1]), .B(N443), .Z(N444) );
  GTECH_OR2 C821 ( .A(a1stg_op[0]), .B(N444), .Z(N445) );
  GTECH_NOT I_81 ( .A(N445), .Z(N446) );
  GTECH_OR2 C826 ( .A(N73), .B(N72), .Z(N447) );
  GTECH_OR2 C827 ( .A(a1stg_op[5]), .B(N447), .Z(N448) );
  GTECH_OR2 C828 ( .A(a1stg_op[4]), .B(N448), .Z(N449) );
  GTECH_OR2 C829 ( .A(a1stg_op[3]), .B(N449), .Z(N450) );
  GTECH_OR2 C830 ( .A(N109), .B(N450), .Z(N451) );
  GTECH_OR2 C831 ( .A(a1stg_op[1]), .B(N451), .Z(N452) );
  GTECH_OR2 C832 ( .A(a1stg_op[0]), .B(N452), .Z(N453) );
  GTECH_NOT I_82 ( .A(N453), .Z(N454) );
  GTECH_OR2 C836 ( .A(a1stg_op[6]), .B(N72), .Z(N455) );
  GTECH_OR2 C837 ( .A(a1stg_op[5]), .B(N455), .Z(N456) );
  GTECH_OR2 C838 ( .A(a1stg_op[4]), .B(N456), .Z(N457) );
  GTECH_OR2 C839 ( .A(a1stg_op[3]), .B(N457), .Z(N458) );
  GTECH_OR2 C840 ( .A(N109), .B(N458), .Z(N459) );
  GTECH_OR2 C841 ( .A(a1stg_op[1]), .B(N459), .Z(N460) );
  GTECH_OR2 C842 ( .A(a1stg_op[0]), .B(N460), .Z(N461) );
  GTECH_NOT I_83 ( .A(N461), .Z(N462) );
  GTECH_OR2 C846 ( .A(a1stg_op[6]), .B(N72), .Z(N463) );
  GTECH_OR2 C847 ( .A(a1stg_op[5]), .B(N463), .Z(N464) );
  GTECH_OR2 C848 ( .A(a1stg_op[4]), .B(N464), .Z(N465) );
  GTECH_OR2 C849 ( .A(N118), .B(N465), .Z(N466) );
  GTECH_OR2 C850 ( .A(a1stg_op[2]), .B(N466), .Z(N467) );
  GTECH_OR2 C851 ( .A(a1stg_op[1]), .B(N467), .Z(N468) );
  GTECH_OR2 C852 ( .A(a1stg_op[0]), .B(N468), .Z(N469) );
  GTECH_NOT I_84 ( .A(N469), .Z(N470) );
  GTECH_OR2 C856 ( .A(N73), .B(a1stg_op[7]), .Z(N471) );
  GTECH_OR2 C857 ( .A(a1stg_op[5]), .B(N471), .Z(N472) );
  GTECH_OR2 C858 ( .A(a1stg_op[4]), .B(N472), .Z(N473) );
  GTECH_OR2 C859 ( .A(a1stg_op[3]), .B(N473), .Z(N474) );
  GTECH_OR2 C860 ( .A(a1stg_op[2]), .B(N474), .Z(N475) );
  GTECH_OR2 C861 ( .A(a1stg_op[1]), .B(N475), .Z(N476) );
  GTECH_OR2 C862 ( .A(N75), .B(N476), .Z(N477) );
  GTECH_NOT I_85 ( .A(N477), .Z(N478) );
  GTECH_OR2 C867 ( .A(N73), .B(a1stg_op[7]), .Z(N479) );
  GTECH_OR2 C868 ( .A(a1stg_op[5]), .B(N479), .Z(N480) );
  GTECH_OR2 C869 ( .A(a1stg_op[4]), .B(N480), .Z(N481) );
  GTECH_OR2 C870 ( .A(a1stg_op[3]), .B(N481), .Z(N482) );
  GTECH_OR2 C871 ( .A(N109), .B(N482), .Z(N483) );
  GTECH_OR2 C872 ( .A(a1stg_op[1]), .B(N483), .Z(N484) );
  GTECH_OR2 C873 ( .A(N75), .B(N484), .Z(N485) );
  GTECH_NOT I_86 ( .A(N485), .Z(N486) );
  GTECH_OR2 C879 ( .A(N73), .B(N72), .Z(N487) );
  GTECH_OR2 C880 ( .A(a1stg_op[5]), .B(N487), .Z(N488) );
  GTECH_OR2 C881 ( .A(a1stg_op[4]), .B(N488), .Z(N489) );
  GTECH_OR2 C882 ( .A(a1stg_op[3]), .B(N489), .Z(N490) );
  GTECH_OR2 C883 ( .A(N109), .B(N490), .Z(N491) );
  GTECH_OR2 C884 ( .A(N92), .B(N491), .Z(N492) );
  GTECH_OR2 C885 ( .A(a1stg_op[0]), .B(N492), .Z(N493) );
  GTECH_NOT I_87 ( .A(N493), .Z(N494) );
  GTECH_OR2 C889 ( .A(N73), .B(a1stg_op[7]), .Z(N495) );
  GTECH_OR2 C890 ( .A(a1stg_op[5]), .B(N495), .Z(N496) );
  GTECH_OR2 C891 ( .A(a1stg_op[4]), .B(N496), .Z(N497) );
  GTECH_OR2 C892 ( .A(a1stg_op[3]), .B(N497), .Z(N498) );
  GTECH_OR2 C893 ( .A(a1stg_op[2]), .B(N498), .Z(N499) );
  GTECH_OR2 C894 ( .A(a1stg_op[1]), .B(N499), .Z(N500) );
  GTECH_OR2 C895 ( .A(N75), .B(N500), .Z(N501) );
  GTECH_NOT I_88 ( .A(N501), .Z(N502) );
  GTECH_OR2 C900 ( .A(N73), .B(a1stg_op[7]), .Z(N503) );
  GTECH_OR2 C901 ( .A(a1stg_op[5]), .B(N503), .Z(N504) );
  GTECH_OR2 C902 ( .A(a1stg_op[4]), .B(N504), .Z(N505) );
  GTECH_OR2 C903 ( .A(a1stg_op[3]), .B(N505), .Z(N506) );
  GTECH_OR2 C904 ( .A(N109), .B(N506), .Z(N507) );
  GTECH_OR2 C905 ( .A(a1stg_op[1]), .B(N507), .Z(N508) );
  GTECH_OR2 C906 ( .A(N75), .B(N508), .Z(N509) );
  GTECH_NOT I_89 ( .A(N509), .Z(N510) );
  GTECH_OR2 C910 ( .A(N73), .B(a1stg_op[7]), .Z(N511) );
  GTECH_OR2 C911 ( .A(a1stg_op[5]), .B(N511), .Z(N512) );
  GTECH_OR2 C912 ( .A(a1stg_op[4]), .B(N512), .Z(N513) );
  GTECH_OR2 C913 ( .A(a1stg_op[3]), .B(N513), .Z(N514) );
  GTECH_OR2 C914 ( .A(a1stg_op[2]), .B(N514), .Z(N515) );
  GTECH_OR2 C915 ( .A(N92), .B(N515), .Z(N516) );
  GTECH_OR2 C916 ( .A(a1stg_op[0]), .B(N516), .Z(N517) );
  GTECH_NOT I_90 ( .A(N517), .Z(N518) );
  GTECH_OR2 C921 ( .A(N73), .B(a1stg_op[7]), .Z(N519) );
  GTECH_OR2 C922 ( .A(a1stg_op[5]), .B(N519), .Z(N520) );
  GTECH_OR2 C923 ( .A(a1stg_op[4]), .B(N520), .Z(N521) );
  GTECH_OR2 C924 ( .A(a1stg_op[3]), .B(N521), .Z(N522) );
  GTECH_OR2 C925 ( .A(N109), .B(N522), .Z(N523) );
  GTECH_OR2 C926 ( .A(N92), .B(N523), .Z(N524) );
  GTECH_OR2 C927 ( .A(a1stg_op[0]), .B(N524), .Z(N525) );
  GTECH_NOT I_91 ( .A(N525), .Z(N526) );
  GTECH_OR2 C932 ( .A(N73), .B(N72), .Z(N527) );
  GTECH_OR2 C933 ( .A(a1stg_op[5]), .B(N527), .Z(N528) );
  GTECH_OR2 C934 ( .A(a1stg_op[4]), .B(N528), .Z(N529) );
  GTECH_OR2 C935 ( .A(N118), .B(N529), .Z(N530) );
  GTECH_OR2 C936 ( .A(a1stg_op[2]), .B(N530), .Z(N531) );
  GTECH_OR2 C937 ( .A(a1stg_op[1]), .B(N531), .Z(N532) );
  GTECH_OR2 C938 ( .A(a1stg_op[0]), .B(N532), .Z(N533) );
  GTECH_NOT I_92 ( .A(N533), .Z(N534) );
  GTECH_OR2 C944 ( .A(N73), .B(N72), .Z(N535) );
  GTECH_OR2 C945 ( .A(a1stg_op[5]), .B(N535), .Z(N536) );
  GTECH_OR2 C946 ( .A(a1stg_op[4]), .B(N536), .Z(N537) );
  GTECH_OR2 C947 ( .A(N118), .B(N537), .Z(N538) );
  GTECH_OR2 C948 ( .A(a1stg_op[2]), .B(N538), .Z(N539) );
  GTECH_OR2 C949 ( .A(a1stg_op[1]), .B(N539), .Z(N540) );
  GTECH_OR2 C950 ( .A(N75), .B(N540), .Z(N541) );
  GTECH_NOT I_93 ( .A(N541), .Z(N542) );
  GTECH_OR2 C955 ( .A(N73), .B(N72), .Z(N543) );
  GTECH_OR2 C956 ( .A(a1stg_op[5]), .B(N543), .Z(N544) );
  GTECH_OR2 C957 ( .A(a1stg_op[4]), .B(N544), .Z(N545) );
  GTECH_OR2 C958 ( .A(a1stg_op[3]), .B(N545), .Z(N546) );
  GTECH_OR2 C959 ( .A(N109), .B(N546), .Z(N547) );
  GTECH_OR2 C960 ( .A(a1stg_op[1]), .B(N547), .Z(N548) );
  GTECH_OR2 C961 ( .A(a1stg_op[0]), .B(N548), .Z(N549) );
  GTECH_NOT I_94 ( .A(N549), .Z(N550) );
  GTECH_OR2 C965 ( .A(a1stg_op[6]), .B(N72), .Z(N551) );
  GTECH_OR2 C966 ( .A(a1stg_op[5]), .B(N551), .Z(N552) );
  GTECH_OR2 C967 ( .A(a1stg_op[4]), .B(N552), .Z(N553) );
  GTECH_OR2 C968 ( .A(a1stg_op[3]), .B(N553), .Z(N554) );
  GTECH_OR2 C969 ( .A(N109), .B(N554), .Z(N555) );
  GTECH_OR2 C970 ( .A(a1stg_op[1]), .B(N555), .Z(N556) );
  GTECH_OR2 C971 ( .A(a1stg_op[0]), .B(N556), .Z(N557) );
  GTECH_NOT I_95 ( .A(N557), .Z(N558) );
  GTECH_OR2 C975 ( .A(N73), .B(a1stg_op[7]), .Z(N559) );
  GTECH_OR2 C976 ( .A(a1stg_op[5]), .B(N559), .Z(N560) );
  GTECH_OR2 C977 ( .A(a1stg_op[4]), .B(N560), .Z(N561) );
  GTECH_OR2 C978 ( .A(a1stg_op[3]), .B(N561), .Z(N562) );
  GTECH_OR2 C979 ( .A(a1stg_op[2]), .B(N562), .Z(N563) );
  GTECH_OR2 C980 ( .A(a1stg_op[1]), .B(N563), .Z(N564) );
  GTECH_OR2 C981 ( .A(N75), .B(N564), .Z(N565) );
  GTECH_NOT I_96 ( .A(N565), .Z(N566) );
  GTECH_OR2 C985 ( .A(N73), .B(a1stg_op[7]), .Z(N567) );
  GTECH_OR2 C986 ( .A(a1stg_op[5]), .B(N567), .Z(N568) );
  GTECH_OR2 C987 ( .A(a1stg_op[4]), .B(N568), .Z(N569) );
  GTECH_OR2 C988 ( .A(a1stg_op[3]), .B(N569), .Z(N570) );
  GTECH_OR2 C989 ( .A(a1stg_op[2]), .B(N570), .Z(N571) );
  GTECH_OR2 C990 ( .A(N92), .B(N571), .Z(N572) );
  GTECH_OR2 C991 ( .A(a1stg_op[0]), .B(N572), .Z(N573) );
  GTECH_NOT I_97 ( .A(N573), .Z(N574) );
  GTECH_OR2 C996 ( .A(N73), .B(a1stg_op[7]), .Z(N575) );
  GTECH_OR2 C997 ( .A(a1stg_op[5]), .B(N575), .Z(N576) );
  GTECH_OR2 C998 ( .A(a1stg_op[4]), .B(N576), .Z(N577) );
  GTECH_OR2 C999 ( .A(a1stg_op[3]), .B(N577), .Z(N578) );
  GTECH_OR2 C1000 ( .A(N109), .B(N578), .Z(N579) );
  GTECH_OR2 C1001 ( .A(a1stg_op[1]), .B(N579), .Z(N580) );
  GTECH_OR2 C1002 ( .A(N75), .B(N580), .Z(N581) );
  GTECH_NOT I_98 ( .A(N581), .Z(N582) );
  GTECH_OR2 C1007 ( .A(N73), .B(a1stg_op[7]), .Z(N583) );
  GTECH_OR2 C1008 ( .A(a1stg_op[5]), .B(N583), .Z(N584) );
  GTECH_OR2 C1009 ( .A(a1stg_op[4]), .B(N584), .Z(N585) );
  GTECH_OR2 C1010 ( .A(a1stg_op[3]), .B(N585), .Z(N586) );
  GTECH_OR2 C1011 ( .A(N109), .B(N586), .Z(N587) );
  GTECH_OR2 C1012 ( .A(N92), .B(N587), .Z(N588) );
  GTECH_OR2 C1013 ( .A(a1stg_op[0]), .B(N588), .Z(N589) );
  GTECH_NOT I_99 ( .A(N589), .Z(N590) );
  GTECH_OR2 C1019 ( .A(N73), .B(a1stg_op[7]), .Z(N591) );
  GTECH_OR2 C1020 ( .A(a1stg_op[5]), .B(N591), .Z(N592) );
  GTECH_OR2 C1021 ( .A(N74), .B(N592), .Z(N593) );
  GTECH_OR2 C1022 ( .A(a1stg_op[3]), .B(N593), .Z(N594) );
  GTECH_OR2 C1023 ( .A(N109), .B(N594), .Z(N595) );
  GTECH_OR2 C1024 ( .A(a1stg_op[1]), .B(N595), .Z(N596) );
  GTECH_OR2 C1025 ( .A(N75), .B(N596), .Z(N597) );
  GTECH_NOT I_100 ( .A(N597), .Z(N598) );
  GTECH_OR2 C1031 ( .A(N73), .B(a1stg_op[7]), .Z(N599) );
  GTECH_OR2 C1032 ( .A(a1stg_op[5]), .B(N599), .Z(N600) );
  GTECH_OR2 C1033 ( .A(N74), .B(N600), .Z(N601) );
  GTECH_OR2 C1034 ( .A(a1stg_op[3]), .B(N601), .Z(N602) );
  GTECH_OR2 C1035 ( .A(N109), .B(N602), .Z(N603) );
  GTECH_OR2 C1036 ( .A(N92), .B(N603), .Z(N604) );
  GTECH_OR2 C1037 ( .A(a1stg_op[0]), .B(N604), .Z(N605) );
  GTECH_NOT I_101 ( .A(N605), .Z(N606) );
  GTECH_OR2 C1042 ( .A(N73), .B(a1stg_op[7]), .Z(N607) );
  GTECH_OR2 C1043 ( .A(a1stg_op[5]), .B(N607), .Z(N608) );
  GTECH_OR2 C1044 ( .A(N74), .B(N608), .Z(N609) );
  GTECH_OR2 C1045 ( .A(a1stg_op[3]), .B(N609), .Z(N610) );
  GTECH_OR2 C1046 ( .A(a1stg_op[2]), .B(N610), .Z(N611) );
  GTECH_OR2 C1047 ( .A(a1stg_op[1]), .B(N611), .Z(N612) );
  GTECH_OR2 C1048 ( .A(N75), .B(N612), .Z(N613) );
  GTECH_NOT I_102 ( .A(N613), .Z(N614) );
  GTECH_OR2 C1053 ( .A(N73), .B(a1stg_op[7]), .Z(N615) );
  GTECH_OR2 C1054 ( .A(a1stg_op[5]), .B(N615), .Z(N616) );
  GTECH_OR2 C1055 ( .A(N74), .B(N616), .Z(N617) );
  GTECH_OR2 C1056 ( .A(a1stg_op[3]), .B(N617), .Z(N618) );
  GTECH_OR2 C1057 ( .A(a1stg_op[2]), .B(N618), .Z(N619) );
  GTECH_OR2 C1058 ( .A(N92), .B(N619), .Z(N620) );
  GTECH_OR2 C1059 ( .A(a1stg_op[0]), .B(N620), .Z(N621) );
  GTECH_NOT I_103 ( .A(N621), .Z(N622) );
  GTECH_OR2 C1064 ( .A(N73), .B(N72), .Z(N623) );
  GTECH_OR2 C1065 ( .A(a1stg_op[5]), .B(N623), .Z(N624) );
  GTECH_OR2 C1066 ( .A(a1stg_op[4]), .B(N624), .Z(N625) );
  GTECH_OR2 C1067 ( .A(a1stg_op[3]), .B(N625), .Z(N626) );
  GTECH_OR2 C1068 ( .A(N109), .B(N626), .Z(N627) );
  GTECH_OR2 C1069 ( .A(a1stg_op[1]), .B(N627), .Z(N628) );
  GTECH_OR2 C1070 ( .A(a1stg_op[0]), .B(N628), .Z(N629) );
  GTECH_NOT I_104 ( .A(N629), .Z(N630) );
  GTECH_OR2 C1075 ( .A(N73), .B(N72), .Z(N631) );
  GTECH_OR2 C1076 ( .A(a1stg_op[5]), .B(N631), .Z(N632) );
  GTECH_OR2 C1077 ( .A(a1stg_op[4]), .B(N632), .Z(N633) );
  GTECH_OR2 C1078 ( .A(N118), .B(N633), .Z(N634) );
  GTECH_OR2 C1079 ( .A(a1stg_op[2]), .B(N634), .Z(N635) );
  GTECH_OR2 C1080 ( .A(a1stg_op[1]), .B(N635), .Z(N636) );
  GTECH_OR2 C1081 ( .A(a1stg_op[0]), .B(N636), .Z(N637) );
  GTECH_NOT I_105 ( .A(N637), .Z(N638) );
  GTECH_OR2 C1085 ( .A(a1stg_op[6]), .B(N72), .Z(N639) );
  GTECH_OR2 C1086 ( .A(a1stg_op[5]), .B(N639), .Z(N640) );
  GTECH_OR2 C1087 ( .A(a1stg_op[4]), .B(N640), .Z(N641) );
  GTECH_OR2 C1088 ( .A(a1stg_op[3]), .B(N641), .Z(N642) );
  GTECH_OR2 C1089 ( .A(N109), .B(N642), .Z(N643) );
  GTECH_OR2 C1090 ( .A(a1stg_op[1]), .B(N643), .Z(N644) );
  GTECH_OR2 C1091 ( .A(a1stg_op[0]), .B(N644), .Z(N645) );
  GTECH_NOT I_106 ( .A(N645), .Z(N646) );
  GTECH_OR2 C1095 ( .A(a1stg_op[6]), .B(N72), .Z(N647) );
  GTECH_OR2 C1096 ( .A(a1stg_op[5]), .B(N647), .Z(N648) );
  GTECH_OR2 C1097 ( .A(a1stg_op[4]), .B(N648), .Z(N649) );
  GTECH_OR2 C1098 ( .A(N118), .B(N649), .Z(N650) );
  GTECH_OR2 C1099 ( .A(a1stg_op[2]), .B(N650), .Z(N651) );
  GTECH_OR2 C1100 ( .A(a1stg_op[1]), .B(N651), .Z(N652) );
  GTECH_OR2 C1101 ( .A(a1stg_op[0]), .B(N652), .Z(N653) );
  GTECH_NOT I_107 ( .A(N653), .Z(N654) );
  GTECH_OR2 C1107 ( .A(N73), .B(N72), .Z(N655) );
  GTECH_OR2 C1108 ( .A(a1stg_op[5]), .B(N655), .Z(N656) );
  GTECH_OR2 C1109 ( .A(N74), .B(N656), .Z(N657) );
  GTECH_OR2 C1110 ( .A(a1stg_op[3]), .B(N657), .Z(N658) );
  GTECH_OR2 C1111 ( .A(a1stg_op[2]), .B(N658), .Z(N659) );
  GTECH_OR2 C1112 ( .A(a1stg_op[1]), .B(N659), .Z(N660) );
  GTECH_OR2 C1113 ( .A(N75), .B(N660), .Z(N661) );
  GTECH_NOT I_108 ( .A(N661), .Z(N662) );
  GTECH_OR2 C1117 ( .A(a1stg_op[6]), .B(N72), .Z(N663) );
  GTECH_OR2 C1118 ( .A(a1stg_op[5]), .B(N663), .Z(N664) );
  GTECH_OR2 C1119 ( .A(a1stg_op[4]), .B(N664), .Z(N665) );
  GTECH_OR2 C1120 ( .A(a1stg_op[3]), .B(N665), .Z(N666) );
  GTECH_OR2 C1121 ( .A(a1stg_op[2]), .B(N666), .Z(N667) );
  GTECH_OR2 C1122 ( .A(a1stg_op[1]), .B(N667), .Z(N668) );
  GTECH_OR2 C1123 ( .A(N75), .B(N668), .Z(N669) );
  GTECH_NOT I_109 ( .A(N669), .Z(N670) );
  GTECH_OR2 C1129 ( .A(N73), .B(N72), .Z(N671) );
  GTECH_OR2 C1130 ( .A(a1stg_op[5]), .B(N671), .Z(N672) );
  GTECH_OR2 C1131 ( .A(N74), .B(N672), .Z(N673) );
  GTECH_OR2 C1132 ( .A(a1stg_op[3]), .B(N673), .Z(N674) );
  GTECH_OR2 C1133 ( .A(a1stg_op[2]), .B(N674), .Z(N675) );
  GTECH_OR2 C1134 ( .A(N92), .B(N675), .Z(N676) );
  GTECH_OR2 C1135 ( .A(a1stg_op[0]), .B(N676), .Z(N677) );
  GTECH_NOT I_110 ( .A(N677), .Z(N678) );
  GTECH_OR2 C1139 ( .A(a1stg_op[6]), .B(N72), .Z(N679) );
  GTECH_OR2 C1140 ( .A(a1stg_op[5]), .B(N679), .Z(N680) );
  GTECH_OR2 C1141 ( .A(a1stg_op[4]), .B(N680), .Z(N681) );
  GTECH_OR2 C1142 ( .A(a1stg_op[3]), .B(N681), .Z(N682) );
  GTECH_OR2 C1143 ( .A(a1stg_op[2]), .B(N682), .Z(N683) );
  GTECH_OR2 C1144 ( .A(N92), .B(N683), .Z(N684) );
  GTECH_OR2 C1145 ( .A(a1stg_op[0]), .B(N684), .Z(N685) );
  GTECH_NOT I_111 ( .A(N685), .Z(N686) );
  GTECH_OR2 C1151 ( .A(N73), .B(N72), .Z(N687) );
  GTECH_OR2 C1152 ( .A(a1stg_op[5]), .B(N687), .Z(N688) );
  GTECH_OR2 C1153 ( .A(a1stg_op[4]), .B(N688), .Z(N689) );
  GTECH_OR2 C1154 ( .A(N118), .B(N689), .Z(N690) );
  GTECH_OR2 C1155 ( .A(a1stg_op[2]), .B(N690), .Z(N691) );
  GTECH_OR2 C1156 ( .A(a1stg_op[1]), .B(N691), .Z(N692) );
  GTECH_OR2 C1157 ( .A(N75), .B(N692), .Z(N693) );
  GTECH_NOT I_112 ( .A(N693), .Z(N694) );
  GTECH_OR2 C1163 ( .A(N73), .B(N72), .Z(N695) );
  GTECH_OR2 C1164 ( .A(a1stg_op[5]), .B(N695), .Z(N696) );
  GTECH_OR2 C1165 ( .A(a1stg_op[4]), .B(N696), .Z(N697) );
  GTECH_OR2 C1166 ( .A(a1stg_op[3]), .B(N697), .Z(N698) );
  GTECH_OR2 C1167 ( .A(N109), .B(N698), .Z(N699) );
  GTECH_OR2 C1168 ( .A(N92), .B(N699), .Z(N700) );
  GTECH_OR2 C1169 ( .A(a1stg_op[0]), .B(N700), .Z(N701) );
  GTECH_NOT I_113 ( .A(N701), .Z(N702) );
  GTECH_AND2 C1171 ( .A(a2stg_rnd_mode[0]), .B(a2stg_rnd_mode[1]), .Z(N703) );
  GTECH_OR2 C1176 ( .A(N73), .B(a1stg_op[7]), .Z(N704) );
  GTECH_OR2 C1177 ( .A(a1stg_op[5]), .B(N704), .Z(N705) );
  GTECH_OR2 C1178 ( .A(N74), .B(N705), .Z(N706) );
  GTECH_OR2 C1179 ( .A(a1stg_op[3]), .B(N706), .Z(N707) );
  GTECH_OR2 C1180 ( .A(N109), .B(N707), .Z(N708) );
  GTECH_OR2 C1181 ( .A(a1stg_op[1]), .B(N708), .Z(N709) );
  GTECH_OR2 C1182 ( .A(N75), .B(N709), .Z(N710) );
  GTECH_NOT I_114 ( .A(N710), .Z(N711) );
  GTECH_OR2 C1188 ( .A(N73), .B(a1stg_op[7]), .Z(N712) );
  GTECH_OR2 C1189 ( .A(a1stg_op[5]), .B(N712), .Z(N713) );
  GTECH_OR2 C1190 ( .A(N74), .B(N713), .Z(N714) );
  GTECH_OR2 C1191 ( .A(a1stg_op[3]), .B(N714), .Z(N715) );
  GTECH_OR2 C1192 ( .A(N109), .B(N715), .Z(N716) );
  GTECH_OR2 C1193 ( .A(N92), .B(N716), .Z(N717) );
  GTECH_OR2 C1194 ( .A(a1stg_op[0]), .B(N717), .Z(N718) );
  GTECH_NOT I_115 ( .A(N718), .Z(N719) );
  GTECH_OR2 C1199 ( .A(N73), .B(a1stg_op[7]), .Z(N720) );
  GTECH_OR2 C1200 ( .A(a1stg_op[5]), .B(N720), .Z(N721) );
  GTECH_OR2 C1201 ( .A(N74), .B(N721), .Z(N722) );
  GTECH_OR2 C1202 ( .A(a1stg_op[3]), .B(N722), .Z(N723) );
  GTECH_OR2 C1203 ( .A(a1stg_op[2]), .B(N723), .Z(N724) );
  GTECH_OR2 C1204 ( .A(a1stg_op[1]), .B(N724), .Z(N725) );
  GTECH_OR2 C1205 ( .A(N75), .B(N725), .Z(N726) );
  GTECH_NOT I_116 ( .A(N726), .Z(N727) );
  GTECH_OR2 C1210 ( .A(N73), .B(a1stg_op[7]), .Z(N728) );
  GTECH_OR2 C1211 ( .A(a1stg_op[5]), .B(N728), .Z(N729) );
  GTECH_OR2 C1212 ( .A(N74), .B(N729), .Z(N730) );
  GTECH_OR2 C1213 ( .A(a1stg_op[3]), .B(N730), .Z(N731) );
  GTECH_OR2 C1214 ( .A(a1stg_op[2]), .B(N731), .Z(N732) );
  GTECH_OR2 C1215 ( .A(N92), .B(N732), .Z(N733) );
  GTECH_OR2 C1216 ( .A(a1stg_op[0]), .B(N733), .Z(N734) );
  GTECH_NOT I_117 ( .A(N734), .Z(N735) );
  GTECH_OR2 C1221 ( .A(N73), .B(N72), .Z(N736) );
  GTECH_OR2 C1222 ( .A(a1stg_op[5]), .B(N736), .Z(N737) );
  GTECH_OR2 C1223 ( .A(a1stg_op[4]), .B(N737), .Z(N738) );
  GTECH_OR2 C1224 ( .A(a1stg_op[3]), .B(N738), .Z(N739) );
  GTECH_OR2 C1225 ( .A(N109), .B(N739), .Z(N740) );
  GTECH_OR2 C1226 ( .A(a1stg_op[1]), .B(N740), .Z(N741) );
  GTECH_OR2 C1227 ( .A(a1stg_op[0]), .B(N741), .Z(N742) );
  GTECH_NOT I_118 ( .A(N742), .Z(N743) );
  GTECH_OR2 C1232 ( .A(N73), .B(N72), .Z(N744) );
  GTECH_OR2 C1233 ( .A(a1stg_op[5]), .B(N744), .Z(N745) );
  GTECH_OR2 C1234 ( .A(a1stg_op[4]), .B(N745), .Z(N746) );
  GTECH_OR2 C1235 ( .A(N118), .B(N746), .Z(N747) );
  GTECH_OR2 C1236 ( .A(a1stg_op[2]), .B(N747), .Z(N748) );
  GTECH_OR2 C1237 ( .A(a1stg_op[1]), .B(N748), .Z(N749) );
  GTECH_OR2 C1238 ( .A(a1stg_op[0]), .B(N749), .Z(N750) );
  GTECH_NOT I_119 ( .A(N750), .Z(N751) );
  GTECH_OR2 C1242 ( .A(a1stg_op[6]), .B(N72), .Z(N752) );
  GTECH_OR2 C1243 ( .A(a1stg_op[5]), .B(N752), .Z(N753) );
  GTECH_OR2 C1244 ( .A(a1stg_op[4]), .B(N753), .Z(N754) );
  GTECH_OR2 C1245 ( .A(a1stg_op[3]), .B(N754), .Z(N755) );
  GTECH_OR2 C1246 ( .A(N109), .B(N755), .Z(N756) );
  GTECH_OR2 C1247 ( .A(a1stg_op[1]), .B(N756), .Z(N757) );
  GTECH_OR2 C1248 ( .A(a1stg_op[0]), .B(N757), .Z(N758) );
  GTECH_NOT I_120 ( .A(N758), .Z(N759) );
  GTECH_OR2 C1252 ( .A(a1stg_op[6]), .B(N72), .Z(N760) );
  GTECH_OR2 C1253 ( .A(a1stg_op[5]), .B(N760), .Z(N761) );
  GTECH_OR2 C1254 ( .A(a1stg_op[4]), .B(N761), .Z(N762) );
  GTECH_OR2 C1255 ( .A(N118), .B(N762), .Z(N763) );
  GTECH_OR2 C1256 ( .A(a1stg_op[2]), .B(N763), .Z(N764) );
  GTECH_OR2 C1257 ( .A(a1stg_op[1]), .B(N764), .Z(N765) );
  GTECH_OR2 C1258 ( .A(a1stg_op[0]), .B(N765), .Z(N766) );
  GTECH_NOT I_121 ( .A(N766), .Z(N767) );
  GTECH_OR2 C1264 ( .A(N73), .B(N72), .Z(N768) );
  GTECH_OR2 C1265 ( .A(a1stg_op[5]), .B(N768), .Z(N769) );
  GTECH_OR2 C1266 ( .A(a1stg_op[4]), .B(N769), .Z(N770) );
  GTECH_OR2 C1267 ( .A(a1stg_op[3]), .B(N770), .Z(N771) );
  GTECH_OR2 C1268 ( .A(N109), .B(N771), .Z(N772) );
  GTECH_OR2 C1269 ( .A(N92), .B(N772), .Z(N773) );
  GTECH_OR2 C1270 ( .A(a1stg_op[0]), .B(N773), .Z(N774) );
  GTECH_NOT I_122 ( .A(N774), .Z(N775) );
  GTECH_OR2 C1275 ( .A(N73), .B(a1stg_op[7]), .Z(N776) );
  GTECH_OR2 C1276 ( .A(a1stg_op[5]), .B(N776), .Z(N777) );
  GTECH_OR2 C1277 ( .A(a1stg_op[4]), .B(N777), .Z(N778) );
  GTECH_OR2 C1278 ( .A(a1stg_op[3]), .B(N778), .Z(N779) );
  GTECH_OR2 C1279 ( .A(N109), .B(N779), .Z(N780) );
  GTECH_OR2 C1280 ( .A(a1stg_op[1]), .B(N780), .Z(N781) );
  GTECH_OR2 C1281 ( .A(N75), .B(N781), .Z(N782) );
  GTECH_NOT I_123 ( .A(N782), .Z(N783) );
  GTECH_OR2 C1286 ( .A(N73), .B(a1stg_op[7]), .Z(N784) );
  GTECH_OR2 C1287 ( .A(a1stg_op[5]), .B(N784), .Z(N785) );
  GTECH_OR2 C1288 ( .A(a1stg_op[4]), .B(N785), .Z(N786) );
  GTECH_OR2 C1289 ( .A(a1stg_op[3]), .B(N786), .Z(N787) );
  GTECH_OR2 C1290 ( .A(N109), .B(N787), .Z(N788) );
  GTECH_OR2 C1291 ( .A(N92), .B(N788), .Z(N789) );
  GTECH_OR2 C1292 ( .A(a1stg_op[0]), .B(N789), .Z(N790) );
  GTECH_NOT I_124 ( .A(N790), .Z(N791) );
  GTECH_OR2 C1298 ( .A(N73), .B(N72), .Z(N792) );
  GTECH_OR2 C1299 ( .A(a1stg_op[5]), .B(N792), .Z(N793) );
  GTECH_OR2 C1300 ( .A(N74), .B(N793), .Z(N794) );
  GTECH_OR2 C1301 ( .A(a1stg_op[3]), .B(N794), .Z(N795) );
  GTECH_OR2 C1302 ( .A(a1stg_op[2]), .B(N795), .Z(N796) );
  GTECH_OR2 C1303 ( .A(a1stg_op[1]), .B(N796), .Z(N797) );
  GTECH_OR2 C1304 ( .A(N75), .B(N797), .Z(N798) );
  GTECH_NOT I_125 ( .A(N798), .Z(N799) );
  GTECH_OR2 C1308 ( .A(a1stg_op[6]), .B(N72), .Z(N800) );
  GTECH_OR2 C1309 ( .A(a1stg_op[5]), .B(N800), .Z(N801) );
  GTECH_OR2 C1310 ( .A(a1stg_op[4]), .B(N801), .Z(N802) );
  GTECH_OR2 C1311 ( .A(a1stg_op[3]), .B(N802), .Z(N803) );
  GTECH_OR2 C1312 ( .A(a1stg_op[2]), .B(N803), .Z(N804) );
  GTECH_OR2 C1313 ( .A(a1stg_op[1]), .B(N804), .Z(N805) );
  GTECH_OR2 C1314 ( .A(N75), .B(N805), .Z(N806) );
  GTECH_NOT I_126 ( .A(N806), .Z(N807) );
  GTECH_OR2 C1320 ( .A(N73), .B(N72), .Z(N808) );
  GTECH_OR2 C1321 ( .A(a1stg_op[5]), .B(N808), .Z(N809) );
  GTECH_OR2 C1322 ( .A(N74), .B(N809), .Z(N810) );
  GTECH_OR2 C1323 ( .A(a1stg_op[3]), .B(N810), .Z(N811) );
  GTECH_OR2 C1324 ( .A(a1stg_op[2]), .B(N811), .Z(N812) );
  GTECH_OR2 C1325 ( .A(N92), .B(N812), .Z(N813) );
  GTECH_OR2 C1326 ( .A(a1stg_op[0]), .B(N813), .Z(N814) );
  GTECH_NOT I_127 ( .A(N814), .Z(N815) );
  GTECH_OR2 C1330 ( .A(a1stg_op[6]), .B(N72), .Z(N816) );
  GTECH_OR2 C1331 ( .A(a1stg_op[5]), .B(N816), .Z(N817) );
  GTECH_OR2 C1332 ( .A(a1stg_op[4]), .B(N817), .Z(N818) );
  GTECH_OR2 C1333 ( .A(a1stg_op[3]), .B(N818), .Z(N819) );
  GTECH_OR2 C1334 ( .A(a1stg_op[2]), .B(N819), .Z(N820) );
  GTECH_OR2 C1335 ( .A(N92), .B(N820), .Z(N821) );
  GTECH_OR2 C1336 ( .A(a1stg_op[0]), .B(N821), .Z(N822) );
  GTECH_NOT I_128 ( .A(N822), .Z(N823) );
  GTECH_OR2 C1339 ( .A(a4stg_rnd_mode[0]), .B(N171), .Z(N824) );
  GTECH_NOT I_129 ( .A(N824), .Z(N825) );
  GTECH_AND2 C1341 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N826) );
  GTECH_OR2 C1342 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N827) );
  GTECH_NOT I_130 ( .A(N827), .Z(N828) );
  GTECH_OR2 C1345 ( .A(a4stg_rnd_mode[0]), .B(N171), .Z(N829) );
  GTECH_NOT I_131 ( .A(N829), .Z(N830) );
  GTECH_AND2 C1347 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N831) );
  GTECH_OR2 C1348 ( .A(a4stg_rnd_mode[0]), .B(a4stg_rnd_mode[1]), .Z(N832) );
  GTECH_NOT I_132 ( .A(N832), .Z(N833) );
  GTECH_OR2 C1352 ( .A(a1stg_op[6]), .B(N72), .Z(N834) );
  GTECH_OR2 C1353 ( .A(a1stg_op[5]), .B(N834), .Z(N835) );
  GTECH_OR2 C1354 ( .A(a1stg_op[4]), .B(N835), .Z(N836) );
  GTECH_OR2 C1355 ( .A(a1stg_op[3]), .B(N836), .Z(N837) );
  GTECH_OR2 C1356 ( .A(a1stg_op[2]), .B(N837), .Z(N838) );
  GTECH_OR2 C1357 ( .A(a1stg_op[1]), .B(N838), .Z(N839) );
  GTECH_OR2 C1358 ( .A(N75), .B(N839), .Z(N840) );
  GTECH_NOT I_133 ( .A(N840), .Z(N841) );
  GTECH_OR2 C1362 ( .A(a1stg_op[6]), .B(N72), .Z(N842) );
  GTECH_OR2 C1363 ( .A(a1stg_op[5]), .B(N842), .Z(N843) );
  GTECH_OR2 C1364 ( .A(a1stg_op[4]), .B(N843), .Z(N844) );
  GTECH_OR2 C1365 ( .A(a1stg_op[3]), .B(N844), .Z(N845) );
  GTECH_OR2 C1366 ( .A(a1stg_op[2]), .B(N845), .Z(N846) );
  GTECH_OR2 C1367 ( .A(N92), .B(N846), .Z(N847) );
  GTECH_OR2 C1368 ( .A(a1stg_op[0]), .B(N847), .Z(N848) );
  GTECH_NOT I_134 ( .A(N848), .Z(N849) );
  GTECH_OR2 C1372 ( .A(N73), .B(a1stg_op[7]), .Z(N850) );
  GTECH_OR2 C1373 ( .A(a1stg_op[5]), .B(N850), .Z(N851) );
  GTECH_OR2 C1374 ( .A(a1stg_op[4]), .B(N851), .Z(N852) );
  GTECH_OR2 C1375 ( .A(a1stg_op[3]), .B(N852), .Z(N853) );
  GTECH_OR2 C1376 ( .A(a1stg_op[2]), .B(N853), .Z(N854) );
  GTECH_OR2 C1377 ( .A(a1stg_op[1]), .B(N854), .Z(N855) );
  GTECH_OR2 C1378 ( .A(N75), .B(N855), .Z(N856) );
  GTECH_NOT I_135 ( .A(N856), .Z(N857) );
  GTECH_OR2 C1382 ( .A(N73), .B(a1stg_op[7]), .Z(N858) );
  GTECH_OR2 C1383 ( .A(a1stg_op[5]), .B(N858), .Z(N859) );
  GTECH_OR2 C1384 ( .A(a1stg_op[4]), .B(N859), .Z(N860) );
  GTECH_OR2 C1385 ( .A(a1stg_op[3]), .B(N860), .Z(N861) );
  GTECH_OR2 C1386 ( .A(a1stg_op[2]), .B(N861), .Z(N862) );
  GTECH_OR2 C1387 ( .A(N92), .B(N862), .Z(N863) );
  GTECH_OR2 C1388 ( .A(a1stg_op[0]), .B(N863), .Z(N864) );
  GTECH_NOT I_136 ( .A(N864), .Z(N865) );
  GTECH_OR2 C1393 ( .A(N73), .B(a1stg_op[7]), .Z(N866) );
  GTECH_OR2 C1394 ( .A(a1stg_op[5]), .B(N866), .Z(N867) );
  GTECH_OR2 C1395 ( .A(a1stg_op[4]), .B(N867), .Z(N868) );
  GTECH_OR2 C1396 ( .A(a1stg_op[3]), .B(N868), .Z(N869) );
  GTECH_OR2 C1397 ( .A(N109), .B(N869), .Z(N870) );
  GTECH_OR2 C1398 ( .A(a1stg_op[1]), .B(N870), .Z(N871) );
  GTECH_OR2 C1399 ( .A(N75), .B(N871), .Z(N872) );
  GTECH_NOT I_137 ( .A(N872), .Z(N873) );
  GTECH_OR2 C1404 ( .A(N73), .B(a1stg_op[7]), .Z(N874) );
  GTECH_OR2 C1405 ( .A(a1stg_op[5]), .B(N874), .Z(N875) );
  GTECH_OR2 C1406 ( .A(a1stg_op[4]), .B(N875), .Z(N876) );
  GTECH_OR2 C1407 ( .A(a1stg_op[3]), .B(N876), .Z(N877) );
  GTECH_OR2 C1408 ( .A(N109), .B(N877), .Z(N878) );
  GTECH_OR2 C1409 ( .A(N92), .B(N878), .Z(N879) );
  GTECH_OR2 C1410 ( .A(a1stg_op[0]), .B(N879), .Z(N880) );
  GTECH_NOT I_138 ( .A(N880), .Z(N881) );
  GTECH_OR2 C1416 ( .A(N73), .B(N72), .Z(N882) );
  GTECH_OR2 C1417 ( .A(a1stg_op[5]), .B(N882), .Z(N883) );
  GTECH_OR2 C1418 ( .A(a1stg_op[4]), .B(N883), .Z(N884) );
  GTECH_OR2 C1419 ( .A(a1stg_op[3]), .B(N884), .Z(N885) );
  GTECH_OR2 C1420 ( .A(N109), .B(N885), .Z(N886) );
  GTECH_OR2 C1421 ( .A(N92), .B(N886), .Z(N887) );
  GTECH_OR2 C1422 ( .A(a1stg_op[0]), .B(N887), .Z(N888) );
  GTECH_NOT I_139 ( .A(N888), .Z(N889) );
  GTECH_OR2 C1426 ( .A(N73), .B(a1stg_op[7]), .Z(N890) );
  GTECH_OR2 C1427 ( .A(a1stg_op[5]), .B(N890), .Z(N891) );
  GTECH_OR2 C1428 ( .A(a1stg_op[4]), .B(N891), .Z(N892) );
  GTECH_OR2 C1429 ( .A(a1stg_op[3]), .B(N892), .Z(N893) );
  GTECH_OR2 C1430 ( .A(a1stg_op[2]), .B(N893), .Z(N894) );
  GTECH_OR2 C1431 ( .A(a1stg_op[1]), .B(N894), .Z(N895) );
  GTECH_OR2 C1432 ( .A(N75), .B(N895), .Z(N896) );
  GTECH_NOT I_140 ( .A(N896), .Z(N897) );
  GTECH_OR2 C1436 ( .A(N73), .B(a1stg_op[7]), .Z(N898) );
  GTECH_OR2 C1437 ( .A(a1stg_op[5]), .B(N898), .Z(N899) );
  GTECH_OR2 C1438 ( .A(a1stg_op[4]), .B(N899), .Z(N900) );
  GTECH_OR2 C1439 ( .A(a1stg_op[3]), .B(N900), .Z(N901) );
  GTECH_OR2 C1440 ( .A(a1stg_op[2]), .B(N901), .Z(N902) );
  GTECH_OR2 C1441 ( .A(N92), .B(N902), .Z(N903) );
  GTECH_OR2 C1442 ( .A(a1stg_op[0]), .B(N903), .Z(N904) );
  GTECH_NOT I_141 ( .A(N904), .Z(N905) );
  GTECH_OR2 C1447 ( .A(N73), .B(a1stg_op[7]), .Z(N906) );
  GTECH_OR2 C1448 ( .A(a1stg_op[5]), .B(N906), .Z(N907) );
  GTECH_OR2 C1449 ( .A(a1stg_op[4]), .B(N907), .Z(N908) );
  GTECH_OR2 C1450 ( .A(a1stg_op[3]), .B(N908), .Z(N909) );
  GTECH_OR2 C1451 ( .A(N109), .B(N909), .Z(N910) );
  GTECH_OR2 C1452 ( .A(a1stg_op[1]), .B(N910), .Z(N911) );
  GTECH_OR2 C1453 ( .A(N75), .B(N911), .Z(N912) );
  GTECH_NOT I_142 ( .A(N912), .Z(N913) );
  GTECH_OR2 C1458 ( .A(N73), .B(a1stg_op[7]), .Z(N914) );
  GTECH_OR2 C1459 ( .A(a1stg_op[5]), .B(N914), .Z(N915) );
  GTECH_OR2 C1460 ( .A(a1stg_op[4]), .B(N915), .Z(N916) );
  GTECH_OR2 C1461 ( .A(a1stg_op[3]), .B(N916), .Z(N917) );
  GTECH_OR2 C1462 ( .A(N109), .B(N917), .Z(N918) );
  GTECH_OR2 C1463 ( .A(N92), .B(N918), .Z(N919) );
  GTECH_OR2 C1464 ( .A(a1stg_op[0]), .B(N919), .Z(N920) );
  GTECH_NOT I_143 ( .A(N920), .Z(N921) );
  GTECH_NOT I_144 ( .A(add_ctl_rst_l), .Z(reset) );
  GTECH_AND2 C1469 ( .A(a1stg_in1_exp_eq_0), .B(a1stg_sngopa[0]), .Z(
        a1stg_denorm_sng_in1) );
  GTECH_AND2 C1470 ( .A(a1stg_in1_exp_eq_0), .B(a1stg_dblopa[0]), .Z(
        a1stg_denorm_dbl_in1) );
  GTECH_AND2 C1471 ( .A(a1stg_in2_exp_eq_0), .B(a1stg_sngopa[0]), .Z(
        a1stg_denorm_sng_in2) );
  GTECH_AND2 C1472 ( .A(a1stg_in2_exp_eq_0), .B(a1stg_dblopa[0]), .Z(
        a1stg_denorm_dbl_in2) );
  GTECH_AND2 C1473 ( .A(N922), .B(a1stg_sngopa[0]), .Z(a1stg_norm_sng_in1) );
  GTECH_NOT I_145 ( .A(a1stg_in1_exp_eq_0), .Z(N922) );
  GTECH_AND2 C1475 ( .A(N922), .B(a1stg_dblopa[0]), .Z(a1stg_norm_dbl_in1) );
  GTECH_AND2 C1477 ( .A(N923), .B(a1stg_sngopa[0]), .Z(a1stg_norm_sng_in2) );
  GTECH_NOT I_146 ( .A(a1stg_in2_exp_eq_0), .Z(N923) );
  GTECH_AND2 C1479 ( .A(N923), .B(a1stg_dblopa[0]), .Z(a1stg_norm_dbl_in2) );
  GTECH_AND2 C1481 ( .A(N927), .B(a1stg_sngopa[1]), .Z(a1stg_snan_sng_in1) );
  GTECH_AND2 C1482 ( .A(N926), .B(a1stg_in1_53_32_neq_0), .Z(N927) );
  GTECH_AND2 C1483 ( .A(N924), .B(N925), .Z(N926) );
  GTECH_NOT I_147 ( .A(a1stg_in1_exp_neq_ffs), .Z(N924) );
  GTECH_NOT I_148 ( .A(a1stg_in1_54), .Z(N925) );
  GTECH_AND2 C1486 ( .A(N930), .B(a1stg_dblopa[1]), .Z(a1stg_snan_dbl_in1) );
  GTECH_AND2 C1487 ( .A(N929), .B(a1stg_in1_50_0_neq_0), .Z(N930) );
  GTECH_AND2 C1488 ( .A(N924), .B(N928), .Z(N929) );
  GTECH_NOT I_149 ( .A(a1stg_in1_51), .Z(N928) );
  GTECH_AND2 C1491 ( .A(N934), .B(a1stg_sngopa[1]), .Z(a1stg_snan_sng_in2) );
  GTECH_AND2 C1492 ( .A(N933), .B(a1stg_in2_53_32_neq_0), .Z(N934) );
  GTECH_AND2 C1493 ( .A(N931), .B(N932), .Z(N933) );
  GTECH_NOT I_150 ( .A(a1stg_in2_exp_neq_ffs), .Z(N931) );
  GTECH_NOT I_151 ( .A(a1stg_in2_54), .Z(N932) );
  GTECH_AND2 C1496 ( .A(N937), .B(a1stg_dblopa[1]), .Z(a1stg_snan_dbl_in2) );
  GTECH_AND2 C1497 ( .A(N936), .B(a1stg_in2_50_0_neq_0), .Z(N937) );
  GTECH_AND2 C1498 ( .A(N931), .B(N935), .Z(N936) );
  GTECH_NOT I_152 ( .A(a1stg_in2_51), .Z(N935) );
  GTECH_AND2 C1501 ( .A(N938), .B(a1stg_sngopa[1]), .Z(a1stg_qnan_sng_in1) );
  GTECH_AND2 C1502 ( .A(N924), .B(a1stg_in1_54), .Z(N938) );
  GTECH_AND2 C1504 ( .A(N939), .B(a1stg_dblopa[1]), .Z(a1stg_qnan_dbl_in1) );
  GTECH_AND2 C1505 ( .A(N924), .B(a1stg_in1_51), .Z(N939) );
  GTECH_AND2 C1507 ( .A(N940), .B(a1stg_sngopa[1]), .Z(a1stg_qnan_sng_in2) );
  GTECH_AND2 C1508 ( .A(N931), .B(a1stg_in2_54), .Z(N940) );
  GTECH_AND2 C1510 ( .A(N941), .B(a1stg_dblopa[1]), .Z(a1stg_qnan_dbl_in2) );
  GTECH_AND2 C1511 ( .A(N931), .B(a1stg_in2_51), .Z(N941) );
  GTECH_OR2 C1513 ( .A(a1stg_snan_sng_in1), .B(a1stg_snan_dbl_in1), .Z(
        a1stg_snan_in1) );
  GTECH_OR2 C1514 ( .A(a1stg_snan_sng_in2), .B(a1stg_snan_dbl_in2), .Z(
        a1stg_snan_in2) );
  GTECH_OR2 C1515 ( .A(a1stg_qnan_sng_in1), .B(a1stg_qnan_dbl_in1), .Z(
        a1stg_qnan_in1) );
  GTECH_OR2 C1516 ( .A(a1stg_qnan_sng_in2), .B(a1stg_qnan_dbl_in2), .Z(
        a1stg_qnan_in2) );
  GTECH_AND2 C1517 ( .A(N943), .B(a1stg_sngopa[2]), .Z(a1stg_nan_sng_in1) );
  GTECH_AND2 C1518 ( .A(N924), .B(N942), .Z(N943) );
  GTECH_OR2 C1520 ( .A(a1stg_in1_54), .B(a1stg_in1_53_32_neq_0), .Z(N942) );
  GTECH_AND2 C1521 ( .A(N945), .B(a1stg_dblopa[2]), .Z(a1stg_nan_dbl_in1) );
  GTECH_AND2 C1522 ( .A(N924), .B(N944), .Z(N945) );
  GTECH_OR2 C1524 ( .A(a1stg_in1_51), .B(a1stg_in1_50_0_neq_0), .Z(N944) );
  GTECH_AND2 C1525 ( .A(N947), .B(a1stg_sngopa[2]), .Z(a1stg_nan_sng_in2) );
  GTECH_AND2 C1526 ( .A(N931), .B(N946), .Z(N947) );
  GTECH_OR2 C1528 ( .A(a1stg_in2_54), .B(a1stg_in2_53_32_neq_0), .Z(N946) );
  GTECH_AND2 C1529 ( .A(N949), .B(a1stg_dblopa[2]), .Z(a1stg_nan_dbl_in2) );
  GTECH_AND2 C1530 ( .A(N931), .B(N948), .Z(N949) );
  GTECH_OR2 C1532 ( .A(a1stg_in2_51), .B(a1stg_in2_50_0_neq_0), .Z(N948) );
  GTECH_OR2 C1533 ( .A(a1stg_nan_sng_in1), .B(a1stg_nan_dbl_in1), .Z(
        a1stg_nan_in1) );
  GTECH_OR2 C1534 ( .A(a1stg_nan_sng_in2), .B(a1stg_nan_dbl_in2), .Z(
        a1stg_nan_in2) );
  GTECH_OR2 C1535 ( .A(a1stg_nan_in1), .B(a1stg_nan_in2), .Z(a1stg_nan_in) );
  GTECH_AND2 C1536 ( .A(a1stg_nan_in1), .B(a1stg_nan_in2), .Z(a1stg_2nan_in)
         );
  GTECH_AND2 C1537 ( .A(N952), .B(a1stg_sngopa[2]), .Z(a1stg_inf_sng_in1) );
  GTECH_AND2 C1538 ( .A(N950), .B(N951), .Z(N952) );
  GTECH_AND2 C1539 ( .A(N924), .B(N925), .Z(N950) );
  GTECH_NOT I_153 ( .A(a1stg_in1_53_32_neq_0), .Z(N951) );
  GTECH_AND2 C1543 ( .A(N955), .B(a1stg_dblopa[2]), .Z(a1stg_inf_dbl_in1) );
  GTECH_AND2 C1544 ( .A(N953), .B(N954), .Z(N955) );
  GTECH_AND2 C1545 ( .A(N924), .B(N928), .Z(N953) );
  GTECH_NOT I_154 ( .A(a1stg_in1_50_0_neq_0), .Z(N954) );
  GTECH_AND2 C1549 ( .A(N958), .B(a1stg_sngopa[2]), .Z(a1stg_inf_sng_in2) );
  GTECH_AND2 C1550 ( .A(N956), .B(N957), .Z(N958) );
  GTECH_AND2 C1551 ( .A(N931), .B(N932), .Z(N956) );
  GTECH_NOT I_155 ( .A(a1stg_in2_53_32_neq_0), .Z(N957) );
  GTECH_AND2 C1555 ( .A(N961), .B(a1stg_dblopa[2]), .Z(a1stg_inf_dbl_in2) );
  GTECH_AND2 C1556 ( .A(N959), .B(N960), .Z(N961) );
  GTECH_AND2 C1557 ( .A(N931), .B(N935), .Z(N959) );
  GTECH_NOT I_156 ( .A(a1stg_in2_50_0_neq_0), .Z(N960) );
  GTECH_OR2 C1561 ( .A(a1stg_inf_sng_in1), .B(a1stg_inf_dbl_in1), .Z(
        a1stg_inf_in1) );
  GTECH_OR2 C1562 ( .A(a1stg_inf_sng_in2), .B(a1stg_inf_dbl_in2), .Z(
        a1stg_inf_in2) );
  GTECH_AND2 C1563 ( .A(a1stg_inf_in1), .B(a1stg_inf_in2), .Z(a1stg_2inf_in)
         );
  GTECH_AND2 C1564 ( .A(N924), .B(a1stg_sngopa[3]), .Z(a1stg_infnan_sng_in1)
         );
  GTECH_AND2 C1566 ( .A(N924), .B(a1stg_dblopa[3]), .Z(a1stg_infnan_dbl_in1)
         );
  GTECH_AND2 C1568 ( .A(N931), .B(a1stg_sngopa[3]), .Z(a1stg_infnan_sng_in2)
         );
  GTECH_AND2 C1570 ( .A(N931), .B(a1stg_dblopa[3]), .Z(a1stg_infnan_dbl_in2)
         );
  GTECH_OR2 C1572 ( .A(a1stg_infnan_sng_in1), .B(a1stg_infnan_dbl_in1), .Z(
        a1stg_infnan_in1) );
  GTECH_OR2 C1573 ( .A(a1stg_infnan_sng_in2), .B(a1stg_infnan_dbl_in2), .Z(
        a1stg_infnan_in2) );
  GTECH_OR2 C1574 ( .A(a1stg_infnan_in1), .B(a1stg_infnan_in2), .Z(
        a1stg_infnan_in) );
  GTECH_AND2 C1575 ( .A(N973), .B(N960), .Z(a1stg_2zero_in) );
  GTECH_AND2 C1576 ( .A(N972), .B(N935), .Z(N973) );
  GTECH_AND2 C1577 ( .A(N970), .B(N971), .Z(N972) );
  GTECH_AND2 C1578 ( .A(N968), .B(N969), .Z(N970) );
  GTECH_AND2 C1579 ( .A(N967), .B(a1stg_in2_exp_eq_0), .Z(N968) );
  GTECH_AND2 C1580 ( .A(N966), .B(N954), .Z(N967) );
  GTECH_AND2 C1581 ( .A(N965), .B(N928), .Z(N966) );
  GTECH_AND2 C1582 ( .A(N963), .B(N964), .Z(N965) );
  GTECH_AND2 C1583 ( .A(a1stg_in1_exp_eq_0), .B(N962), .Z(N963) );
  GTECH_OR2 C1584 ( .A(N925), .B(a1stg_dblopa[3]), .Z(N962) );
  GTECH_OR2 C1586 ( .A(N951), .B(a1stg_dblopa[3]), .Z(N964) );
  GTECH_OR2 C1590 ( .A(N932), .B(a1stg_dblopa[3]), .Z(N969) );
  GTECH_OR2 C1592 ( .A(N957), .B(a1stg_dblopa[3]), .Z(N971) );
  GTECH_AND2 C1596 ( .A(N974), .B(N975), .Z(a1stg_step) );
  GTECH_NOT I_157 ( .A(fixtosd_hold), .Z(N974) );
  GTECH_NOT I_158 ( .A(a6stg_hold), .Z(N975) );
  GTECH_AND2 C1599 ( .A(inq_add), .B(inq_op[7]), .Z(a1stg_op_in[7]) );
  GTECH_AND2 C1600 ( .A(inq_add), .B(inq_op[6]), .Z(a1stg_op_in[6]) );
  GTECH_AND2 C1601 ( .A(inq_add), .B(inq_op[5]), .Z(a1stg_op_in[5]) );
  GTECH_AND2 C1602 ( .A(inq_add), .B(inq_op[4]), .Z(a1stg_op_in[4]) );
  GTECH_AND2 C1603 ( .A(inq_add), .B(inq_op[3]), .Z(a1stg_op_in[3]) );
  GTECH_AND2 C1604 ( .A(inq_add), .B(inq_op[2]), .Z(a1stg_op_in[2]) );
  GTECH_AND2 C1605 ( .A(inq_add), .B(inq_op[1]), .Z(a1stg_op_in[1]) );
  GTECH_AND2 C1606 ( .A(inq_add), .B(inq_op[0]), .Z(a1stg_op_in[0]) );
  GTECH_OR2 C1607 ( .A(N991), .B(N702), .Z(a1stg_opdec[34]) );
  GTECH_OR2 C1608 ( .A(N990), .B(N694), .Z(N991) );
  GTECH_OR2 C1609 ( .A(N989), .B(N686), .Z(N990) );
  GTECH_OR2 C1610 ( .A(N988), .B(N678), .Z(N989) );
  GTECH_OR2 C1611 ( .A(N987), .B(N670), .Z(N988) );
  GTECH_OR2 C1612 ( .A(N986), .B(N662), .Z(N987) );
  GTECH_OR2 C1613 ( .A(N985), .B(N654), .Z(N986) );
  GTECH_OR2 C1614 ( .A(N984), .B(N646), .Z(N985) );
  GTECH_OR2 C1615 ( .A(N983), .B(N638), .Z(N984) );
  GTECH_OR2 C1616 ( .A(N982), .B(N630), .Z(N983) );
  GTECH_OR2 C1617 ( .A(N981), .B(N622), .Z(N982) );
  GTECH_OR2 C1618 ( .A(N980), .B(N614), .Z(N981) );
  GTECH_OR2 C1619 ( .A(N979), .B(N606), .Z(N980) );
  GTECH_OR2 C1620 ( .A(N978), .B(N598), .Z(N979) );
  GTECH_OR2 C1621 ( .A(N977), .B(N590), .Z(N978) );
  GTECH_OR2 C1622 ( .A(N976), .B(N582), .Z(N977) );
  GTECH_OR2 C1623 ( .A(N566), .B(N574), .Z(N976) );
  GTECH_OR2 C1624 ( .A(N994), .B(N214), .Z(a1stg_opdec[33]) );
  GTECH_OR2 C1625 ( .A(N993), .B(N206), .Z(N994) );
  GTECH_OR2 C1626 ( .A(N992), .B(N198), .Z(N993) );
  GTECH_OR2 C1627 ( .A(N182), .B(N190), .Z(N992) );
  GTECH_OR2 C1628 ( .A(N997), .B(N254), .Z(a1stg_opdec[32]) );
  GTECH_OR2 C1629 ( .A(N996), .B(N246), .Z(N997) );
  GTECH_OR2 C1630 ( .A(N995), .B(N238), .Z(N996) );
  GTECH_OR2 C1631 ( .A(N222), .B(N230), .Z(N995) );
  GTECH_OR2 C1632 ( .A(N262), .B(N270), .Z(a1stg_opdec[31]) );
  GTECH_OR2 C1633 ( .A(N278), .B(N286), .Z(a1stg_opdec[30]) );
  GTECH_NOT I_159 ( .A(N998), .Z(a1stg_intlngop) );
  GTECH_OR2 C1635 ( .A(a1stg_sngopa[3]), .B(a1stg_dblop), .Z(N998) );
  GTECH_OR2 C1636 ( .A(N1000), .B(N921), .Z(a1stg_opdec[29]) );
  GTECH_OR2 C1637 ( .A(N999), .B(N913), .Z(N1000) );
  GTECH_OR2 C1638 ( .A(N897), .B(N905), .Z(N999) );
  GTECH_OR2 C1639 ( .A(N783), .B(N791), .Z(a1stg_opdec[28]) );
  GTECH_OR2 C1640 ( .A(N841), .B(N849), .Z(a1stg_fsdtox) );
  GTECH_OR2 C1641 ( .A(N711), .B(N719), .Z(a1stg_fcmpesd) );
  GTECH_OR2 C1642 ( .A(N727), .B(N735), .Z(a1stg_fcmpsd) );
  GTECH_OR2 C1643 ( .A(N1003), .B(N889), .Z(a1stg_opdec_24_21[3]) );
  GTECH_OR2 C1644 ( .A(N1002), .B(N881), .Z(N1003) );
  GTECH_OR2 C1645 ( .A(N1001), .B(N873), .Z(N1002) );
  GTECH_OR2 C1646 ( .A(N857), .B(N865), .Z(N1001) );
  GTECH_OR2 C1647 ( .A(N294), .B(N302), .Z(a1stg_opdec_24_21[2]) );
  GTECH_OR2 C1648 ( .A(N310), .B(N318), .Z(a1stg_opdec_24_21[1]) );
  GTECH_OR2 C1649 ( .A(N1005), .B(N823), .Z(a1stg_fsdtoix) );
  GTECH_OR2 C1650 ( .A(N1004), .B(N815), .Z(N1005) );
  GTECH_OR2 C1651 ( .A(N799), .B(N807), .Z(N1004) );
  GTECH_OR2 C1652 ( .A(N1007), .B(N767), .Z(a1stg_fixtosd) );
  GTECH_OR2 C1653 ( .A(N1006), .B(N759), .Z(N1007) );
  GTECH_OR2 C1654 ( .A(N743), .B(N751), .Z(N1006) );
  GTECH_OR2 C1655 ( .A(N1010), .B(N358), .Z(a1stg_opdec_19_11[3]) );
  GTECH_OR2 C1656 ( .A(N1009), .B(N350), .Z(N1010) );
  GTECH_OR2 C1657 ( .A(N1008), .B(N342), .Z(N1009) );
  GTECH_OR2 C1658 ( .A(N326), .B(N334), .Z(N1008) );
  GTECH_OR2 C1659 ( .A(N1012), .B(N390), .Z(a1stg_opdec_9_0[9]) );
  GTECH_OR2 C1660 ( .A(N1011), .B(N382), .Z(N1012) );
  GTECH_OR2 C1661 ( .A(N366), .B(N374), .Z(N1011) );
  GTECH_OR2 C1662 ( .A(N1017), .B(N446), .Z(a1stg_opdec_9_0[8]) );
  GTECH_OR2 C1663 ( .A(N1016), .B(N438), .Z(N1017) );
  GTECH_OR2 C1664 ( .A(N1015), .B(N430), .Z(N1016) );
  GTECH_OR2 C1665 ( .A(N1014), .B(N422), .Z(N1015) );
  GTECH_OR2 C1666 ( .A(N1013), .B(N414), .Z(N1014) );
  GTECH_OR2 C1667 ( .A(N398), .B(N406), .Z(N1013) );
  GTECH_OR2 C1668 ( .A(N1018), .B(N470), .Z(a1stg_opdec_9_0[7]) );
  GTECH_OR2 C1669 ( .A(N454), .B(N462), .Z(N1018) );
  GTECH_OR2 C1670 ( .A(N1019), .B(N494), .Z(a1stg_opdec_9_0[6]) );
  GTECH_OR2 C1671 ( .A(N478), .B(N486), .Z(N1019) );
  GTECH_OR2 C1672 ( .A(N502), .B(N510), .Z(a1stg_faddsubs) );
  GTECH_OR2 C1673 ( .A(N518), .B(N526), .Z(a1stg_faddsubd) );
  GTECH_OR2 C1674 ( .A(N534), .B(N542), .Z(a1stg_opdec_9_0_2) );
  GTECH_OR2 C1675 ( .A(N550), .B(N558), .Z(a1stg_opdec_9_0_1) );
  GTECH_AND2 C1676 ( .A(a2stg_opdec_9_0[7]), .B(N1024), .Z(fixtosd_hold) );
  GTECH_NOT I_160 ( .A(N1023), .Z(N1024) );
  GTECH_AND2 C1678 ( .A(N1021), .B(N1022), .Z(N1023) );
  GTECH_AND2 C1679 ( .A(N1020), .B(N75), .Z(N1021) );
  GTECH_AND2 C1680 ( .A(a1stg_op[7]), .B(N92), .Z(N1020) );
  GTECH_OR2 C1683 ( .A(a1stg_op[2]), .B(N73), .Z(N1022) );
  GTECH_AND2 C1685 ( .A(N974), .B(a1stg_dblop), .Z(a2stg_opdec_in[30]) );
  GTECH_AND2 C1687 ( .A(N974), .B(a1stg_opdec[34]), .Z(a2stg_opdec_in[29]) );
  GTECH_AND2 C1689 ( .A(N974), .B(a1stg_opdec[33]), .Z(a2stg_opdec_in[28]) );
  GTECH_AND2 C1691 ( .A(N974), .B(a1stg_opdec[32]), .Z(a2stg_opdec_in[27]) );
  GTECH_AND2 C1693 ( .A(N974), .B(a1stg_opdec[31]), .Z(a2stg_opdec_in[26]) );
  GTECH_AND2 C1695 ( .A(N974), .B(a1stg_opdec[30]), .Z(a2stg_opdec_in[25]) );
  GTECH_AND2 C1697 ( .A(N974), .B(a1stg_opdec[29]), .Z(a2stg_opdec_in[24]) );
  GTECH_AND2 C1699 ( .A(N974), .B(a1stg_opdec[28]), .Z(a2stg_opdec_in[23]) );
  GTECH_AND2 C1701 ( .A(N974), .B(a1stg_opdec_24_21[3]), .Z(a2stg_opdec_in[22]) );
  GTECH_AND2 C1703 ( .A(N974), .B(a1stg_opdec_24_21[2]), .Z(a2stg_opdec_in[21]) );
  GTECH_AND2 C1705 ( .A(N974), .B(a1stg_opdec_24_21[1]), .Z(a2stg_opdec_in[20]) );
  GTECH_AND2 C1707 ( .A(N974), .B(a1stg_fsdtoix), .Z(a2stg_opdec_in[19]) );
  GTECH_AND2 C1709 ( .A(N974), .B(N168), .Z(a2stg_opdec_in[18]) );
  GTECH_AND2 C1711 ( .A(N974), .B(N83), .Z(a2stg_opdec_in[17]) );
  GTECH_AND2 C1713 ( .A(N974), .B(N91), .Z(a2stg_opdec_in[16]) );
  GTECH_AND2 C1715 ( .A(N974), .B(N100), .Z(a2stg_opdec_in[15]) );
  GTECH_AND2 C1717 ( .A(N974), .B(N108), .Z(a2stg_opdec_in[14]) );
  GTECH_AND2 C1719 ( .A(N974), .B(a1stg_opdec_19_11[3]), .Z(a2stg_opdec_in[13]) );
  GTECH_AND2 C1721 ( .A(N974), .B(N117), .Z(a2stg_opdec_in[12]) );
  GTECH_AND2 C1723 ( .A(N974), .B(N126), .Z(a2stg_opdec_in[11]) );
  GTECH_AND2 C1725 ( .A(N974), .B(N134), .Z(a2stg_opdec_in[10]) );
  GTECH_AND2 C1727 ( .A(N974), .B(a1stg_opdec_9_0[9]), .Z(a2stg_opdec_in[9])
         );
  GTECH_AND2 C1729 ( .A(N974), .B(a1stg_opdec_9_0[8]), .Z(a2stg_opdec_in[8])
         );
  GTECH_AND2 C1731 ( .A(N974), .B(a1stg_opdec_9_0[7]), .Z(a2stg_opdec_in[7])
         );
  GTECH_AND2 C1733 ( .A(N974), .B(a1stg_opdec_9_0[6]), .Z(a2stg_opdec_in[6])
         );
  GTECH_AND2 C1735 ( .A(N974), .B(a1stg_faddsubs), .Z(a2stg_opdec_in[5]) );
  GTECH_AND2 C1737 ( .A(N974), .B(a1stg_faddsubd), .Z(a2stg_opdec_in[4]) );
  GTECH_AND2 C1739 ( .A(N974), .B(N775), .Z(a2stg_opdec_in[3]) );
  GTECH_AND2 C1741 ( .A(N974), .B(a1stg_opdec_9_0_2), .Z(a2stg_opdec_in[2]) );
  GTECH_AND2 C1743 ( .A(N974), .B(a1stg_opdec_9_0_1), .Z(a2stg_opdec_in[1]) );
  GTECH_AND2 C1745 ( .A(N974), .B(N142), .Z(a2stg_opdec_in[0]) );
  GTECH_OR2 C1747 ( .A(N1025), .B(N1027), .Z(a4stg_rnd_mode_in[1]) );
  GTECH_AND2 C1748 ( .A(a3stg_opdec_9_0[8]), .B(a3stg_rnd_mode[1]), .Z(N1025)
         );
  GTECH_AND2 C1749 ( .A(N1026), .B(a4stg_rnd_mode2[1]), .Z(N1027) );
  GTECH_NOT I_161 ( .A(a3stg_opdec_9_0[8]), .Z(N1026) );
  GTECH_OR2 C1751 ( .A(N1028), .B(N1029), .Z(a4stg_rnd_mode_in[0]) );
  GTECH_AND2 C1752 ( .A(a3stg_opdec_9_0[8]), .B(a3stg_rnd_mode[0]), .Z(N1028)
         );
  GTECH_AND2 C1753 ( .A(N1026), .B(a4stg_rnd_mode2[0]), .Z(N1029) );
  GTECH_OR2 C1755 ( .A(N1030), .B(N1034), .Z(a6stg_opdec_in[34]) );
  GTECH_AND2 C1756 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec[34]), .Z(N1030) );
  GTECH_AND2 C1757 ( .A(N1033), .B(a4stg_opdec[34]), .Z(N1034) );
  GTECH_AND2 C1758 ( .A(N1031), .B(N1032), .Z(N1033) );
  GTECH_NOT I_162 ( .A(a4stg_opdec_7_0[7]), .Z(N1031) );
  GTECH_NOT I_163 ( .A(a5stg_fixtos_fxtod), .Z(N1032) );
  GTECH_OR2 C1761 ( .A(N1035), .B(N1038), .Z(a6stg_opdec_in[33]) );
  GTECH_AND2 C1762 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec[33]), .Z(N1035) );
  GTECH_AND2 C1763 ( .A(N1037), .B(a4stg_opdec[33]), .Z(N1038) );
  GTECH_AND2 C1764 ( .A(N1036), .B(N1032), .Z(N1037) );
  GTECH_NOT I_164 ( .A(a4stg_opdec_7_0[7]), .Z(N1036) );
  GTECH_OR2 C1767 ( .A(N1039), .B(N1042), .Z(a6stg_opdec_in[32]) );
  GTECH_AND2 C1768 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec[32]), .Z(N1039) );
  GTECH_AND2 C1769 ( .A(N1041), .B(a4stg_opdec[32]), .Z(N1042) );
  GTECH_AND2 C1770 ( .A(N1040), .B(N1032), .Z(N1041) );
  GTECH_NOT I_165 ( .A(a4stg_opdec_7_0[7]), .Z(N1040) );
  GTECH_OR2 C1773 ( .A(N1043), .B(N1046), .Z(a6stg_opdec_in[31]) );
  GTECH_AND2 C1774 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec[31]), .Z(N1043) );
  GTECH_AND2 C1775 ( .A(N1045), .B(a4stg_opdec[31]), .Z(N1046) );
  GTECH_AND2 C1776 ( .A(N1044), .B(N1032), .Z(N1045) );
  GTECH_NOT I_166 ( .A(a4stg_opdec_7_0[7]), .Z(N1044) );
  GTECH_OR2 C1779 ( .A(N1047), .B(N1050), .Z(a6stg_opdec_in[30]) );
  GTECH_AND2 C1780 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec[30]), .Z(N1047) );
  GTECH_AND2 C1781 ( .A(N1049), .B(a4stg_opdec[30]), .Z(N1050) );
  GTECH_AND2 C1782 ( .A(N1048), .B(N1032), .Z(N1049) );
  GTECH_NOT I_167 ( .A(a4stg_opdec_7_0[7]), .Z(N1048) );
  GTECH_OR2 C1785 ( .A(N1051), .B(N1054), .Z(a6stg_opdec_in_9) );
  GTECH_AND2 C1786 ( .A(a5stg_fixtos_fxtod), .B(a5stg_opdec_9), .Z(N1051) );
  GTECH_AND2 C1787 ( .A(N1053), .B(a4stg_fcmpop), .Z(N1054) );
  GTECH_AND2 C1788 ( .A(N1052), .B(N1032), .Z(N1053) );
  GTECH_NOT I_168 ( .A(a4stg_opdec_7_0[7]), .Z(N1052) );
  GTECH_NOT I_169 ( .A(reset), .Z(N0) );
  GTECH_OR2 C1792 ( .A(N1063), .B(N1066), .Z(a6stg_fadd_in) );
  GTECH_OR2 C1793 ( .A(N1057), .B(N1062), .Z(N1063) );
  GTECH_AND2 C1794 ( .A(N1056), .B(a5stg_opdec[34]), .Z(N1057) );
  GTECH_AND2 C1795 ( .A(N1055), .B(N0), .Z(N1056) );
  GTECH_AND2 C1796 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1055) );
  GTECH_AND2 C1797 ( .A(N1061), .B(a4stg_opdec[34]), .Z(N1062) );
  GTECH_AND2 C1798 ( .A(N1060), .B(N0), .Z(N1061) );
  GTECH_AND2 C1799 ( .A(N1059), .B(a6stg_step), .Z(N1060) );
  GTECH_AND2 C1800 ( .A(N1058), .B(N1032), .Z(N1059) );
  GTECH_NOT I_170 ( .A(a4stg_opdec_7_0[7]), .Z(N1058) );
  GTECH_AND2 C1803 ( .A(N1065), .B(a6stg_opdec[34]), .Z(N1066) );
  GTECH_AND2 C1804 ( .A(N1064), .B(N0), .Z(N1065) );
  GTECH_NOT I_171 ( .A(a6stg_step), .Z(N1064) );
  GTECH_OR2 C1806 ( .A(N1071), .B(N1073), .Z(add_id_out_in[9]) );
  GTECH_OR2 C1807 ( .A(N1068), .B(N1070), .Z(N1071) );
  GTECH_AND2 C1808 ( .A(N1067), .B(a4stg_id[9]), .Z(N1068) );
  GTECH_AND2 C1809 ( .A(N1032), .B(a6stg_step), .Z(N1067) );
  GTECH_AND2 C1811 ( .A(N1069), .B(a5stg_id[9]), .Z(N1070) );
  GTECH_AND2 C1812 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1069) );
  GTECH_AND2 C1813 ( .A(N1072), .B(add_id_out[9]), .Z(N1073) );
  GTECH_NOT I_172 ( .A(a6stg_step), .Z(N1072) );
  GTECH_OR2 C1815 ( .A(N1078), .B(N1080), .Z(add_id_out_in[8]) );
  GTECH_OR2 C1816 ( .A(N1075), .B(N1077), .Z(N1078) );
  GTECH_AND2 C1817 ( .A(N1074), .B(a4stg_id[8]), .Z(N1075) );
  GTECH_AND2 C1818 ( .A(N1032), .B(a6stg_step), .Z(N1074) );
  GTECH_AND2 C1820 ( .A(N1076), .B(a5stg_id[8]), .Z(N1077) );
  GTECH_AND2 C1821 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1076) );
  GTECH_AND2 C1822 ( .A(N1079), .B(add_id_out[8]), .Z(N1080) );
  GTECH_NOT I_173 ( .A(a6stg_step), .Z(N1079) );
  GTECH_OR2 C1824 ( .A(N1085), .B(N1087), .Z(add_id_out_in[7]) );
  GTECH_OR2 C1825 ( .A(N1082), .B(N1084), .Z(N1085) );
  GTECH_AND2 C1826 ( .A(N1081), .B(a4stg_id[7]), .Z(N1082) );
  GTECH_AND2 C1827 ( .A(N1032), .B(a6stg_step), .Z(N1081) );
  GTECH_AND2 C1829 ( .A(N1083), .B(a5stg_id[7]), .Z(N1084) );
  GTECH_AND2 C1830 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1083) );
  GTECH_AND2 C1831 ( .A(N1086), .B(add_id_out[7]), .Z(N1087) );
  GTECH_NOT I_174 ( .A(a6stg_step), .Z(N1086) );
  GTECH_OR2 C1833 ( .A(N1092), .B(N1094), .Z(add_id_out_in[6]) );
  GTECH_OR2 C1834 ( .A(N1089), .B(N1091), .Z(N1092) );
  GTECH_AND2 C1835 ( .A(N1088), .B(a4stg_id[6]), .Z(N1089) );
  GTECH_AND2 C1836 ( .A(N1032), .B(a6stg_step), .Z(N1088) );
  GTECH_AND2 C1838 ( .A(N1090), .B(a5stg_id[6]), .Z(N1091) );
  GTECH_AND2 C1839 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1090) );
  GTECH_AND2 C1840 ( .A(N1093), .B(add_id_out[6]), .Z(N1094) );
  GTECH_NOT I_175 ( .A(a6stg_step), .Z(N1093) );
  GTECH_OR2 C1842 ( .A(N1099), .B(N1101), .Z(add_id_out_in[5]) );
  GTECH_OR2 C1843 ( .A(N1096), .B(N1098), .Z(N1099) );
  GTECH_AND2 C1844 ( .A(N1095), .B(a4stg_id[5]), .Z(N1096) );
  GTECH_AND2 C1845 ( .A(N1032), .B(a6stg_step), .Z(N1095) );
  GTECH_AND2 C1847 ( .A(N1097), .B(a5stg_id[5]), .Z(N1098) );
  GTECH_AND2 C1848 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1097) );
  GTECH_AND2 C1849 ( .A(N1100), .B(add_id_out[5]), .Z(N1101) );
  GTECH_NOT I_176 ( .A(a6stg_step), .Z(N1100) );
  GTECH_OR2 C1851 ( .A(N1106), .B(N1108), .Z(add_id_out_in[4]) );
  GTECH_OR2 C1852 ( .A(N1103), .B(N1105), .Z(N1106) );
  GTECH_AND2 C1853 ( .A(N1102), .B(a4stg_id[4]), .Z(N1103) );
  GTECH_AND2 C1854 ( .A(N1032), .B(a6stg_step), .Z(N1102) );
  GTECH_AND2 C1856 ( .A(N1104), .B(a5stg_id[4]), .Z(N1105) );
  GTECH_AND2 C1857 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1104) );
  GTECH_AND2 C1858 ( .A(N1107), .B(add_id_out[4]), .Z(N1108) );
  GTECH_NOT I_177 ( .A(a6stg_step), .Z(N1107) );
  GTECH_OR2 C1860 ( .A(N1113), .B(N1115), .Z(add_id_out_in[3]) );
  GTECH_OR2 C1861 ( .A(N1110), .B(N1112), .Z(N1113) );
  GTECH_AND2 C1862 ( .A(N1109), .B(a4stg_id[3]), .Z(N1110) );
  GTECH_AND2 C1863 ( .A(N1032), .B(a6stg_step), .Z(N1109) );
  GTECH_AND2 C1865 ( .A(N1111), .B(a5stg_id[3]), .Z(N1112) );
  GTECH_AND2 C1866 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1111) );
  GTECH_AND2 C1867 ( .A(N1114), .B(add_id_out[3]), .Z(N1115) );
  GTECH_NOT I_178 ( .A(a6stg_step), .Z(N1114) );
  GTECH_OR2 C1869 ( .A(N1120), .B(N1122), .Z(add_id_out_in[2]) );
  GTECH_OR2 C1870 ( .A(N1117), .B(N1119), .Z(N1120) );
  GTECH_AND2 C1871 ( .A(N1116), .B(a4stg_id[2]), .Z(N1117) );
  GTECH_AND2 C1872 ( .A(N1032), .B(a6stg_step), .Z(N1116) );
  GTECH_AND2 C1874 ( .A(N1118), .B(a5stg_id[2]), .Z(N1119) );
  GTECH_AND2 C1875 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1118) );
  GTECH_AND2 C1876 ( .A(N1121), .B(add_id_out[2]), .Z(N1122) );
  GTECH_NOT I_179 ( .A(a6stg_step), .Z(N1121) );
  GTECH_OR2 C1878 ( .A(N1127), .B(N1129), .Z(add_id_out_in[1]) );
  GTECH_OR2 C1879 ( .A(N1124), .B(N1126), .Z(N1127) );
  GTECH_AND2 C1880 ( .A(N1123), .B(a4stg_id[1]), .Z(N1124) );
  GTECH_AND2 C1881 ( .A(N1032), .B(a6stg_step), .Z(N1123) );
  GTECH_AND2 C1883 ( .A(N1125), .B(a5stg_id[1]), .Z(N1126) );
  GTECH_AND2 C1884 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1125) );
  GTECH_AND2 C1885 ( .A(N1128), .B(add_id_out[1]), .Z(N1129) );
  GTECH_NOT I_180 ( .A(a6stg_step), .Z(N1128) );
  GTECH_OR2 C1887 ( .A(N1134), .B(N1136), .Z(add_id_out_in[0]) );
  GTECH_OR2 C1888 ( .A(N1131), .B(N1133), .Z(N1134) );
  GTECH_AND2 C1889 ( .A(N1130), .B(a4stg_id[0]), .Z(N1131) );
  GTECH_AND2 C1890 ( .A(N1032), .B(a6stg_step), .Z(N1130) );
  GTECH_AND2 C1892 ( .A(N1132), .B(a5stg_id[0]), .Z(N1133) );
  GTECH_AND2 C1893 ( .A(a5stg_fixtos_fxtod), .B(a6stg_step), .Z(N1132) );
  GTECH_AND2 C1894 ( .A(N1135), .B(add_id_out[0]), .Z(N1136) );
  GTECH_NOT I_181 ( .A(a6stg_step), .Z(N1135) );
  GTECH_AND2 C1896 ( .A(a4stg_fcmpop), .B(a4stg_fcc[1]), .Z(add_fcc_out_in[1])
         );
  GTECH_AND2 C1897 ( .A(a4stg_fcmpop), .B(a4stg_fcc[0]), .Z(add_fcc_out_in[0])
         );
  GTECH_AND2 C1898 ( .A(a6stg_opdec[34]), .B(N1137), .Z(a6stg_hold) );
  GTECH_NOT I_182 ( .A(add_dest_rdy), .Z(N1137) );
  GTECH_NOT I_183 ( .A(a6stg_hold), .Z(a6stg_step) );
  GTECH_OR2 C1901 ( .A(N1141), .B(a6stg_opdec[34]), .Z(add_pipe_active_in) );
  GTECH_OR2 C1902 ( .A(N1140), .B(a5stg_opdec[34]), .Z(N1141) );
  GTECH_OR2 C1903 ( .A(N1139), .B(a4stg_opdec[34]), .Z(N1140) );
  GTECH_OR2 C1904 ( .A(N1138), .B(a3stg_opdec[34]), .Z(N1139) );
  GTECH_OR2 C1905 ( .A(a1stg_opdec[34]), .B(a2stg_opdec[34]), .Z(N1138) );
  GTECH_AND2 C1906 ( .A(N1144), .B(N1146), .Z(a1stg_sub) );
  GTECH_AND2 C1907 ( .A(N1143), .B(N774), .Z(N1144) );
  GTECH_XOR2 C1908 ( .A(a1stg_opdec[28]), .B(N1142), .Z(N1143) );
  GTECH_XOR2 C1909 ( .A(a1stg_in1_63), .B(a1stg_in2_63), .Z(N1142) );
  GTECH_NOT I_184 ( .A(N1145), .Z(N1146) );
  GTECH_AND2 C1912 ( .A(a1stg_opdec[29]), .B(a1stg_nan_in), .Z(N1145) );
  GTECH_AND2 C1913 ( .A(a2stg_in2_eq_in1_exp), .B(N1147), .Z(a2stg_in2_eq_in1)
         );
  GTECH_NOT I_185 ( .A(a2stg_in2_neq_in1_frac), .Z(N1147) );
  GTECH_OR2 C1915 ( .A(a2stg_in2_gt_in1_exp), .B(N1149), .Z(a2stg_in2_gt_in1)
         );
  GTECH_AND2 C1916 ( .A(N1148), .B(a2stg_in2_gt_in1_frac), .Z(N1149) );
  GTECH_AND2 C1917 ( .A(a2stg_in2_eq_in1_exp), .B(a2stg_in2_neq_in1_frac), .Z(
        N1148) );
  GTECH_AND2 C1918 ( .A(N1151), .B(N1154), .Z(a3stg_sub_in) );
  GTECH_AND2 C1919 ( .A(a2stg_sub), .B(N1150), .Z(N1151) );
  GTECH_NOT I_186 ( .A(a2stg_nan_in), .Z(N1150) );
  GTECH_NOT I_187 ( .A(N1153), .Z(N1154) );
  GTECH_AND2 C1922 ( .A(a2stg_opdec_24_21[0]), .B(N1152), .Z(N1153) );
  GTECH_NOT I_188 ( .A(a2stg_expadd[11]), .Z(N1152) );
  GTECH_AND2 C1925 ( .A(a2stg_sign1), .B(N1150), .Z(N1) );
  GTECH_XOR2 C1926 ( .A(a2stg_sign2), .B(a2stg_opdec_28), .Z(N2) );
  GTECH_NOT I_189 ( .A(N1155), .Z(N3) );
  GTECH_AND2 C1928 ( .A(a2stg_2inf_in), .B(a2stg_sub), .Z(N1155) );
  GTECH_NOT I_190 ( .A(a2stg_in2_eq_in1), .Z(N4) );
  GTECH_OR2 C1930 ( .A(N1179), .B(N1185), .Z(a2stg_faddsub_sign) );
  GTECH_OR2 C1931 ( .A(N1172), .B(N1178), .Z(N1179) );
  GTECH_OR2 C1932 ( .A(N1167), .B(N1171), .Z(N1172) );
  GTECH_OR2 C1933 ( .A(N1162), .B(N1166), .Z(N1167) );
  GTECH_OR2 C1934 ( .A(N1157), .B(N1161), .Z(N1162) );
  GTECH_AND2 C1935 ( .A(N1156), .B(N3), .Z(N1157) );
  GTECH_AND2 C1936 ( .A(N1), .B(N2), .Z(N1156) );
  GTECH_AND2 C1937 ( .A(N1160), .B(N3), .Z(N1161) );
  GTECH_AND2 C1938 ( .A(N1158), .B(N1159), .Z(N1160) );
  GTECH_AND2 C1939 ( .A(N1), .B(N4), .Z(N1158) );
  GTECH_NOT I_191 ( .A(a2stg_in2_gt_in1), .Z(N1159) );
  GTECH_AND2 C1941 ( .A(N1165), .B(N3), .Z(N1166) );
  GTECH_AND2 C1942 ( .A(N1164), .B(N2), .Z(N1165) );
  GTECH_AND2 C1943 ( .A(N1163), .B(N1150), .Z(N1164) );
  GTECH_AND2 C1944 ( .A(N4), .B(a2stg_in2_gt_in1), .Z(N1163) );
  GTECH_AND2 C1945 ( .A(a2stg_sign2), .B(N1170), .Z(N1171) );
  GTECH_OR2 C1946 ( .A(a2stg_snan_in2), .B(N1169), .Z(N1170) );
  GTECH_AND2 C1947 ( .A(a2stg_qnan_in2), .B(N1168), .Z(N1169) );
  GTECH_NOT I_192 ( .A(a2stg_snan_in1), .Z(N1168) );
  GTECH_AND2 C1949 ( .A(a2stg_sign1), .B(N1177), .Z(N1178) );
  GTECH_OR2 C1950 ( .A(N1174), .B(N1176), .Z(N1177) );
  GTECH_AND2 C1951 ( .A(a2stg_snan_in1), .B(N1173), .Z(N1174) );
  GTECH_NOT I_193 ( .A(a2stg_snan_in2), .Z(N1173) );
  GTECH_AND2 C1953 ( .A(a2stg_qnan_in1), .B(N1175), .Z(N1176) );
  GTECH_NOT I_194 ( .A(a2stg_nan_in2), .Z(N1175) );
  GTECH_AND2 C1955 ( .A(N1183), .B(N1184), .Z(N1185) );
  GTECH_AND2 C1956 ( .A(N1182), .B(N1150), .Z(N1183) );
  GTECH_AND2 C1957 ( .A(N1180), .B(N1181), .Z(N1182) );
  GTECH_AND2 C1958 ( .A(N703), .B(a2stg_in2_eq_in1), .Z(N1180) );
  GTECH_XOR2 C1959 ( .A(a2stg_sign1), .B(N2), .Z(N1181) );
  GTECH_NOT I_195 ( .A(a2stg_2inf_in), .Z(N1184) );
  GTECH_OR2 C1961 ( .A(N1186), .B(N1188), .Z(a3stg_sign_in) );
  GTECH_AND2 C1962 ( .A(a2stg_faddsubop), .B(a2stg_faddsub_sign), .Z(N1186) );
  GTECH_AND2 C1963 ( .A(N1187), .B(a2stg_sign2), .Z(N1188) );
  GTECH_NOT I_196 ( .A(a2stg_faddsubop), .Z(N1187) );
  GTECH_AND2 C1965 ( .A(N1198), .B(a2stg_opdec_9_0[9]), .Z(a2stg_cc[1]) );
  GTECH_OR2 C1966 ( .A(N1197), .B(a2stg_nan_in), .Z(N1198) );
  GTECH_OR2 C1967 ( .A(N1191), .B(N1196), .Z(N1197) );
  GTECH_AND2 C1968 ( .A(N1190), .B(a2stg_sub), .Z(N1191) );
  GTECH_AND2 C1969 ( .A(a2stg_sign2), .B(N1189), .Z(N1190) );
  GTECH_NOT I_197 ( .A(a2stg_2zero_in), .Z(N1189) );
  GTECH_AND2 C1971 ( .A(N1193), .B(N1195), .Z(N1196) );
  GTECH_AND2 C1972 ( .A(N4), .B(N1192), .Z(N1193) );
  GTECH_NOT I_198 ( .A(a2stg_sub), .Z(N1192) );
  GTECH_XOR2 C1975 ( .A(a2stg_in2_gt_in1), .B(N1194), .Z(N1195) );
  GTECH_NOT I_199 ( .A(a2stg_sign2), .Z(N1194) );
  GTECH_AND2 C1977 ( .A(N1205), .B(a2stg_opdec_9_0[9]), .Z(a2stg_cc[0]) );
  GTECH_OR2 C1978 ( .A(N1204), .B(a2stg_nan_in), .Z(N1205) );
  GTECH_OR2 C1979 ( .A(N1200), .B(N1203), .Z(N1204) );
  GTECH_AND2 C1980 ( .A(N1199), .B(a2stg_sub), .Z(N1200) );
  GTECH_AND2 C1981 ( .A(N1194), .B(N1189), .Z(N1199) );
  GTECH_AND2 C1984 ( .A(N1201), .B(N1202), .Z(N1203) );
  GTECH_AND2 C1985 ( .A(N4), .B(N1192), .Z(N1201) );
  GTECH_XOR2 C1988 ( .A(a2stg_in2_gt_in1), .B(a2stg_sign2), .Z(N1202) );
  GTECH_OR2 C1989 ( .A(N1206), .B(N1207), .Z(a4stg_sign_in) );
  GTECH_AND2 C1990 ( .A(a3stg_opdec_9_0[8]), .B(a3stg_sign), .Z(N1206) );
  GTECH_AND2 C1991 ( .A(N1026), .B(a4stg_sign2), .Z(N1207) );
  GTECH_AND2 C1993 ( .A(a4stg_fcmpop), .B(a4stg_cc[1]), .Z(add_cc_out_in[1])
         );
  GTECH_AND2 C1994 ( .A(a4stg_fcmpop), .B(a4stg_cc[0]), .Z(add_cc_out_in[0])
         );
  GTECH_OR2 C1995 ( .A(N1217), .B(N1219), .Z(a1stg_nv) );
  GTECH_OR2 C1996 ( .A(N1215), .B(N1216), .Z(N1217) );
  GTECH_OR2 C1997 ( .A(N1213), .B(N1214), .Z(N1215) );
  GTECH_OR2 C1998 ( .A(N1211), .B(N1212), .Z(N1213) );
  GTECH_AND2 C1999 ( .A(a1stg_opdec[29]), .B(N1210), .Z(N1211) );
  GTECH_OR2 C2000 ( .A(N1209), .B(a1stg_snan_in2), .Z(N1210) );
  GTECH_OR2 C2001 ( .A(N1208), .B(a1stg_snan_in1), .Z(N1209) );
  GTECH_AND2 C2002 ( .A(a1stg_2inf_in), .B(a1stg_sub), .Z(N1208) );
  GTECH_AND2 C2003 ( .A(N168), .B(a1stg_snan_in2), .Z(N1212) );
  GTECH_AND2 C2004 ( .A(N775), .B(a1stg_snan_in2), .Z(N1214) );
  GTECH_AND2 C2005 ( .A(a1stg_fcmpesd), .B(a1stg_nan_in), .Z(N1216) );
  GTECH_AND2 C2006 ( .A(a1stg_fcmpsd), .B(N1218), .Z(N1219) );
  GTECH_OR2 C2007 ( .A(a1stg_snan_in1), .B(a1stg_snan_in2), .Z(N1218) );
  GTECH_NOT I_200 ( .A(N1220), .Z(a1stg_of_mask) );
  GTECH_AND2 C2009 ( .A(a1stg_opdec_24_21[3]), .B(a1stg_infnan_in), .Z(N1220)
         );
  GTECH_OR2 C2010 ( .A(N1237), .B(a2stg_nv), .Z(a3stg_nv_in) );
  GTECH_AND2 C2011 ( .A(N1222), .B(N1236), .Z(N1237) );
  GTECH_AND2 C2012 ( .A(N1221), .B(a2stg_opdec_24_21[0]), .Z(N1222) );
  GTECH_NOT I_201 ( .A(a2stg_expadd[11]), .Z(N1221) );
  GTECH_OR2 C2014 ( .A(N1234), .B(N1235), .Z(N1236) );
  GTECH_OR2 C2015 ( .A(N1233), .B(a2stg_frac2hi_neq_0), .Z(N1234) );
  GTECH_OR2 C2016 ( .A(N1194), .B(N1232), .Z(N1233) );
  GTECH_OR2 C2018 ( .A(N1231), .B(a2stg_expadd[0]), .Z(N1232) );
  GTECH_OR2 C2019 ( .A(N1230), .B(a2stg_expadd[1]), .Z(N1231) );
  GTECH_OR2 C2020 ( .A(N1229), .B(a2stg_expadd[2]), .Z(N1230) );
  GTECH_OR2 C2021 ( .A(N1228), .B(a2stg_expadd[3]), .Z(N1229) );
  GTECH_OR2 C2022 ( .A(N1227), .B(a2stg_expadd[4]), .Z(N1228) );
  GTECH_OR2 C2023 ( .A(N1226), .B(a2stg_expadd[5]), .Z(N1227) );
  GTECH_OR2 C2024 ( .A(N1225), .B(a2stg_expadd[6]), .Z(N1226) );
  GTECH_OR2 C2025 ( .A(N1224), .B(a2stg_expadd[7]), .Z(N1225) );
  GTECH_OR2 C2026 ( .A(N1223), .B(a2stg_expadd[8]), .Z(N1224) );
  GTECH_OR2 C2027 ( .A(a2stg_expadd[10]), .B(a2stg_expadd[9]), .Z(N1223) );
  GTECH_AND2 C2028 ( .A(a2stg_opdec[31]), .B(a2stg_frac2lo_neq_0), .Z(N1235)
         );
  GTECH_OR2 C2029 ( .A(N1239), .B(N1243), .Z(a2stg_nx_tmp1) );
  GTECH_AND2 C2030 ( .A(a2stg_opdec_24_21[2]), .B(N1238), .Z(N1239) );
  GTECH_OR2 C2031 ( .A(a2stg_exp[11]), .B(a2stg_exp[10]), .Z(N1238) );
  GTECH_AND2 C2032 ( .A(a2stg_opdec_24_21[1]), .B(N1242), .Z(N1243) );
  GTECH_OR2 C2033 ( .A(N1241), .B(a2stg_exp[7]), .Z(N1242) );
  GTECH_OR2 C2034 ( .A(N1240), .B(a2stg_exp[8]), .Z(N1241) );
  GTECH_OR2 C2035 ( .A(N1238), .B(a2stg_exp[9]), .Z(N1240) );
  GTECH_AND2 C2037 ( .A(N1252), .B(N1264), .Z(a2stg_nx_tmp2) );
  GTECH_OR2 C2038 ( .A(N1246), .B(N1251), .Z(N1252) );
  GTECH_AND2 C2039 ( .A(a2stg_opdec_24_21[2]), .B(N1245), .Z(N1246) );
  GTECH_NOT I_202 ( .A(N1244), .Z(N1245) );
  GTECH_OR2 C2041 ( .A(a2stg_exp[11]), .B(a2stg_exp[10]), .Z(N1244) );
  GTECH_AND2 C2042 ( .A(a2stg_opdec_24_21[1]), .B(N1250), .Z(N1251) );
  GTECH_NOT I_203 ( .A(N1249), .Z(N1250) );
  GTECH_OR2 C2044 ( .A(N1248), .B(a2stg_exp[7]), .Z(N1249) );
  GTECH_OR2 C2045 ( .A(N1247), .B(a2stg_exp[8]), .Z(N1248) );
  GTECH_OR2 C2046 ( .A(N1244), .B(a2stg_exp[9]), .Z(N1247) );
  GTECH_OR2 C2048 ( .A(N1263), .B(a2stg_frac2_63), .Z(N1264) );
  GTECH_OR2 C2049 ( .A(N1262), .B(a2stg_frac2lo_neq_0), .Z(N1263) );
  GTECH_OR2 C2050 ( .A(N1261), .B(a2stg_frac2hi_neq_0), .Z(N1262) );
  GTECH_OR2 C2051 ( .A(N1260), .B(a2stg_exp[1]), .Z(N1261) );
  GTECH_OR2 C2052 ( .A(N1259), .B(a2stg_exp[2]), .Z(N1260) );
  GTECH_OR2 C2053 ( .A(N1258), .B(a2stg_exp[3]), .Z(N1259) );
  GTECH_OR2 C2054 ( .A(N1257), .B(a2stg_exp[4]), .Z(N1258) );
  GTECH_OR2 C2055 ( .A(N1256), .B(a2stg_exp[5]), .Z(N1257) );
  GTECH_OR2 C2056 ( .A(N1255), .B(a2stg_exp[6]), .Z(N1256) );
  GTECH_OR2 C2057 ( .A(N1254), .B(a2stg_exp[7]), .Z(N1255) );
  GTECH_OR2 C2058 ( .A(N1253), .B(a2stg_exp[8]), .Z(N1254) );
  GTECH_OR2 C2059 ( .A(a2stg_exp[10]), .B(a2stg_exp[9]), .Z(N1253) );
  GTECH_AND2 C2060 ( .A(N1268), .B(a2stg_opdec_19_11[5]), .Z(a2stg_nx_tmp3) );
  GTECH_AND2 C2061 ( .A(N1267), .B(a2stg_frac2lo_neq_0), .Z(N1268) );
  GTECH_AND2 C2062 ( .A(N1265), .B(N1266), .Z(N1267) );
  GTECH_AND2 C2063 ( .A(N160), .B(a2stg_sign2), .Z(N1265) );
  GTECH_NOT I_204 ( .A(a2stg_frac2hi_neq_0), .Z(N1266) );
  GTECH_OR2 C2065 ( .A(N1273), .B(a3stg_nx_tmp3), .Z(a3stg_nx) );
  GTECH_AND2 C2066 ( .A(a3stg_a2_expadd_11), .B(N1272), .Z(N1273) );
  GTECH_OR2 C2067 ( .A(N1271), .B(a3stg_nx_tmp2), .Z(N1272) );
  GTECH_AND2 C2068 ( .A(a3stg_nx_tmp1), .B(N1270), .Z(N1271) );
  GTECH_OR2 C2069 ( .A(N1269), .B(a3stg_fsdtoix_nx), .Z(N1270) );
  GTECH_AND2 C2070 ( .A(a3stg_fsdtoi_nx), .B(a3stg_opdec[30]), .Z(N1269) );
  GTECH_AND2 C2071 ( .A(a3stg_opdec[34]), .B(N1274), .Z(N5) );
  GTECH_NOT I_205 ( .A(a3stg_opdec_9_0[7]), .Z(N1274) );
  GTECH_OR2 C2073 ( .A(N1275), .B(N1277), .Z(a4stg_nv_in) );
  GTECH_AND2 C2074 ( .A(N5), .B(a3stg_nv), .Z(N1275) );
  GTECH_AND2 C2075 ( .A(N1276), .B(a4stg_nv2), .Z(N1277) );
  GTECH_NOT I_206 ( .A(N5), .Z(N1276) );
  GTECH_AND2 C2077 ( .A(a3stg_opdec[34]), .B(N1278), .Z(N6) );
  GTECH_NOT I_207 ( .A(a3stg_opdec_9_0[7]), .Z(N1278) );
  GTECH_OR2 C2079 ( .A(N1279), .B(N1281), .Z(a4stg_of_mask_in) );
  GTECH_AND2 C2080 ( .A(N6), .B(a3stg_of_mask), .Z(N1279) );
  GTECH_AND2 C2081 ( .A(N1280), .B(a4stg_of_mask2), .Z(N1281) );
  GTECH_NOT I_208 ( .A(N6), .Z(N1280) );
  GTECH_AND2 C2083 ( .A(a3stg_opdec[34]), .B(N1282), .Z(N7) );
  GTECH_NOT I_209 ( .A(a3stg_opdec_9_0[7]), .Z(N1282) );
  GTECH_OR2 C2085 ( .A(N1283), .B(N1285), .Z(a4stg_nx_in) );
  GTECH_AND2 C2086 ( .A(N7), .B(a3stg_nx), .Z(N1283) );
  GTECH_AND2 C2087 ( .A(N1284), .B(a4stg_nx2), .Z(N1285) );
  GTECH_NOT I_210 ( .A(N7), .Z(N1284) );
  GTECH_OR2 C2089 ( .A(N1298), .B(N1311), .Z(a4stg_in_of) );
  GTECH_AND2 C2090 ( .A(N1297), .B(a4stg_of_mask), .Z(N1298) );
  GTECH_AND2 C2091 ( .A(N1296), .B(a4stg_opdec_7_0[4]), .Z(N1297) );
  GTECH_OR2 C2092 ( .A(a4stg_exp[11]), .B(N1295), .Z(N1296) );
  GTECH_AND2 C2093 ( .A(N1294), .B(a4stg_exp[0]), .Z(N1295) );
  GTECH_AND2 C2094 ( .A(N1293), .B(a4stg_exp[1]), .Z(N1294) );
  GTECH_AND2 C2095 ( .A(N1292), .B(a4stg_exp[2]), .Z(N1293) );
  GTECH_AND2 C2096 ( .A(N1291), .B(a4stg_exp[3]), .Z(N1292) );
  GTECH_AND2 C2097 ( .A(N1290), .B(a4stg_exp[4]), .Z(N1291) );
  GTECH_AND2 C2098 ( .A(N1289), .B(a4stg_exp[5]), .Z(N1290) );
  GTECH_AND2 C2099 ( .A(N1288), .B(a4stg_exp[6]), .Z(N1289) );
  GTECH_AND2 C2100 ( .A(N1287), .B(a4stg_exp[7]), .Z(N1288) );
  GTECH_AND2 C2101 ( .A(N1286), .B(a4stg_exp[8]), .Z(N1287) );
  GTECH_AND2 C2102 ( .A(a4stg_exp[10]), .B(a4stg_exp[9]), .Z(N1286) );
  GTECH_AND2 C2103 ( .A(N1310), .B(a4stg_of_mask), .Z(N1311) );
  GTECH_AND2 C2104 ( .A(N1309), .B(a4stg_opdec_7_0[6]), .Z(N1310) );
  GTECH_OR2 C2105 ( .A(N1301), .B(N1308), .Z(N1309) );
  GTECH_OR2 C2106 ( .A(N1300), .B(a4stg_exp[8]), .Z(N1301) );
  GTECH_OR2 C2107 ( .A(N1299), .B(a4stg_exp[9]), .Z(N1300) );
  GTECH_OR2 C2108 ( .A(a4stg_exp[11]), .B(a4stg_exp[10]), .Z(N1299) );
  GTECH_AND2 C2109 ( .A(N1307), .B(a4stg_exp[0]), .Z(N1308) );
  GTECH_AND2 C2110 ( .A(N1306), .B(a4stg_exp[1]), .Z(N1307) );
  GTECH_AND2 C2111 ( .A(N1305), .B(a4stg_exp[2]), .Z(N1306) );
  GTECH_AND2 C2112 ( .A(N1304), .B(a4stg_exp[3]), .Z(N1305) );
  GTECH_AND2 C2113 ( .A(N1303), .B(a4stg_exp[4]), .Z(N1304) );
  GTECH_AND2 C2114 ( .A(N1302), .B(a4stg_exp[5]), .Z(N1303) );
  GTECH_AND2 C2115 ( .A(a4stg_exp[7]), .B(a4stg_exp[6]), .Z(N1302) );
  GTECH_OR2 C2116 ( .A(N1324), .B(N1335), .Z(add_of_out_tmp1_in) );
  GTECH_AND2 C2117 ( .A(N1323), .B(a4stg_of_mask), .Z(N1324) );
  GTECH_AND2 C2118 ( .A(N1322), .B(a4stg_opdec_7_0[4]), .Z(N1323) );
  GTECH_AND2 C2119 ( .A(N1321), .B(a4stg_round), .Z(N1322) );
  GTECH_AND2 C2120 ( .A(N1320), .B(a4stg_rndup), .Z(N1321) );
  GTECH_AND2 C2121 ( .A(N1319), .B(a4stg_exp[1]), .Z(N1320) );
  GTECH_AND2 C2122 ( .A(N1318), .B(a4stg_exp[2]), .Z(N1319) );
  GTECH_AND2 C2123 ( .A(N1317), .B(a4stg_exp[3]), .Z(N1318) );
  GTECH_AND2 C2124 ( .A(N1316), .B(a4stg_exp[4]), .Z(N1317) );
  GTECH_AND2 C2125 ( .A(N1315), .B(a4stg_exp[5]), .Z(N1316) );
  GTECH_AND2 C2126 ( .A(N1314), .B(a4stg_exp[6]), .Z(N1315) );
  GTECH_AND2 C2127 ( .A(N1313), .B(a4stg_exp[7]), .Z(N1314) );
  GTECH_AND2 C2128 ( .A(N1312), .B(a4stg_exp[8]), .Z(N1313) );
  GTECH_AND2 C2129 ( .A(a4stg_exp[10]), .B(a4stg_exp[9]), .Z(N1312) );
  GTECH_AND2 C2130 ( .A(N1334), .B(a4stg_of_mask), .Z(N1335) );
  GTECH_AND2 C2131 ( .A(N1333), .B(a4stg_opdec_7_0[6]), .Z(N1334) );
  GTECH_AND2 C2132 ( .A(N1331), .B(N1332), .Z(N1333) );
  GTECH_AND2 C2133 ( .A(N1330), .B(a4stg_rndup), .Z(N1331) );
  GTECH_AND2 C2134 ( .A(N1329), .B(a4stg_exp[1]), .Z(N1330) );
  GTECH_AND2 C2135 ( .A(N1328), .B(a4stg_exp[2]), .Z(N1329) );
  GTECH_AND2 C2136 ( .A(N1327), .B(a4stg_exp[3]), .Z(N1328) );
  GTECH_AND2 C2137 ( .A(N1326), .B(a4stg_exp[4]), .Z(N1327) );
  GTECH_AND2 C2138 ( .A(N1325), .B(a4stg_exp[5]), .Z(N1326) );
  GTECH_AND2 C2139 ( .A(a4stg_exp[7]), .B(a4stg_exp[6]), .Z(N1325) );
  GTECH_OR2 C2140 ( .A(a4stg_round), .B(a4stg_opdec_7_0[3]), .Z(N1332) );
  GTECH_OR2 C2141 ( .A(add_of_out_tmp2), .B(N1336), .Z(add_exc_out[3]) );
  GTECH_AND2 C2142 ( .A(add_of_out_tmp1), .B(add_of_out_cout), .Z(N1336) );
  GTECH_OR2 C2143 ( .A(a4stg_round), .B(a4stg_opdec_7_0[3]), .Z(N8) );
  GTECH_OR2 C2144 ( .A(N1350), .B(N1355), .Z(a4stg_uf) );
  GTECH_AND2 C2145 ( .A(N1349), .B(a4stg_faddsub_dtosop), .Z(N1350) );
  GTECH_AND2 C2146 ( .A(N1348), .B(N8), .Z(N1349) );
  GTECH_AND2 C2147 ( .A(N1347), .B(a4stg_frac_neq_0), .Z(N1348) );
  GTECH_NOT I_211 ( .A(N1346), .Z(N1347) );
  GTECH_OR2 C2149 ( .A(N1345), .B(a4stg_exp[0]), .Z(N1346) );
  GTECH_OR2 C2150 ( .A(N1344), .B(a4stg_exp[1]), .Z(N1345) );
  GTECH_OR2 C2151 ( .A(N1343), .B(a4stg_exp[2]), .Z(N1344) );
  GTECH_OR2 C2152 ( .A(N1342), .B(a4stg_exp[3]), .Z(N1343) );
  GTECH_OR2 C2153 ( .A(N1341), .B(a4stg_exp[4]), .Z(N1342) );
  GTECH_OR2 C2154 ( .A(N1340), .B(a4stg_exp[5]), .Z(N1341) );
  GTECH_OR2 C2155 ( .A(N1339), .B(a4stg_exp[6]), .Z(N1340) );
  GTECH_OR2 C2156 ( .A(N1338), .B(a4stg_exp[7]), .Z(N1339) );
  GTECH_OR2 C2157 ( .A(N1337), .B(a4stg_exp[8]), .Z(N1338) );
  GTECH_OR2 C2158 ( .A(a4stg_exp[10]), .B(a4stg_exp[9]), .Z(N1337) );
  GTECH_AND2 C2159 ( .A(N1354), .B(a4stg_shl_data_neq_0), .Z(N1355) );
  GTECH_AND2 C2160 ( .A(N1352), .B(N1353), .Z(N1354) );
  GTECH_AND2 C2161 ( .A(a4stg_opdec[29]), .B(N1351), .Z(N1352) );
  GTECH_NOT I_212 ( .A(N8), .Z(N1351) );
  GTECH_NOT I_213 ( .A(a4stg_denorm_inv), .Z(N1353) );
  GTECH_OR2 C2164 ( .A(N1368), .B(a4stg_nx), .Z(add_nx_out_in) );
  GTECH_OR2 C2165 ( .A(N1361), .B(N1367), .Z(N1368) );
  GTECH_AND2 C2166 ( .A(N1358), .B(N1360), .Z(N1361) );
  GTECH_AND2 C2167 ( .A(N1356), .B(N1357), .Z(N1358) );
  GTECH_AND2 C2168 ( .A(a4stg_of_mask), .B(a4stg_frac_dbl_nx), .Z(N1356) );
  GTECH_OR2 C2169 ( .A(a4stg_opdec_7_0[4]), .B(a5stg_fxtod), .Z(N1357) );
  GTECH_OR2 C2170 ( .A(N1359), .B(a4stg_round), .Z(N1360) );
  GTECH_NOT I_214 ( .A(a4stg_opdec_7_0[4]), .Z(N1359) );
  GTECH_AND2 C2172 ( .A(N1364), .B(N1366), .Z(N1367) );
  GTECH_AND2 C2173 ( .A(N1362), .B(N1363), .Z(N1364) );
  GTECH_AND2 C2174 ( .A(a4stg_of_mask), .B(a4stg_frac_sng_nx), .Z(N1362) );
  GTECH_OR2 C2175 ( .A(a4stg_opdec_7_0[6]), .B(a5stg_fixtos), .Z(N1363) );
  GTECH_OR2 C2176 ( .A(N1365), .B(a4stg_round), .Z(N1366) );
  GTECH_NOT I_215 ( .A(a4stg_opdec_7_0[5]), .Z(N1365) );
  GTECH_OR2 C2178 ( .A(add_nx_out), .B(add_exc_out[3]), .Z(add_exc_out_0) );
  GTECH_OR2 C2179 ( .A(a1stg_snan_in2), .B(N1370), .Z(a2stg_frac1_in_frac1) );
  GTECH_AND2 C2180 ( .A(a1stg_qnan_in2), .B(N1369), .Z(N1370) );
  GTECH_NOT I_216 ( .A(a1stg_snan_in1), .Z(N1369) );
  GTECH_AND2 C2182 ( .A(a1stg_opdec[29]), .B(N1375), .Z(a2stg_frac1_in_frac2)
         );
  GTECH_OR2 C2183 ( .A(N1372), .B(N1374), .Z(N1375) );
  GTECH_OR2 C2184 ( .A(N1371), .B(a1stg_snan_in2), .Z(N1372) );
  GTECH_NOT I_217 ( .A(a1stg_2nan_in), .Z(N1371) );
  GTECH_AND2 C2186 ( .A(a1stg_qnan_in2), .B(N1373), .Z(N1374) );
  GTECH_NOT I_218 ( .A(a1stg_snan_in1), .Z(N1373) );
  GTECH_NOT I_219 ( .A(a1stg_2nan_in), .Z(a1stg_2nan_in_inv) );
  GTECH_NOT I_220 ( .A(a1stg_opdec[29]), .Z(a1stg_faddsubop_inv) );
  GTECH_AND2 C2190 ( .A(N1377), .B(a1stg_opdec[29]), .Z(a2stg_frac1_in_qnan)
         );
  GTECH_OR2 C2191 ( .A(a1stg_nan_in), .B(N1376), .Z(N1377) );
  GTECH_AND2 C2192 ( .A(a1stg_2inf_in), .B(a1stg_sub), .Z(N1376) );
  GTECH_AND2 C2193 ( .A(N1378), .B(a1stg_opdec[29]), .Z(a2stg_frac1_in_nv) );
  GTECH_AND2 C2194 ( .A(a1stg_2inf_in), .B(a1stg_sub), .Z(N1378) );
  GTECH_AND2 C2195 ( .A(N1379), .B(a1stg_faddsubd), .Z(a2stg_frac1_in_nv_dbl)
         );
  GTECH_AND2 C2196 ( .A(a1stg_2inf_in), .B(a1stg_sub), .Z(N1379) );
  GTECH_AND2 C2197 ( .A(a1stg_opdec[29]), .B(N1380), .Z(a2stg_frac2_in_frac1)
         );
  GTECH_NOT I_221 ( .A(a1stg_infnan_in), .Z(N1380) );
  GTECH_AND2 C2199 ( .A(a1stg_snan_in2), .B(N1381), .Z(a2stg_frac2_in_qnan) );
  GTECH_NOT I_222 ( .A(a1stg_opdec[29]), .Z(N1381) );
  GTECH_AND2 C2201 ( .A(a1stg_opdec_24_21[3]), .B(N1382), .Z(
        a1stg_exp_diff_add1) );
  GTECH_NOT I_223 ( .A(a1stg_expadd1[11]), .Z(N1382) );
  GTECH_AND2 C2203 ( .A(a1stg_opdec[29]), .B(a1stg_expadd1[11]), .Z(
        a1stg_exp_diff_add2) );
  GTECH_AND2 C2204 ( .A(N1383), .B(a1stg_fsdtox), .Z(a1stg_exp_diff_5) );
  GTECH_NOT I_224 ( .A(a1stg_expadd2[5]), .Z(N1383) );
  GTECH_OR2 C2206 ( .A(N1384), .B(N1386), .Z(a1stg_exp_diff[10]) );
  GTECH_AND2 C2207 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[10]), .Z(N1384)
         );
  GTECH_AND2 C2208 ( .A(a1stg_exp_diff_add2), .B(N1385), .Z(N1386) );
  GTECH_NOT I_225 ( .A(a1stg_expadd4_inv[10]), .Z(N1385) );
  GTECH_OR2 C2210 ( .A(N1387), .B(N1389), .Z(a1stg_exp_diff[9]) );
  GTECH_AND2 C2211 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[9]), .Z(N1387)
         );
  GTECH_AND2 C2212 ( .A(a1stg_exp_diff_add2), .B(N1388), .Z(N1389) );
  GTECH_NOT I_226 ( .A(a1stg_expadd4_inv[9]), .Z(N1388) );
  GTECH_OR2 C2214 ( .A(N1390), .B(N1392), .Z(a1stg_exp_diff[8]) );
  GTECH_AND2 C2215 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[8]), .Z(N1390)
         );
  GTECH_AND2 C2216 ( .A(a1stg_exp_diff_add2), .B(N1391), .Z(N1392) );
  GTECH_NOT I_227 ( .A(a1stg_expadd4_inv[8]), .Z(N1391) );
  GTECH_OR2 C2218 ( .A(N1393), .B(N1395), .Z(a1stg_exp_diff[7]) );
  GTECH_AND2 C2219 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[7]), .Z(N1393)
         );
  GTECH_AND2 C2220 ( .A(a1stg_exp_diff_add2), .B(N1394), .Z(N1395) );
  GTECH_NOT I_228 ( .A(a1stg_expadd4_inv[7]), .Z(N1394) );
  GTECH_OR2 C2222 ( .A(N1396), .B(N1398), .Z(a1stg_exp_diff[6]) );
  GTECH_AND2 C2223 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[6]), .Z(N1396)
         );
  GTECH_AND2 C2224 ( .A(a1stg_exp_diff_add2), .B(N1397), .Z(N1398) );
  GTECH_NOT I_229 ( .A(a1stg_expadd4_inv[6]), .Z(N1397) );
  GTECH_OR2 C2226 ( .A(N1402), .B(N1403), .Z(a1stg_exp_diff[5]) );
  GTECH_OR2 C2227 ( .A(N1399), .B(N1401), .Z(N1402) );
  GTECH_AND2 C2228 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[5]), .Z(N1399)
         );
  GTECH_AND2 C2229 ( .A(a1stg_exp_diff_add2), .B(N1400), .Z(N1401) );
  GTECH_NOT I_230 ( .A(a1stg_expadd4_inv[5]), .Z(N1400) );
  GTECH_AND2 C2231 ( .A(a1stg_fsdtoix), .B(a1stg_exp_diff_5), .Z(N1403) );
  GTECH_OR2 C2232 ( .A(N1407), .B(N1409), .Z(a1stg_exp_diff[4]) );
  GTECH_OR2 C2233 ( .A(N1404), .B(N1406), .Z(N1407) );
  GTECH_AND2 C2234 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[4]), .Z(N1404)
         );
  GTECH_AND2 C2235 ( .A(a1stg_exp_diff_add2), .B(N1405), .Z(N1406) );
  GTECH_NOT I_231 ( .A(a1stg_expadd4_inv[4]), .Z(N1405) );
  GTECH_AND2 C2237 ( .A(a1stg_fsdtoix), .B(N1408), .Z(N1409) );
  GTECH_NOT I_232 ( .A(a1stg_expadd2[4]), .Z(N1408) );
  GTECH_OR2 C2239 ( .A(N1413), .B(N1415), .Z(a1stg_exp_diff[3]) );
  GTECH_OR2 C2240 ( .A(N1410), .B(N1412), .Z(N1413) );
  GTECH_AND2 C2241 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[3]), .Z(N1410)
         );
  GTECH_AND2 C2242 ( .A(a1stg_exp_diff_add2), .B(N1411), .Z(N1412) );
  GTECH_NOT I_233 ( .A(a1stg_expadd4_inv[3]), .Z(N1411) );
  GTECH_AND2 C2244 ( .A(a1stg_fsdtoix), .B(N1414), .Z(N1415) );
  GTECH_NOT I_234 ( .A(a1stg_expadd2[3]), .Z(N1414) );
  GTECH_OR2 C2246 ( .A(N1419), .B(N1421), .Z(a1stg_exp_diff[2]) );
  GTECH_OR2 C2247 ( .A(N1416), .B(N1418), .Z(N1419) );
  GTECH_AND2 C2248 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[2]), .Z(N1416)
         );
  GTECH_AND2 C2249 ( .A(a1stg_exp_diff_add2), .B(N1417), .Z(N1418) );
  GTECH_NOT I_235 ( .A(a1stg_expadd4_inv[2]), .Z(N1417) );
  GTECH_AND2 C2251 ( .A(a1stg_fsdtoix), .B(N1420), .Z(N1421) );
  GTECH_NOT I_236 ( .A(a1stg_expadd2[2]), .Z(N1420) );
  GTECH_OR2 C2253 ( .A(N1425), .B(N1427), .Z(a1stg_exp_diff[1]) );
  GTECH_OR2 C2254 ( .A(N1422), .B(N1424), .Z(N1425) );
  GTECH_AND2 C2255 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[1]), .Z(N1422)
         );
  GTECH_AND2 C2256 ( .A(a1stg_exp_diff_add2), .B(N1423), .Z(N1424) );
  GTECH_NOT I_237 ( .A(a1stg_expadd4_inv[1]), .Z(N1423) );
  GTECH_AND2 C2258 ( .A(a1stg_fsdtoix), .B(N1426), .Z(N1427) );
  GTECH_NOT I_238 ( .A(a1stg_expadd2[1]), .Z(N1426) );
  GTECH_OR2 C2260 ( .A(N1431), .B(N1433), .Z(a1stg_exp_diff[0]) );
  GTECH_OR2 C2261 ( .A(N1428), .B(N1430), .Z(N1431) );
  GTECH_AND2 C2262 ( .A(a1stg_exp_diff_add1), .B(a1stg_expadd1[0]), .Z(N1428)
         );
  GTECH_AND2 C2263 ( .A(a1stg_exp_diff_add2), .B(N1429), .Z(N1430) );
  GTECH_NOT I_239 ( .A(a1stg_expadd4_inv[0]), .Z(N1429) );
  GTECH_AND2 C2265 ( .A(a1stg_fsdtoix), .B(N1432), .Z(N1433) );
  GTECH_NOT I_240 ( .A(a1stg_expadd2[0]), .Z(N1432) );
  GTECH_OR2 C2267 ( .A(a1stg_exp_diff[5]), .B(N1437), .Z(a2stg_shr_cnt_in[5])
         );
  GTECH_OR2 C2268 ( .A(N1436), .B(a1stg_exp_diff[6]), .Z(N1437) );
  GTECH_OR2 C2269 ( .A(N1435), .B(a1stg_exp_diff[7]), .Z(N1436) );
  GTECH_OR2 C2270 ( .A(N1434), .B(a1stg_exp_diff[8]), .Z(N1435) );
  GTECH_OR2 C2271 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1434)
         );
  GTECH_OR2 C2272 ( .A(a1stg_exp_diff[4]), .B(N1441), .Z(a2stg_shr_cnt_in[4])
         );
  GTECH_OR2 C2273 ( .A(N1440), .B(a1stg_exp_diff[6]), .Z(N1441) );
  GTECH_OR2 C2274 ( .A(N1439), .B(a1stg_exp_diff[7]), .Z(N1440) );
  GTECH_OR2 C2275 ( .A(N1438), .B(a1stg_exp_diff[8]), .Z(N1439) );
  GTECH_OR2 C2276 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1438)
         );
  GTECH_OR2 C2277 ( .A(a1stg_exp_diff[3]), .B(N1445), .Z(a2stg_shr_cnt_in[3])
         );
  GTECH_OR2 C2278 ( .A(N1444), .B(a1stg_exp_diff[6]), .Z(N1445) );
  GTECH_OR2 C2279 ( .A(N1443), .B(a1stg_exp_diff[7]), .Z(N1444) );
  GTECH_OR2 C2280 ( .A(N1442), .B(a1stg_exp_diff[8]), .Z(N1443) );
  GTECH_OR2 C2281 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1442)
         );
  GTECH_OR2 C2282 ( .A(a1stg_exp_diff[2]), .B(N1449), .Z(a2stg_shr_cnt_in[2])
         );
  GTECH_OR2 C2283 ( .A(N1448), .B(a1stg_exp_diff[6]), .Z(N1449) );
  GTECH_OR2 C2284 ( .A(N1447), .B(a1stg_exp_diff[7]), .Z(N1448) );
  GTECH_OR2 C2285 ( .A(N1446), .B(a1stg_exp_diff[8]), .Z(N1447) );
  GTECH_OR2 C2286 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1446)
         );
  GTECH_OR2 C2287 ( .A(a1stg_exp_diff[1]), .B(N1453), .Z(a2stg_shr_cnt_in[1])
         );
  GTECH_OR2 C2288 ( .A(N1452), .B(a1stg_exp_diff[6]), .Z(N1453) );
  GTECH_OR2 C2289 ( .A(N1451), .B(a1stg_exp_diff[7]), .Z(N1452) );
  GTECH_OR2 C2290 ( .A(N1450), .B(a1stg_exp_diff[8]), .Z(N1451) );
  GTECH_OR2 C2291 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1450)
         );
  GTECH_OR2 C2292 ( .A(a1stg_exp_diff[0]), .B(N1457), .Z(a2stg_shr_cnt_in[0])
         );
  GTECH_OR2 C2293 ( .A(N1456), .B(a1stg_exp_diff[6]), .Z(N1457) );
  GTECH_OR2 C2294 ( .A(N1455), .B(a1stg_exp_diff[7]), .Z(N1456) );
  GTECH_OR2 C2295 ( .A(N1454), .B(a1stg_exp_diff[8]), .Z(N1455) );
  GTECH_OR2 C2296 ( .A(a1stg_exp_diff[10]), .B(a1stg_exp_diff[9]), .Z(N1454)
         );
  GTECH_NOT I_241 ( .A(a2stg_shr_cnt_in[5]), .Z(a2stg_shr_cnt_5_inv_in) );
  GTECH_AND2 C2298 ( .A(a2stg_opdec_24_21[3]), .B(a6stg_step), .Z(
        a2stg_shr_frac2_shr_int) );
  GTECH_AND2 C2299 ( .A(N1464), .B(a6stg_step), .Z(a2stg_shr_frac2_shr_dbl) );
  GTECH_OR2 C2300 ( .A(N1459), .B(N1463), .Z(N1464) );
  GTECH_AND2 C2301 ( .A(a2stg_opdec_19_11[4]), .B(N1458), .Z(N1459) );
  GTECH_OR2 C2302 ( .A(a2stg_exp[11]), .B(a2stg_exp[10]), .Z(N1458) );
  GTECH_AND2 C2303 ( .A(a2stg_opdec_19_11[6]), .B(N1462), .Z(N1463) );
  GTECH_OR2 C2304 ( .A(N1461), .B(a2stg_exp[7]), .Z(N1462) );
  GTECH_OR2 C2305 ( .A(N1460), .B(a2stg_exp[8]), .Z(N1461) );
  GTECH_OR2 C2306 ( .A(N1458), .B(a2stg_exp[9]), .Z(N1460) );
  GTECH_AND2 C2308 ( .A(N1471), .B(a6stg_step), .Z(a2stg_shr_frac2_shr_sng) );
  GTECH_OR2 C2309 ( .A(N1466), .B(N1470), .Z(N1471) );
  GTECH_AND2 C2310 ( .A(a2stg_opdec_19_11[5]), .B(N1465), .Z(N1466) );
  GTECH_OR2 C2311 ( .A(a2stg_exp[11]), .B(a2stg_exp[10]), .Z(N1465) );
  GTECH_AND2 C2312 ( .A(a2stg_opdec_19_11[7]), .B(N1469), .Z(N1470) );
  GTECH_OR2 C2313 ( .A(N1468), .B(a2stg_exp[7]), .Z(N1469) );
  GTECH_OR2 C2314 ( .A(N1467), .B(a2stg_exp[8]), .Z(N1468) );
  GTECH_OR2 C2315 ( .A(N1465), .B(a2stg_exp[9]), .Z(N1467) );
  GTECH_AND2 C2317 ( .A(a2stg_opdec_24_21[0]), .B(a6stg_step), .Z(
        a2stg_shr_frac2_max) );
  GTECH_AND2 C2318 ( .A(a2stg_sub), .B(a6stg_step), .Z(a2stg_sub_step) );
  GTECH_OR2 C2319 ( .A(N1491), .B(N1494), .Z(a1stg_faddsub_clamp63_0) );
  GTECH_OR2 C2320 ( .A(N1487), .B(N1490), .Z(N1491) );
  GTECH_OR2 C2321 ( .A(N1483), .B(N1486), .Z(N1487) );
  GTECH_OR2 C2322 ( .A(N1479), .B(N1482), .Z(N1483) );
  GTECH_OR2 C2323 ( .A(N1475), .B(N1478), .Z(N1479) );
  GTECH_OR2 C2324 ( .A(N1472), .B(N1474), .Z(N1475) );
  GTECH_AND2 C2325 ( .A(a1stg_expadd1[11]), .B(N1385), .Z(N1472) );
  GTECH_AND2 C2327 ( .A(N1473), .B(a1stg_expadd1[10]), .Z(N1474) );
  GTECH_NOT I_242 ( .A(a1stg_expadd1[11]), .Z(N1473) );
  GTECH_OR2 C2329 ( .A(N1476), .B(N1477), .Z(N1478) );
  GTECH_AND2 C2330 ( .A(a1stg_expadd1[11]), .B(N1388), .Z(N1476) );
  GTECH_AND2 C2332 ( .A(N1473), .B(a1stg_expadd1[9]), .Z(N1477) );
  GTECH_OR2 C2334 ( .A(N1480), .B(N1481), .Z(N1482) );
  GTECH_AND2 C2335 ( .A(a1stg_expadd1[11]), .B(N1391), .Z(N1480) );
  GTECH_AND2 C2337 ( .A(N1473), .B(a1stg_expadd1[8]), .Z(N1481) );
  GTECH_OR2 C2339 ( .A(N1484), .B(N1485), .Z(N1486) );
  GTECH_AND2 C2340 ( .A(a1stg_expadd1[11]), .B(N1394), .Z(N1484) );
  GTECH_AND2 C2342 ( .A(N1473), .B(a1stg_expadd1[7]), .Z(N1485) );
  GTECH_OR2 C2344 ( .A(N1488), .B(N1489), .Z(N1490) );
  GTECH_AND2 C2345 ( .A(a1stg_expadd1[11]), .B(N1397), .Z(N1488) );
  GTECH_AND2 C2347 ( .A(N1473), .B(a1stg_expadd1[6]), .Z(N1489) );
  GTECH_OR2 C2349 ( .A(N1492), .B(N1493), .Z(N1494) );
  GTECH_AND2 C2350 ( .A(a1stg_expadd1[11]), .B(N1429), .Z(N1492) );
  GTECH_AND2 C2352 ( .A(N1473), .B(a1stg_expadd1[0]), .Z(N1493) );
  GTECH_OR2 C2354 ( .A(N1495), .B(N1498), .Z(a2stg_fracadd_frac2_inv_in) );
  GTECH_AND2 C2355 ( .A(a1stg_fixtosd), .B(a1stg_in2_63), .Z(N1495) );
  GTECH_AND2 C2356 ( .A(N1496), .B(N1497), .Z(N1498) );
  GTECH_AND2 C2357 ( .A(a1stg_opdec[29]), .B(a1stg_sub), .Z(N1496) );
  GTECH_NOT I_243 ( .A(a1stg_faddsub_clamp63_0), .Z(N1497) );
  GTECH_AND2 C2359 ( .A(N1499), .B(a1stg_faddsub_clamp63_0), .Z(
        a2stg_fracadd_frac2_inv_shr1_in) );
  GTECH_AND2 C2360 ( .A(a1stg_opdec[29]), .B(a1stg_sub), .Z(N1499) );
  GTECH_OR2 C2361 ( .A(N1502), .B(N1504), .Z(a2stg_fracadd_frac2_in) );
  GTECH_OR2 C2362 ( .A(N1501), .B(N168), .Z(N1502) );
  GTECH_AND2 C2363 ( .A(a1stg_fixtosd), .B(N1500), .Z(N1501) );
  GTECH_NOT I_244 ( .A(a1stg_in2_63), .Z(N1500) );
  GTECH_AND2 C2365 ( .A(a1stg_opdec[29]), .B(N1503), .Z(N1504) );
  GTECH_NOT I_245 ( .A(a1stg_sub), .Z(N1503) );
  GTECH_OR2 C2367 ( .A(N1505), .B(N1506), .Z(a2stg_fracadd_cin_in) );
  GTECH_AND2 C2368 ( .A(a1stg_fixtosd), .B(a1stg_in2_63), .Z(N1505) );
  GTECH_AND2 C2369 ( .A(a1stg_opdec[29]), .B(a1stg_sub), .Z(N1506) );
  GTECH_AND2 C2370 ( .A(a2stg_opdec_19_11[8]), .B(N1513), .Z(a3stg_exp_7ff) );
  GTECH_AND2 C2371 ( .A(N1512), .B(a2stg_exp[0]), .Z(N1513) );
  GTECH_AND2 C2372 ( .A(N1511), .B(a2stg_exp[1]), .Z(N1512) );
  GTECH_AND2 C2373 ( .A(N1510), .B(a2stg_exp[2]), .Z(N1511) );
  GTECH_AND2 C2374 ( .A(N1509), .B(a2stg_exp[3]), .Z(N1510) );
  GTECH_AND2 C2375 ( .A(N1508), .B(a2stg_exp[4]), .Z(N1509) );
  GTECH_AND2 C2376 ( .A(N1507), .B(a2stg_exp[5]), .Z(N1508) );
  GTECH_AND2 C2377 ( .A(a2stg_exp[7]), .B(a2stg_exp[6]), .Z(N1507) );
  GTECH_AND2 C2378 ( .A(a2stg_opdec_9_0[3]), .B(N1523), .Z(a3stg_exp_ff) );
  GTECH_AND2 C2379 ( .A(N1522), .B(a2stg_exp[0]), .Z(N1523) );
  GTECH_AND2 C2380 ( .A(N1521), .B(a2stg_exp[1]), .Z(N1522) );
  GTECH_AND2 C2381 ( .A(N1520), .B(a2stg_exp[2]), .Z(N1521) );
  GTECH_AND2 C2382 ( .A(N1519), .B(a2stg_exp[3]), .Z(N1520) );
  GTECH_AND2 C2383 ( .A(N1518), .B(a2stg_exp[4]), .Z(N1519) );
  GTECH_AND2 C2384 ( .A(N1517), .B(a2stg_exp[5]), .Z(N1518) );
  GTECH_AND2 C2385 ( .A(N1516), .B(a2stg_exp[6]), .Z(N1517) );
  GTECH_AND2 C2386 ( .A(N1515), .B(a2stg_exp[7]), .Z(N1516) );
  GTECH_AND2 C2387 ( .A(N1514), .B(a2stg_exp[8]), .Z(N1515) );
  GTECH_AND2 C2388 ( .A(a2stg_exp[10]), .B(a2stg_exp[9]), .Z(N1514) );
  GTECH_OR2 C2389 ( .A(N1532), .B(N1544), .Z(a3stg_exp_add) );
  GTECH_AND2 C2390 ( .A(a2stg_opdec_19_11[8]), .B(N1531), .Z(N1532) );
  GTECH_NOT I_246 ( .A(N1530), .Z(N1531) );
  GTECH_AND2 C2392 ( .A(N1529), .B(a2stg_exp[0]), .Z(N1530) );
  GTECH_AND2 C2393 ( .A(N1528), .B(a2stg_exp[1]), .Z(N1529) );
  GTECH_AND2 C2394 ( .A(N1527), .B(a2stg_exp[2]), .Z(N1528) );
  GTECH_AND2 C2395 ( .A(N1526), .B(a2stg_exp[3]), .Z(N1527) );
  GTECH_AND2 C2396 ( .A(N1525), .B(a2stg_exp[4]), .Z(N1526) );
  GTECH_AND2 C2397 ( .A(N1524), .B(a2stg_exp[5]), .Z(N1525) );
  GTECH_AND2 C2398 ( .A(a2stg_exp[7]), .B(a2stg_exp[6]), .Z(N1524) );
  GTECH_AND2 C2399 ( .A(a2stg_opdec_9_0[3]), .B(N1543), .Z(N1544) );
  GTECH_NOT I_247 ( .A(N1542), .Z(N1543) );
  GTECH_AND2 C2401 ( .A(N1541), .B(a2stg_exp[0]), .Z(N1542) );
  GTECH_AND2 C2402 ( .A(N1540), .B(a2stg_exp[1]), .Z(N1541) );
  GTECH_AND2 C2403 ( .A(N1539), .B(a2stg_exp[2]), .Z(N1540) );
  GTECH_AND2 C2404 ( .A(N1538), .B(a2stg_exp[3]), .Z(N1539) );
  GTECH_AND2 C2405 ( .A(N1537), .B(a2stg_exp[4]), .Z(N1538) );
  GTECH_AND2 C2406 ( .A(N1536), .B(a2stg_exp[5]), .Z(N1537) );
  GTECH_AND2 C2407 ( .A(N1535), .B(a2stg_exp[6]), .Z(N1536) );
  GTECH_AND2 C2408 ( .A(N1534), .B(a2stg_exp[7]), .Z(N1535) );
  GTECH_AND2 C2409 ( .A(N1533), .B(a2stg_exp[8]), .Z(N1534) );
  GTECH_AND2 C2410 ( .A(a2stg_exp[10]), .B(a2stg_exp[9]), .Z(N1533) );
  GTECH_AND2 C2411 ( .A(a2stg_faddsubop), .B(N9), .Z(a2stg_expdec_neq_0) );
  GTECH_NOT I_248 ( .A(a3stg_opdec_9_0[3]), .Z(a3stg_fdtos_inv) );
  GTECH_NOT I_249 ( .A(a4stg_opdec_7_0[7]), .Z(a4stg_fixtos_fxtod_inv) );
  GTECH_NOT I_250 ( .A(N1546), .Z(a4stg_rnd_frac_add_inv) );
  GTECH_OR2 C2415 ( .A(a3stg_fsdtoix), .B(N1545), .Z(N1546) );
  GTECH_AND2 C2416 ( .A(a3stg_faddsubop), .B(N53), .Z(N1545) );
  GTECH_OR2 C2417 ( .A(N1547), .B(N1548), .Z(a4stg_shl_cnt_in[9]) );
  GTECH_AND2 C2418 ( .A(a3stg_denorm), .B(N54), .Z(N1547) );
  GTECH_AND2 C2419 ( .A(a3stg_denorm_inv), .B(N55), .Z(N1548) );
  GTECH_OR2 C2420 ( .A(N1549), .B(N1550), .Z(a4stg_shl_cnt_in[8]) );
  GTECH_AND2 C2421 ( .A(a3stg_denorm), .B(N58), .Z(N1549) );
  GTECH_AND2 C2422 ( .A(a3stg_denorm_inv), .B(N61), .Z(N1550) );
  GTECH_OR2 C2423 ( .A(N1551), .B(N1552), .Z(a4stg_shl_cnt_in[7]) );
  GTECH_AND2 C2424 ( .A(a3stg_denorm), .B(N64), .Z(N1551) );
  GTECH_AND2 C2425 ( .A(a3stg_denorm_inv), .B(N67), .Z(N1552) );
  GTECH_OR2 C2426 ( .A(N1553), .B(N1554), .Z(a4stg_shl_cnt_in[6]) );
  GTECH_AND2 C2427 ( .A(a3stg_denorm), .B(N69), .Z(N1553) );
  GTECH_AND2 C2428 ( .A(a3stg_denorm_inv), .B(N71), .Z(N1554) );
  GTECH_OR2 C2429 ( .A(N1555), .B(N1556), .Z(a4stg_shl_cnt_in[5]) );
  GTECH_AND2 C2430 ( .A(a3stg_denorm), .B(a3stg_exp[5]), .Z(N1555) );
  GTECH_AND2 C2431 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[5]), .Z(N1556) );
  GTECH_OR2 C2432 ( .A(N1557), .B(N1558), .Z(a4stg_shl_cnt_in[4]) );
  GTECH_AND2 C2433 ( .A(a3stg_denorm), .B(a3stg_exp[4]), .Z(N1557) );
  GTECH_AND2 C2434 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[4]), .Z(N1558) );
  GTECH_OR2 C2435 ( .A(N1559), .B(N1560), .Z(a4stg_shl_cnt_in[3]) );
  GTECH_AND2 C2436 ( .A(a3stg_denorm), .B(a3stg_exp[3]), .Z(N1559) );
  GTECH_AND2 C2437 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[3]), .Z(N1560) );
  GTECH_OR2 C2438 ( .A(N1561), .B(N1562), .Z(a4stg_shl_cnt_in[2]) );
  GTECH_AND2 C2439 ( .A(a3stg_denorm), .B(a3stg_exp[2]), .Z(N1561) );
  GTECH_AND2 C2440 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[2]), .Z(N1562) );
  GTECH_OR2 C2441 ( .A(N1563), .B(N1564), .Z(a4stg_shl_cnt_in[1]) );
  GTECH_AND2 C2442 ( .A(a3stg_denorm), .B(a3stg_exp[1]), .Z(N1563) );
  GTECH_AND2 C2443 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[1]), .Z(N1564) );
  GTECH_OR2 C2444 ( .A(N1565), .B(N1566), .Z(a4stg_shl_cnt_in[0]) );
  GTECH_AND2 C2445 ( .A(a3stg_denorm), .B(a3stg_exp[0]), .Z(N1565) );
  GTECH_AND2 C2446 ( .A(a3stg_denorm_inv), .B(a3stg_lead0[0]), .Z(N1566) );
  GTECH_OR2 C2447 ( .A(a5stg_fixtos), .B(a4stg_opdec_7_0[6]), .Z(a4stg_rnd_sng) );
  GTECH_OR2 C2448 ( .A(a5stg_fxtod), .B(a4stg_opdec_7_0[4]), .Z(a4stg_rnd_dbl)
         );
  GTECH_OR2 C2449 ( .A(N1572), .B(N1575), .Z(a4stg_rndup_sng) );
  GTECH_OR2 C2450 ( .A(N1569), .B(N1571), .Z(N1572) );
  GTECH_AND2 C2451 ( .A(N1568), .B(a4stg_frac_sng_nx), .Z(N1569) );
  GTECH_AND2 C2452 ( .A(N830), .B(N1567), .Z(N1568) );
  GTECH_NOT I_251 ( .A(a4stg_sign), .Z(N1567) );
  GTECH_AND2 C2454 ( .A(N1570), .B(a4stg_frac_sng_nx), .Z(N1571) );
  GTECH_AND2 C2455 ( .A(N831), .B(a4stg_sign), .Z(N1570) );
  GTECH_AND2 C2456 ( .A(N1573), .B(N1574), .Z(N1575) );
  GTECH_AND2 C2457 ( .A(N833), .B(a4stg_rnd_frac_39), .Z(N1573) );
  GTECH_OR2 C2458 ( .A(a4stg_frac_38_0_nx), .B(a4stg_rnd_frac_40), .Z(N1574)
         );
  GTECH_OR2 C2459 ( .A(N1581), .B(N1584), .Z(a4stg_rndup_dbl) );
  GTECH_OR2 C2460 ( .A(N1578), .B(N1580), .Z(N1581) );
  GTECH_AND2 C2461 ( .A(N1577), .B(a4stg_frac_dbl_nx), .Z(N1578) );
  GTECH_AND2 C2462 ( .A(N825), .B(N1576), .Z(N1577) );
  GTECH_NOT I_252 ( .A(a4stg_sign), .Z(N1576) );
  GTECH_AND2 C2464 ( .A(N1579), .B(a4stg_frac_dbl_nx), .Z(N1580) );
  GTECH_AND2 C2465 ( .A(N826), .B(a4stg_sign), .Z(N1579) );
  GTECH_AND2 C2466 ( .A(N1582), .B(N1583), .Z(N1584) );
  GTECH_AND2 C2467 ( .A(N828), .B(a4stg_rnd_frac_10), .Z(N1582) );
  GTECH_OR2 C2468 ( .A(a4stg_frac_9_0_nx), .B(a4stg_rnd_frac_11), .Z(N1583) );
  GTECH_OR2 C2469 ( .A(N1587), .B(N1589), .Z(a4stg_rndup) );
  GTECH_OR2 C2470 ( .A(N1585), .B(N1586), .Z(N1587) );
  GTECH_AND2 C2471 ( .A(a4stg_opdec_7_0[4]), .B(a4stg_rndup_dbl), .Z(N1585) );
  GTECH_AND2 C2472 ( .A(a4stg_opdec_7_0[5]), .B(a4stg_rndup_sng), .Z(N1586) );
  GTECH_AND2 C2473 ( .A(N1588), .B(a4stg_of_mask), .Z(N1589) );
  GTECH_AND2 C2474 ( .A(a4stg_opdec_7_0[3]), .B(a4stg_rndup_sng), .Z(N1588) );
  GTECH_OR2 C2475 ( .A(N1590), .B(N1591), .Z(a5stg_rndup) );
  GTECH_AND2 C2476 ( .A(a5stg_fxtod), .B(a4stg_rndup_dbl), .Z(N1590) );
  GTECH_AND2 C2477 ( .A(a5stg_fixtos), .B(a4stg_rndup_sng), .Z(N1591) );
  GTECH_NOT I_253 ( .A(a4stg_in_of), .Z(N10) );
  GTECH_OR2 C2479 ( .A(N1597), .B(N1598), .Z(add_frac_out_rndadd) );
  GTECH_OR2 C2480 ( .A(N1594), .B(N1596), .Z(N1597) );
  GTECH_AND2 C2481 ( .A(N1593), .B(N10), .Z(N1594) );
  GTECH_AND2 C2482 ( .A(N1592), .B(a4stg_rndup), .Z(N1593) );
  GTECH_AND2 C2483 ( .A(a4stg_opdec[29]), .B(a4stg_round), .Z(N1592) );
  GTECH_AND2 C2484 ( .A(N1595), .B(N10), .Z(N1596) );
  GTECH_AND2 C2485 ( .A(a4stg_opdec_7_0[3]), .B(a4stg_rndup), .Z(N1595) );
  GTECH_AND2 C2486 ( .A(a5stg_fixtos_fxtod), .B(a5stg_rndup), .Z(N1598) );
  GTECH_NOT I_254 ( .A(a4stg_rndup), .Z(N11) );
  GTECH_NOT I_255 ( .A(a4stg_in_of), .Z(N12) );
  GTECH_OR2 C2489 ( .A(N1607), .B(a4stg_fsdtoix), .Z(add_frac_out_rnd_frac) );
  GTECH_OR2 C2490 ( .A(N1604), .B(N1606), .Z(N1607) );
  GTECH_OR2 C2491 ( .A(N1601), .B(N1603), .Z(N1604) );
  GTECH_AND2 C2492 ( .A(N1600), .B(N12), .Z(N1601) );
  GTECH_AND2 C2493 ( .A(N1599), .B(N11), .Z(N1600) );
  GTECH_AND2 C2494 ( .A(a4stg_opdec[29]), .B(a4stg_round), .Z(N1599) );
  GTECH_AND2 C2495 ( .A(N1602), .B(N12), .Z(N1603) );
  GTECH_AND2 C2496 ( .A(a4stg_opdec_7_0[3]), .B(N11), .Z(N1602) );
  GTECH_AND2 C2497 ( .A(a5stg_fixtos_fxtod), .B(N1605), .Z(N1606) );
  GTECH_NOT I_256 ( .A(a5stg_rndup), .Z(N1605) );
  GTECH_OR2 C2499 ( .A(N1611), .B(a4stg_opdec_7_0[2]), .Z(add_frac_out_shl) );
  GTECH_AND2 C2500 ( .A(N1609), .B(N1610), .Z(N1611) );
  GTECH_AND2 C2501 ( .A(a4stg_opdec[29]), .B(N1608), .Z(N1609) );
  GTECH_NOT I_257 ( .A(a4stg_round), .Z(N1608) );
  GTECH_NOT I_258 ( .A(a4stg_in_of), .Z(N1610) );
  GTECH_NOT I_259 ( .A(N1616), .Z(a4stg_to_0) );
  GTECH_OR2 C2505 ( .A(N1614), .B(N1615), .Z(N1616) );
  GTECH_OR2 C2506 ( .A(N170), .B(N1613), .Z(N1614) );
  GTECH_AND2 C2507 ( .A(N173), .B(N1612), .Z(N1613) );
  GTECH_NOT I_260 ( .A(a4stg_sign), .Z(N1612) );
  GTECH_AND2 C2509 ( .A(N174), .B(a4stg_sign), .Z(N1615) );
  GTECH_NOT I_261 ( .A(a4stg_in_of), .Z(N13) );
  GTECH_OR2 C2511 ( .A(N1622), .B(N1623), .Z(add_exp_out_expinc) );
  GTECH_OR2 C2512 ( .A(N1619), .B(N1621), .Z(N1622) );
  GTECH_AND2 C2513 ( .A(N1618), .B(N13), .Z(N1619) );
  GTECH_AND2 C2514 ( .A(N1617), .B(a4stg_rndup), .Z(N1618) );
  GTECH_AND2 C2515 ( .A(a4stg_opdec[29]), .B(a4stg_round), .Z(N1617) );
  GTECH_AND2 C2516 ( .A(N1620), .B(N13), .Z(N1621) );
  GTECH_AND2 C2517 ( .A(a4stg_opdec_7_0[3]), .B(a4stg_rndup), .Z(N1620) );
  GTECH_AND2 C2518 ( .A(a5stg_fixtos_fxtod), .B(a5stg_rndup), .Z(N1623) );
  GTECH_NOT I_262 ( .A(a4stg_in_of), .Z(N14) );
  GTECH_OR2 C2520 ( .A(N1627), .B(a5stg_fixtos_fxtod), .Z(add_exp_out_exp) );
  GTECH_OR2 C2521 ( .A(N1625), .B(N1626), .Z(N1627) );
  GTECH_AND2 C2522 ( .A(N1624), .B(N14), .Z(N1625) );
  GTECH_AND2 C2523 ( .A(a4stg_opdec[29]), .B(a4stg_round), .Z(N1624) );
  GTECH_AND2 C2524 ( .A(a4stg_opdec_7_0[3]), .B(N14), .Z(N1626) );
  GTECH_NOT I_263 ( .A(a4stg_in_of), .Z(N15) );
  GTECH_OR2 C2527 ( .A(N1633), .B(N1634), .Z(add_exp_out_exp1) );
  GTECH_OR2 C2528 ( .A(N1630), .B(N1632), .Z(N1633) );
  GTECH_AND2 C2529 ( .A(N1629), .B(N15), .Z(N1630) );
  GTECH_AND2 C2530 ( .A(N1628), .B(N11), .Z(N1629) );
  GTECH_AND2 C2531 ( .A(a4stg_opdec[29]), .B(a4stg_round), .Z(N1628) );
  GTECH_AND2 C2532 ( .A(N1631), .B(N15), .Z(N1632) );
  GTECH_AND2 C2533 ( .A(a4stg_opdec_7_0[3]), .B(N11), .Z(N1631) );
  GTECH_AND2 C2534 ( .A(a5stg_fixtos_fxtod), .B(N1605), .Z(N1634) );
  GTECH_OR2 C2536 ( .A(N1637), .B(a4stg_opdec_7_0[2]), .Z(add_exp_out_expadd)
         );
  GTECH_AND2 C2537 ( .A(N1635), .B(N1636), .Z(N1637) );
  GTECH_AND2 C2538 ( .A(a4stg_opdec[29]), .B(N1608), .Z(N1635) );
  GTECH_NOT I_264 ( .A(a4stg_in_of), .Z(N1636) );
  GTECH_NOT I_265 ( .A(a4stg_to_0), .Z(a4stg_to_0_inv) );
endmodule


module dffe_SIZE11 ( din, en, clk, q, se, si, so );
  input [10:0] din;
  output [10:0] q;
  input [10:0] si;
  output [10:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16;
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N16) );
  SELECT_OP C59 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C67 ( .A(N3), .B(N2), .Z(N15) );
  GTECH_NOT I_2 ( .A(N15), .Z(N16) );
endmodule


module dffe_SIZE13 ( din, en, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18;
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N18) );
  SELECT_OP C67 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C75 ( .A(N3), .B(N2), .Z(N17) );
  GTECH_NOT I_2 ( .A(N17), .Z(N18) );
endmodule


module dffe_SIZE12 ( din, en, clk, q, se, si, so );
  input [11:0] din;
  output [11:0] q;
  input [11:0] si;
  output [11:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17;
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N17) );
  SELECT_OP C63 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C71 ( .A(N3), .B(N2), .Z(N16) );
  GTECH_NOT I_2 ( .A(N16), .Z(N17) );
endmodule


module dff_SIZE13 ( din, clk, q, se, si, so );
  input [12:0] din;
  output [12:0] q;
  input [12:0] si;
  output [12:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15;
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C23 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module fpu_add_exp_dp ( inq_in1, inq_in2, inq_op, inq_op_7, a1stg_step, 
        a1stg_faddsubd, a1stg_faddsubs, a1stg_fsdtoix, a6stg_step, a1stg_fstod, 
        a1stg_fdtos, a1stg_fstoi, a1stg_fstox, a1stg_fdtoi, a1stg_fdtox, 
        a2stg_fsdtoix_fdtos, a2stg_faddsubop, a2stg_fitos, a2stg_fitod, 
        a2stg_fxtos, a2stg_fxtod, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add, 
        a3stg_inc_exp_inv, a3stg_same_exp_inv, a3stg_dec_exp_inv, 
        a3stg_faddsubop, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, 
        a4stg_shl_cnt, a4stg_denorm_inv, a4stg_rndadd_cout, add_exp_out_expinc, 
        add_exp_out_exp, add_exp_out_exp1, a4stg_in_of, add_exp_out_expadd, 
        a4stg_dblop, a4stg_to_0_inv, fadd_clken_l, rclk, a1stg_expadd3_11, 
        a1stg_expadd1_11_0, a1stg_expadd4_inv, a1stg_expadd2_5_0, a2stg_exp, 
        a2stg_expadd, a3stg_exp_10_0, a4stg_exp_11_0, add_exp_out, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [1:0] inq_op;
  input [5:0] a4stg_shl_cnt;
  output [11:0] a1stg_expadd1_11_0;
  output [10:0] a1stg_expadd4_inv;
  output [5:0] a1stg_expadd2_5_0;
  output [11:0] a2stg_exp;
  output [12:0] a2stg_expadd;
  output [10:0] a3stg_exp_10_0;
  output [11:0] a4stg_exp_11_0;
  output [10:0] add_exp_out;
  input inq_op_7, a1stg_step, a1stg_faddsubd, a1stg_faddsubs, a1stg_fsdtoix,
         a6stg_step, a1stg_fstod, a1stg_fdtos, a1stg_fstoi, a1stg_fstox,
         a1stg_fdtoi, a1stg_fdtox, a2stg_fsdtoix_fdtos, a2stg_faddsubop,
         a2stg_fitos, a2stg_fitod, a2stg_fxtos, a2stg_fxtod, a3stg_exp_7ff,
         a3stg_exp_ff, a3stg_exp_add, a3stg_inc_exp_inv, a3stg_same_exp_inv,
         a3stg_dec_exp_inv, a3stg_faddsubop, a3stg_fdtos_inv,
         a4stg_fixtos_fxtod_inv, a4stg_denorm_inv, a4stg_rndadd_cout,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1, a4stg_in_of,
         add_exp_out_expadd, a4stg_dblop, a4stg_to_0_inv, fadd_clken_l, rclk,
         se, si;
  output a1stg_expadd3_11, so;
  wire   se_l, clk, a1stg_op_7_0, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458,
         N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667,
         N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678,
         N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689,
         N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722,
         N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733,
         N734, N735, N736, net15823, net15824, net15825, net15826, net15827,
         net15828, net15829, net15830, net15831, net15832, net15833, net15834,
         net15835, net15836, net15837, net15838, net15839, net15840, net15841,
         net15842, net15843, net15844, net15845, net15846, net15847, net15848,
         net15849, net15850, net15851, net15852, net15853, net15854, net15855,
         net15856, net15857, net15858, net15859, net15860, net15861, net15862,
         net15863, net15864, net15865, net15866, net15867, net15868, net15869,
         net15870, net15871, net15872, net15873, net15874, net15875, net15876,
         net15877, net15878, net15879, net15880, net15881, net15882, net15883,
         net15884, net15885, net15886, net15887, net15888, net15889, net15890,
         net15891, net15892, net15893, net15894, net15895, net15896, net15897,
         net15898, net15899, net15900, net15901, net15902, net15903, net15904,
         net15905, net15906, net15907, net15908, net15909, net15910, net15911,
         net15912, net15913, net15914, net15915, net15916, net15917, net15918,
         net15919, net15920, net15921, net15922, net15923, net15924, net15925,
         net15926, net15927, net15928, net15929, net15930, net15931, net15932,
         net15933, net15934, net15935, net15936, net15937, net15938, net15939,
         net15940, net15941, net15942, net15943, net15944, net15945, net15946,
         net15947, net15948, net15949, net15950, net15951, net15952, net15953,
         net15954, net15955, net15956, net15957, net15958, net15959, net15960,
         net15961, net15962, net15963, net15964, net15965, net15966, net15967,
         net15968, net15969, net15970, net15971, net15972, net15973, net15974,
         net15975, net15976, net15977, net15978, net15979, net15980, net15981,
         net15982, net15983, net15984, net15985, net15986, net15987, net15988,
         net15989, net15990, net15991, net15992, net15993, net15994, net15995,
         net15996, net15997, net15998, net15999, net16000, net16001, net16002,
         net16003, net16004, net16005, net16006, net16007, net16008, net16009,
         net16010, net16011, net16012, net16013, net16014, net16015, net16016,
         net16017, net16018, net16019, net16020, net16021, net16022, net16023,
         net16024, net16025, net16026, net16027, net16028, net16029, net16030,
         net16031, net16032, net16033, net16034, net16035, net16036, net16037,
         net16038, net16039, net16040, net16041, net16042, net16043, net16044,
         net16045, net16046, net16047, net16048, net16049, net16050, net16051,
         net16052, net16053, net16054, net16055, net16056, net16057, net16058,
         net16059, net16060, net16061, net16062, net16063, net16064, net16065,
         net16066, net16067, net16068, net16069, net16070, net16071, net16072,
         net16073, net16074, net16075, net16076, net16077, net16078, net16079,
         net16080, net16081, net16082, net16083, net16084, net16085, net16086,
         net16087, net16088, net16089, net16090, net16091, net16092, net16093,
         net16094, net16095, net16096, net16097, net16098, net16099, net16100,
         net16101, net16102, net16103, net16104, net16105, net16881, net16882,
         net16883, net16884, net16885, net16886, net16887, net16888, net16889,
         net16890, net16891;
  wire   [62:52] a1stg_in1;
  wire   [62:52] a1stg_in1a;
  wire   [62:52] a1stg_in2;
  wire   [62:52] a1stg_in2a;
  wire   [12:0] a1stg_dp_sngop;
  wire   [12:0] a1stg_dp_sngopa;
  wire   [12:0] a1stg_dp_dblop;
  wire   [12:0] a1stg_dp_dblopa;
  wire   [9:7] a1stg_op_7;
  wire   [10:0] a1stg_expadd3_in1;
  wire   [10:0] a1stg_expadd3_in2_in;
  wire   [10:0] a1stg_expadd3_in2;
  wire   [10:0] a1stg_expadd1_in1;
  wire   [10:0] a1stg_expadd1_in2;
  wire   [12:12] a1stg_expadd1;
  wire   [10:0] a1stg_expadd4_in1;
  wire   [10:0] a1stg_expadd4_in2;
  wire   [10:0] a1stg_expadd4;
  wire   [10:0] a1stg_expadd2_in1;
  wire   [11:6] a1stg_expadd2;
  wire   [12:0] a2stg_exp_in;
  wire   [12:0] a2stg_expa;
  wire   [12:5] a2stg_expadd_in2_in;
  wire   [12:0] a2stg_expadd_in2;
  wire   [12:0] a3stg_exp_in;
  wire   [12:11] a3stg_exp;
  wire   [12:0] a3stg_exp_plus1;
  wire   [12:0] a3stg_exp_minus1;
  wire   [12:0] a4stg_exp_pre1_in;
  wire   [12:0] a4stg_exp_pre1;
  wire   [12:0] a4stg_exp_pre3_in;
  wire   [12:0] a4stg_exp_pre3;
  wire   [12:0] a4stg_expshl;
  wire   [12:12] a4stg_exp;
  wire   [12:0] a4stg_exp_pre2_in;
  wire   [12:0] a4stg_exp_pre2;
  wire   [12:0] a4stg_exp_pre4_in;
  wire   [12:0] a4stg_exp_pre4;
  wire   [12:0] a4stg_exp2;
  wire   [10:0] a4stg_expinc;
  wire   [5:0] a4stg_expadd_in2;
  wire   [12:0] a4stg_expadd;
  wire   [10:0] add_exp_out_in1;
  wire   [10:0] add_exp_out1;
  wire   [10:0] add_exp_out_in2;
  wire   [10:0] add_exp_out2;
  wire   [10:0] add_exp_out_in3;
  wire   [10:0] add_exp_out3;
  wire   [10:0] add_exp_out4;

  clken_buf ckbuf_add_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fadd_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE11 i_a1stg_in1 ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1), .se(se), .si({net16095, net16096, net16097, net16098, 
        net16099, net16100, net16101, net16102, net16103, net16104, net16105})
         );
  dffe_SIZE11 i_a1stg_in1a ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1a), .se(se), .si({net16084, net16085, net16086, net16087, 
        net16088, net16089, net16090, net16091, net16092, net16093, net16094})
         );
  dffe_SIZE11 i_a1stg_in2 ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2), .se(se), .si({net16073, net16074, net16075, net16076, 
        net16077, net16078, net16079, net16080, net16081, net16082, net16083})
         );
  dffe_SIZE11 i_a1stg_in2a ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2a), .se(se), .si({net16062, net16063, net16064, net16065, 
        net16066, net16067, net16068, net16069, net16070, net16071, net16072})
         );
  dffe_SIZE13 i_a1stg_dp_sngop ( .din({inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0]}), .en(a1stg_step), .clk(
        clk), .q(a1stg_dp_sngop), .se(se), .si({net16049, net16050, net16051, 
        net16052, net16053, net16054, net16055, net16056, net16057, net16058, 
        net16059, net16060, net16061}) );
  dffe_SIZE13 i_a1stg_dp_sngopa ( .din({inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0], inq_op[0], inq_op[0], inq_op[0]}), .en(a1stg_step), .clk(
        clk), .q(a1stg_dp_sngopa), .se(se), .si({net16036, net16037, net16038, 
        net16039, net16040, net16041, net16042, net16043, net16044, net16045, 
        net16046, net16047, net16048}) );
  dffe_SIZE13 i_a1stg_dp_dblop ( .din({inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1]}), .en(a1stg_step), .clk(
        clk), .q(a1stg_dp_dblop), .se(se), .si({net16023, net16024, net16025, 
        net16026, net16027, net16028, net16029, net16030, net16031, net16032, 
        net16033, net16034, net16035}) );
  dffe_SIZE13 i_a1stg_dp_dblopa ( .din({inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1], inq_op[1], inq_op[1], inq_op[1]}), .en(a1stg_step), .clk(
        clk), .q(a1stg_dp_dblopa), .se(se), .si({net16010, net16011, net16012, 
        net16013, net16014, net16015, net16016, net16017, net16018, net16019, 
        net16020, net16021, net16022}) );
  dffe_SIZE4 i_a1stg_op_7 ( .din({inq_op_7, inq_op_7, inq_op_7, inq_op_7}), 
        .en(a1stg_step), .clk(clk), .q({a1stg_op_7, a1stg_op_7_0}), .se(se), 
        .si({net16006, net16007, net16008, net16009}) );
  dffe_SIZE11 i_a1stg_expadd3_in1 ( .din(inq_in1), .en(a1stg_step), .clk(clk), 
        .q(a1stg_expadd3_in1), .se(se), .si({net15995, net15996, net15997, 
        net15998, net15999, net16000, net16001, net16002, net16003, net16004, 
        net16005}) );
  dffe_SIZE11 i_a1stg_expadd3_in2 ( .din(a1stg_expadd3_in2_in), .en(a1stg_step), .clk(clk), .q(a1stg_expadd3_in2), .se(se), .si({net15984, net15985, net15986, 
        net15987, net15988, net15989, net15990, net15991, net15992, net15993, 
        net15994}) );
  dffe_SIZE12 i_a2stg_exp ( .din(a2stg_exp_in[11:0]), .en(a6stg_step), .clk(
        clk), .q(a2stg_exp), .se(se), .si({net15972, net15973, net15974, 
        net15975, net15976, net15977, net15978, net15979, net15980, net15981, 
        net15982, net15983}) );
  dffe_SIZE13 i_a2stg_expa ( .din(a2stg_exp_in), .en(a6stg_step), .clk(clk), 
        .q(a2stg_expa), .se(se), .si({net15959, net15960, net15961, net15962, 
        net15963, net15964, net15965, net15966, net15967, net15968, net15969, 
        net15970, net15971}) );
  dffe_SIZE13 i_a2stg_expadd2_in2 ( .din({a2stg_expadd_in2_in, a1stg_fdtos, 
        a1stg_fdtos, a1stg_fdtos, a1stg_fdtos, a1stg_fdtos}), .en(a6stg_step), 
        .clk(clk), .q(a2stg_expadd_in2), .se(se), .si({net15946, net15947, 
        net15948, net15949, net15950, net15951, net15952, net15953, net15954, 
        net15955, net15956, net15957, net15958}) );
  dffe_SIZE13 i_a3stg_exp ( .din(a3stg_exp_in), .en(a6stg_step), .clk(clk), 
        .q({a3stg_exp, a3stg_exp_10_0}), .se(se), .si({net15933, net15934, 
        net15935, net15936, net15937, net15938, net15939, net15940, net15941, 
        net15942, net15943, net15944, net15945}) );
  dff_SIZE13 i_a4stg_exp_pre1 ( .din(a4stg_exp_pre1_in), .clk(clk), .q(
        a4stg_exp_pre1), .se(se), .si({net15920, net15921, net15922, net15923, 
        net15924, net15925, net15926, net15927, net15928, net15929, net15930, 
        net15931, net15932}) );
  dff_SIZE13 i_a4stg_exp_pre3 ( .din(a4stg_exp_pre3_in), .clk(clk), .q(
        a4stg_exp_pre3), .se(se), .si({net15907, net15908, net15909, net15910, 
        net15911, net15912, net15913, net15914, net15915, net15916, net15917, 
        net15918, net15919}) );
  dff_SIZE13 i_a4stg_exp_pre2 ( .din(a4stg_exp_pre2_in), .clk(clk), .q(
        a4stg_exp_pre2), .se(se), .si({net15894, net15895, net15896, net15897, 
        net15898, net15899, net15900, net15901, net15902, net15903, net15904, 
        net15905, net15906}) );
  dff_SIZE13 i_a4stg_exp_pre4 ( .din(a4stg_exp_pre4_in), .clk(clk), .q(
        a4stg_exp_pre4), .se(se), .si({net15881, net15882, net15883, net15884, 
        net15885, net15886, net15887, net15888, net15889, net15890, net15891, 
        net15892, net15893}) );
  dffe_SIZE13 i_a4stg_exp2 ( .din({a3stg_exp, a3stg_exp_10_0}), .en(a6stg_step), .clk(clk), .q(a4stg_exp2), .se(se), .si({net15868, net15869, net15870, 
        net15871, net15872, net15873, net15874, net15875, net15876, net15877, 
        net15878, net15879, net15880}) );
  dffe_SIZE11 i_add_exp_out1 ( .din(add_exp_out_in1), .en(a6stg_step), .clk(
        clk), .q(add_exp_out1), .se(se), .si({net15857, net15858, net15859, 
        net15860, net15861, net15862, net15863, net15864, net15865, net15866, 
        net15867}) );
  dffe_SIZE11 i_add_exp_out2 ( .din(add_exp_out_in2), .en(a6stg_step), .clk(
        clk), .q(add_exp_out2), .se(se), .si({net15846, net15847, net15848, 
        net15849, net15850, net15851, net15852, net15853, net15854, net15855, 
        net15856}) );
  dffe_SIZE11 i_add_exp_out3 ( .din(add_exp_out_in3), .en(a6stg_step), .clk(
        clk), .q(add_exp_out3), .se(se), .si({net15835, net15836, net15837, 
        net15838, net15839, net15840, net15841, net15842, net15843, net15844, 
        net15845}) );
  dffe_SIZE11 i_add_exp_out4 ( .din({a4stg_rndadd_cout, a4stg_rndadd_cout, 
        a4stg_rndadd_cout, a4stg_rndadd_cout, a4stg_rndadd_cout, 
        a4stg_rndadd_cout, a4stg_rndadd_cout, a4stg_rndadd_cout, 
        a4stg_rndadd_cout, a4stg_rndadd_cout, a4stg_rndadd_cout}), .en(
        a6stg_step), .clk(clk), .q(add_exp_out4), .se(se), .si({net15824, 
        net15825, net15826, net15827, net15828, net15829, net15830, net15831, 
        net15832, net15833, net15834}) );
  ADD_UNS_OP add_501 ( .A(a2stg_expa), .B(a2stg_expadd_in2), .Z({N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39, N38, N37}) );
  ADD_UNS_OP add_501_2 ( .A({N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37}), .B(a2stg_fsdtoix_fdtos), .Z(a2stg_expadd) );
  ADD_UNS_OP add_405 ( .A(a1stg_expadd4_in1), .B(a1stg_expadd4_in2), .Z({N35, 
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25}) );
  ADD_UNS_OP add_415 ( .A(a1stg_expadd2_in1), .B(1'b1), .Z({a1stg_expadd2, 
        a1stg_expadd2_5_0}) );
  ADD_UNS_OP add_546 ( .A({a3stg_exp, a3stg_exp_10_0}), .B(1'b1), .Z(
        a3stg_exp_plus1) );
  SUB_UNS_OP sub_548 ( .A({a3stg_exp, a3stg_exp_10_0}), .B(1'b1), .Z(
        a3stg_exp_minus1) );
  ADD_UNS_OP add_390 ( .A(a1stg_expadd1_in1), .B({1'b1, 1'b1, 
        a1stg_expadd1_in2}), .Z({N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12}) );
  ADD_UNS_OP add_654 ( .A(a4stg_exp2), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, a4stg_expadd_in2}), .Z({N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50}) );
  ADD_UNS_OP add_373 ( .A(a1stg_expadd3_in1), .B({1'b1, a1stg_expadd3_in2}), 
        .Z({N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  ADD_UNS_OP add_641 ( .A(a4stg_exp_11_0[10:0]), .B(1'b1), .Z(a4stg_expinc) );
  ADD_UNS_OP add_405_2 ( .A({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25}), .B(1'b1), .Z(a1stg_expadd4) );
  ADD_UNS_OP add_390_2 ( .A({N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12}), .B(1'b1), .Z({a1stg_expadd1[12], a1stg_expadd1_11_0})
         );
  ADD_UNS_OP add_654_2 ( .A({N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50}), .B(1'b1), .Z(a4stg_expadd) );
  ADD_UNS_OP add_373_2 ( .A({N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), .B(1'b1), .Z({a1stg_expadd3_11, net16881, net16882, net16883, net16884, 
        net16885, net16886, net16887, net16888, net16889, net16890, net16891})
         );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_NOT I_1 ( .A(inq_in2[62]), .Z(a1stg_expadd3_in2_in[10]) );
  GTECH_NOT I_2 ( .A(inq_in2[61]), .Z(a1stg_expadd3_in2_in[9]) );
  GTECH_NOT I_3 ( .A(inq_in2[60]), .Z(a1stg_expadd3_in2_in[8]) );
  GTECH_NOT I_4 ( .A(inq_in2[59]), .Z(a1stg_expadd3_in2_in[7]) );
  GTECH_NOT I_5 ( .A(inq_in2[58]), .Z(a1stg_expadd3_in2_in[6]) );
  GTECH_NOT I_6 ( .A(inq_in2[57]), .Z(a1stg_expadd3_in2_in[5]) );
  GTECH_NOT I_7 ( .A(inq_in2[56]), .Z(a1stg_expadd3_in2_in[4]) );
  GTECH_NOT I_8 ( .A(inq_in2[55]), .Z(a1stg_expadd3_in2_in[3]) );
  GTECH_NOT I_9 ( .A(N63), .Z(a1stg_expadd3_in2_in[2]) );
  GTECH_AND2 C258 ( .A(inq_in2[54]), .B(inq_op[1]), .Z(N63) );
  GTECH_NOT I_10 ( .A(N64), .Z(a1stg_expadd3_in2_in[1]) );
  GTECH_AND2 C260 ( .A(inq_in2[53]), .B(inq_op[1]), .Z(N64) );
  GTECH_NOT I_11 ( .A(N65), .Z(a1stg_expadd3_in2_in[0]) );
  GTECH_AND2 C262 ( .A(inq_in2[52]), .B(inq_op[1]), .Z(N65) );
  GTECH_AND2 C263 ( .A(a1stg_dp_dblopa[10]), .B(a1stg_in1[62]), .Z(
        a1stg_expadd1_in1[10]) );
  GTECH_OR2 C264 ( .A(N66), .B(a1stg_op_7[9]), .Z(a1stg_expadd1_in1[9]) );
  GTECH_AND2 C265 ( .A(a1stg_dp_dblopa[9]), .B(a1stg_in1[61]), .Z(N66) );
  GTECH_OR2 C266 ( .A(N67), .B(a1stg_op_7[8]), .Z(a1stg_expadd1_in1[8]) );
  GTECH_AND2 C267 ( .A(a1stg_dp_dblopa[8]), .B(a1stg_in1[60]), .Z(N67) );
  GTECH_OR2 C268 ( .A(N70), .B(a1stg_op_7[7]), .Z(a1stg_expadd1_in1[7]) );
  GTECH_OR2 C269 ( .A(N68), .B(N69), .Z(N70) );
  GTECH_AND2 C270 ( .A(a1stg_dp_dblopa[7]), .B(a1stg_in1[59]), .Z(N68) );
  GTECH_AND2 C271 ( .A(a1stg_dp_sngopa[7]), .B(a1stg_in1[62]), .Z(N69) );
  GTECH_OR2 C272 ( .A(N71), .B(N72), .Z(a1stg_expadd1_in1[6]) );
  GTECH_AND2 C273 ( .A(a1stg_dp_dblopa[6]), .B(a1stg_in1[58]), .Z(N71) );
  GTECH_AND2 C274 ( .A(a1stg_dp_sngopa[6]), .B(a1stg_in1[61]), .Z(N72) );
  GTECH_OR2 C275 ( .A(N73), .B(N74), .Z(a1stg_expadd1_in1[5]) );
  GTECH_AND2 C276 ( .A(a1stg_dp_dblopa[5]), .B(a1stg_in1[57]), .Z(N73) );
  GTECH_AND2 C277 ( .A(a1stg_dp_sngopa[5]), .B(a1stg_in1[60]), .Z(N74) );
  GTECH_OR2 C278 ( .A(N75), .B(N76), .Z(a1stg_expadd1_in1[4]) );
  GTECH_AND2 C279 ( .A(a1stg_dp_dblopa[4]), .B(a1stg_in1[56]), .Z(N75) );
  GTECH_AND2 C280 ( .A(a1stg_dp_sngopa[4]), .B(a1stg_in1[59]), .Z(N76) );
  GTECH_OR2 C281 ( .A(N77), .B(N78), .Z(a1stg_expadd1_in1[3]) );
  GTECH_AND2 C282 ( .A(a1stg_dp_dblopa[3]), .B(a1stg_in1[55]), .Z(N77) );
  GTECH_AND2 C283 ( .A(a1stg_dp_sngopa[3]), .B(a1stg_in1[58]), .Z(N78) );
  GTECH_OR2 C284 ( .A(N79), .B(N80), .Z(a1stg_expadd1_in1[2]) );
  GTECH_AND2 C285 ( .A(a1stg_dp_dblopa[2]), .B(a1stg_in1[54]), .Z(N79) );
  GTECH_AND2 C286 ( .A(a1stg_dp_sngopa[2]), .B(a1stg_in1[57]), .Z(N80) );
  GTECH_OR2 C287 ( .A(N81), .B(N82), .Z(a1stg_expadd1_in1[1]) );
  GTECH_AND2 C288 ( .A(a1stg_dp_dblopa[1]), .B(a1stg_in1[53]), .Z(N81) );
  GTECH_AND2 C289 ( .A(a1stg_dp_sngopa[1]), .B(a1stg_in1[56]), .Z(N82) );
  GTECH_OR2 C290 ( .A(N85), .B(a1stg_op_7_0), .Z(a1stg_expadd1_in1[0]) );
  GTECH_OR2 C291 ( .A(N83), .B(N84), .Z(N85) );
  GTECH_AND2 C292 ( .A(a1stg_dp_dblopa[0]), .B(a1stg_in1[52]), .Z(N83) );
  GTECH_AND2 C293 ( .A(a1stg_dp_sngopa[0]), .B(a1stg_in1[55]), .Z(N84) );
  GTECH_NOT I_12 ( .A(N86), .Z(a1stg_expadd1_in2[10]) );
  GTECH_AND2 C295 ( .A(a1stg_dp_dblop[10]), .B(a1stg_in2[62]), .Z(N86) );
  GTECH_NOT I_13 ( .A(N87), .Z(a1stg_expadd1_in2[9]) );
  GTECH_AND2 C297 ( .A(a1stg_dp_dblop[9]), .B(a1stg_in2[61]), .Z(N87) );
  GTECH_NOT I_14 ( .A(N88), .Z(a1stg_expadd1_in2[8]) );
  GTECH_AND2 C299 ( .A(a1stg_dp_dblop[8]), .B(a1stg_in2[60]), .Z(N88) );
  GTECH_NOT I_15 ( .A(N91), .Z(a1stg_expadd1_in2[7]) );
  GTECH_OR2 C301 ( .A(N89), .B(N90), .Z(N91) );
  GTECH_AND2 C302 ( .A(a1stg_dp_dblop[7]), .B(a1stg_in2[59]), .Z(N89) );
  GTECH_AND2 C303 ( .A(a1stg_dp_sngop[7]), .B(a1stg_in2[62]), .Z(N90) );
  GTECH_NOT I_16 ( .A(N94), .Z(a1stg_expadd1_in2[6]) );
  GTECH_OR2 C305 ( .A(N92), .B(N93), .Z(N94) );
  GTECH_AND2 C306 ( .A(a1stg_dp_dblop[6]), .B(a1stg_in2[58]), .Z(N92) );
  GTECH_AND2 C307 ( .A(a1stg_dp_sngop[6]), .B(a1stg_in2[61]), .Z(N93) );
  GTECH_NOT I_17 ( .A(N97), .Z(a1stg_expadd1_in2[5]) );
  GTECH_OR2 C309 ( .A(N95), .B(N96), .Z(N97) );
  GTECH_AND2 C310 ( .A(a1stg_dp_dblop[5]), .B(a1stg_in2[57]), .Z(N95) );
  GTECH_AND2 C311 ( .A(a1stg_dp_sngop[5]), .B(a1stg_in2[60]), .Z(N96) );
  GTECH_NOT I_18 ( .A(N100), .Z(a1stg_expadd1_in2[4]) );
  GTECH_OR2 C313 ( .A(N98), .B(N99), .Z(N100) );
  GTECH_AND2 C314 ( .A(a1stg_dp_dblop[4]), .B(a1stg_in2[56]), .Z(N98) );
  GTECH_AND2 C315 ( .A(a1stg_dp_sngop[4]), .B(a1stg_in2[59]), .Z(N99) );
  GTECH_NOT I_19 ( .A(N103), .Z(a1stg_expadd1_in2[3]) );
  GTECH_OR2 C317 ( .A(N101), .B(N102), .Z(N103) );
  GTECH_AND2 C318 ( .A(a1stg_dp_dblop[3]), .B(a1stg_in2[55]), .Z(N101) );
  GTECH_AND2 C319 ( .A(a1stg_dp_sngop[3]), .B(a1stg_in2[58]), .Z(N102) );
  GTECH_NOT I_20 ( .A(N106), .Z(a1stg_expadd1_in2[2]) );
  GTECH_OR2 C321 ( .A(N104), .B(N105), .Z(N106) );
  GTECH_AND2 C322 ( .A(a1stg_dp_dblop[2]), .B(a1stg_in2[54]), .Z(N104) );
  GTECH_AND2 C323 ( .A(a1stg_dp_sngop[2]), .B(a1stg_in2[57]), .Z(N105) );
  GTECH_NOT I_21 ( .A(N109), .Z(a1stg_expadd1_in2[1]) );
  GTECH_OR2 C325 ( .A(N107), .B(N108), .Z(N109) );
  GTECH_AND2 C326 ( .A(a1stg_dp_dblop[1]), .B(a1stg_in2[53]), .Z(N107) );
  GTECH_AND2 C327 ( .A(a1stg_dp_sngop[1]), .B(a1stg_in2[56]), .Z(N108) );
  GTECH_NOT I_22 ( .A(N112), .Z(a1stg_expadd1_in2[0]) );
  GTECH_OR2 C329 ( .A(N110), .B(N111), .Z(N112) );
  GTECH_AND2 C330 ( .A(a1stg_dp_dblop[0]), .B(a1stg_in2[52]), .Z(N110) );
  GTECH_AND2 C331 ( .A(a1stg_dp_sngop[0]), .B(a1stg_in2[55]), .Z(N111) );
  GTECH_AND2 C332 ( .A(a1stg_dp_dblopa[10]), .B(a1stg_in2a[62]), .Z(
        a1stg_expadd4_in1[10]) );
  GTECH_AND2 C333 ( .A(a1stg_dp_dblopa[9]), .B(a1stg_in2a[61]), .Z(
        a1stg_expadd4_in1[9]) );
  GTECH_AND2 C334 ( .A(a1stg_dp_dblopa[8]), .B(a1stg_in2a[60]), .Z(
        a1stg_expadd4_in1[8]) );
  GTECH_OR2 C335 ( .A(N113), .B(N114), .Z(a1stg_expadd4_in1[7]) );
  GTECH_AND2 C336 ( .A(a1stg_dp_dblopa[7]), .B(a1stg_in2a[59]), .Z(N113) );
  GTECH_AND2 C337 ( .A(a1stg_dp_sngopa[7]), .B(a1stg_in2a[62]), .Z(N114) );
  GTECH_OR2 C338 ( .A(N115), .B(N116), .Z(a1stg_expadd4_in1[6]) );
  GTECH_AND2 C339 ( .A(a1stg_dp_dblopa[6]), .B(a1stg_in2a[58]), .Z(N115) );
  GTECH_AND2 C340 ( .A(a1stg_dp_sngopa[6]), .B(a1stg_in2a[61]), .Z(N116) );
  GTECH_OR2 C341 ( .A(N117), .B(N118), .Z(a1stg_expadd4_in1[5]) );
  GTECH_AND2 C342 ( .A(a1stg_dp_dblopa[5]), .B(a1stg_in2a[57]), .Z(N117) );
  GTECH_AND2 C343 ( .A(a1stg_dp_sngopa[5]), .B(a1stg_in2a[60]), .Z(N118) );
  GTECH_OR2 C344 ( .A(N119), .B(N120), .Z(a1stg_expadd4_in1[4]) );
  GTECH_AND2 C345 ( .A(a1stg_dp_dblopa[4]), .B(a1stg_in2a[56]), .Z(N119) );
  GTECH_AND2 C346 ( .A(a1stg_dp_sngopa[4]), .B(a1stg_in2a[59]), .Z(N120) );
  GTECH_OR2 C347 ( .A(N121), .B(N122), .Z(a1stg_expadd4_in1[3]) );
  GTECH_AND2 C348 ( .A(a1stg_dp_dblopa[3]), .B(a1stg_in2a[55]), .Z(N121) );
  GTECH_AND2 C349 ( .A(a1stg_dp_sngopa[3]), .B(a1stg_in2a[58]), .Z(N122) );
  GTECH_OR2 C350 ( .A(N123), .B(N124), .Z(a1stg_expadd4_in1[2]) );
  GTECH_AND2 C351 ( .A(a1stg_dp_dblopa[2]), .B(a1stg_in2a[54]), .Z(N123) );
  GTECH_AND2 C352 ( .A(a1stg_dp_sngopa[2]), .B(a1stg_in2a[57]), .Z(N124) );
  GTECH_OR2 C353 ( .A(N125), .B(N126), .Z(a1stg_expadd4_in1[1]) );
  GTECH_AND2 C354 ( .A(a1stg_dp_dblopa[1]), .B(a1stg_in2a[53]), .Z(N125) );
  GTECH_AND2 C355 ( .A(a1stg_dp_sngopa[1]), .B(a1stg_in2a[56]), .Z(N126) );
  GTECH_OR2 C356 ( .A(N127), .B(N128), .Z(a1stg_expadd4_in1[0]) );
  GTECH_AND2 C357 ( .A(a1stg_dp_dblopa[0]), .B(a1stg_in2a[52]), .Z(N127) );
  GTECH_AND2 C358 ( .A(a1stg_dp_sngopa[0]), .B(a1stg_in2a[55]), .Z(N128) );
  GTECH_NOT I_23 ( .A(N129), .Z(a1stg_expadd4_in2[10]) );
  GTECH_AND2 C360 ( .A(a1stg_dp_dblop[10]), .B(a1stg_in1a[62]), .Z(N129) );
  GTECH_NOT I_24 ( .A(N130), .Z(a1stg_expadd4_in2[9]) );
  GTECH_AND2 C362 ( .A(a1stg_dp_dblop[9]), .B(a1stg_in1a[61]), .Z(N130) );
  GTECH_NOT I_25 ( .A(N131), .Z(a1stg_expadd4_in2[8]) );
  GTECH_AND2 C364 ( .A(a1stg_dp_dblop[8]), .B(a1stg_in1a[60]), .Z(N131) );
  GTECH_NOT I_26 ( .A(N134), .Z(a1stg_expadd4_in2[7]) );
  GTECH_OR2 C366 ( .A(N132), .B(N133), .Z(N134) );
  GTECH_AND2 C367 ( .A(a1stg_dp_dblop[7]), .B(a1stg_in1a[59]), .Z(N132) );
  GTECH_AND2 C368 ( .A(a1stg_dp_sngop[7]), .B(a1stg_in1a[62]), .Z(N133) );
  GTECH_NOT I_27 ( .A(N137), .Z(a1stg_expadd4_in2[6]) );
  GTECH_OR2 C370 ( .A(N135), .B(N136), .Z(N137) );
  GTECH_AND2 C371 ( .A(a1stg_dp_dblop[6]), .B(a1stg_in1a[58]), .Z(N135) );
  GTECH_AND2 C372 ( .A(a1stg_dp_sngop[6]), .B(a1stg_in1a[61]), .Z(N136) );
  GTECH_NOT I_28 ( .A(N140), .Z(a1stg_expadd4_in2[5]) );
  GTECH_OR2 C374 ( .A(N138), .B(N139), .Z(N140) );
  GTECH_AND2 C375 ( .A(a1stg_dp_dblop[5]), .B(a1stg_in1a[57]), .Z(N138) );
  GTECH_AND2 C376 ( .A(a1stg_dp_sngop[5]), .B(a1stg_in1a[60]), .Z(N139) );
  GTECH_NOT I_29 ( .A(N143), .Z(a1stg_expadd4_in2[4]) );
  GTECH_OR2 C378 ( .A(N141), .B(N142), .Z(N143) );
  GTECH_AND2 C379 ( .A(a1stg_dp_dblop[4]), .B(a1stg_in1a[56]), .Z(N141) );
  GTECH_AND2 C380 ( .A(a1stg_dp_sngop[4]), .B(a1stg_in1a[59]), .Z(N142) );
  GTECH_NOT I_30 ( .A(N146), .Z(a1stg_expadd4_in2[3]) );
  GTECH_OR2 C382 ( .A(N144), .B(N145), .Z(N146) );
  GTECH_AND2 C383 ( .A(a1stg_dp_dblop[3]), .B(a1stg_in1a[55]), .Z(N144) );
  GTECH_AND2 C384 ( .A(a1stg_dp_sngop[3]), .B(a1stg_in1a[58]), .Z(N145) );
  GTECH_NOT I_31 ( .A(N149), .Z(a1stg_expadd4_in2[2]) );
  GTECH_OR2 C386 ( .A(N147), .B(N148), .Z(N149) );
  GTECH_AND2 C387 ( .A(a1stg_dp_dblop[2]), .B(a1stg_in1a[54]), .Z(N147) );
  GTECH_AND2 C388 ( .A(a1stg_dp_sngop[2]), .B(a1stg_in1a[57]), .Z(N148) );
  GTECH_NOT I_32 ( .A(N152), .Z(a1stg_expadd4_in2[1]) );
  GTECH_OR2 C390 ( .A(N150), .B(N151), .Z(N152) );
  GTECH_AND2 C391 ( .A(a1stg_dp_dblop[1]), .B(a1stg_in1a[53]), .Z(N150) );
  GTECH_AND2 C392 ( .A(a1stg_dp_sngop[1]), .B(a1stg_in1a[56]), .Z(N151) );
  GTECH_NOT I_33 ( .A(N155), .Z(a1stg_expadd4_in2[0]) );
  GTECH_OR2 C394 ( .A(N153), .B(N154), .Z(N155) );
  GTECH_AND2 C395 ( .A(a1stg_dp_dblop[0]), .B(a1stg_in1a[52]), .Z(N153) );
  GTECH_AND2 C396 ( .A(a1stg_dp_sngop[0]), .B(a1stg_in1a[55]), .Z(N154) );
  GTECH_NOT I_34 ( .A(a1stg_expadd4[10]), .Z(a1stg_expadd4_inv[10]) );
  GTECH_NOT I_35 ( .A(a1stg_expadd4[9]), .Z(a1stg_expadd4_inv[9]) );
  GTECH_NOT I_36 ( .A(a1stg_expadd4[8]), .Z(a1stg_expadd4_inv[8]) );
  GTECH_NOT I_37 ( .A(a1stg_expadd4[7]), .Z(a1stg_expadd4_inv[7]) );
  GTECH_NOT I_38 ( .A(a1stg_expadd4[6]), .Z(a1stg_expadd4_inv[6]) );
  GTECH_NOT I_39 ( .A(a1stg_expadd4[5]), .Z(a1stg_expadd4_inv[5]) );
  GTECH_NOT I_40 ( .A(a1stg_expadd4[4]), .Z(a1stg_expadd4_inv[4]) );
  GTECH_NOT I_41 ( .A(a1stg_expadd4[3]), .Z(a1stg_expadd4_inv[3]) );
  GTECH_NOT I_42 ( .A(a1stg_expadd4[2]), .Z(a1stg_expadd4_inv[2]) );
  GTECH_NOT I_43 ( .A(a1stg_expadd4[1]), .Z(a1stg_expadd4_inv[1]) );
  GTECH_NOT I_44 ( .A(a1stg_expadd4[0]), .Z(a1stg_expadd4_inv[0]) );
  GTECH_AND2 C408 ( .A(a1stg_dp_dblopa[10]), .B(a1stg_in2a[62]), .Z(
        a1stg_expadd2_in1[10]) );
  GTECH_AND2 C409 ( .A(a1stg_dp_dblopa[9]), .B(a1stg_in2a[61]), .Z(
        a1stg_expadd2_in1[9]) );
  GTECH_AND2 C410 ( .A(a1stg_dp_dblopa[8]), .B(a1stg_in2a[60]), .Z(
        a1stg_expadd2_in1[8]) );
  GTECH_OR2 C411 ( .A(N156), .B(N157), .Z(a1stg_expadd2_in1[7]) );
  GTECH_AND2 C412 ( .A(a1stg_dp_dblopa[7]), .B(a1stg_in2a[59]), .Z(N156) );
  GTECH_AND2 C413 ( .A(a1stg_dp_sngopa[7]), .B(a1stg_in2a[62]), .Z(N157) );
  GTECH_OR2 C414 ( .A(N158), .B(N159), .Z(a1stg_expadd2_in1[6]) );
  GTECH_AND2 C415 ( .A(a1stg_dp_dblopa[6]), .B(a1stg_in2a[58]), .Z(N158) );
  GTECH_AND2 C416 ( .A(a1stg_dp_sngopa[6]), .B(a1stg_in2a[61]), .Z(N159) );
  GTECH_OR2 C417 ( .A(N160), .B(N161), .Z(a1stg_expadd2_in1[5]) );
  GTECH_AND2 C418 ( .A(a1stg_dp_dblopa[5]), .B(a1stg_in2a[57]), .Z(N160) );
  GTECH_AND2 C419 ( .A(a1stg_dp_sngopa[5]), .B(a1stg_in2a[60]), .Z(N161) );
  GTECH_OR2 C420 ( .A(N162), .B(N163), .Z(a1stg_expadd2_in1[4]) );
  GTECH_AND2 C421 ( .A(a1stg_dp_dblopa[4]), .B(a1stg_in2a[56]), .Z(N162) );
  GTECH_AND2 C422 ( .A(a1stg_dp_sngopa[4]), .B(a1stg_in2a[59]), .Z(N163) );
  GTECH_OR2 C423 ( .A(N164), .B(N165), .Z(a1stg_expadd2_in1[3]) );
  GTECH_AND2 C424 ( .A(a1stg_dp_dblopa[3]), .B(a1stg_in2a[55]), .Z(N164) );
  GTECH_AND2 C425 ( .A(a1stg_dp_sngopa[3]), .B(a1stg_in2a[58]), .Z(N165) );
  GTECH_OR2 C426 ( .A(N166), .B(N167), .Z(a1stg_expadd2_in1[2]) );
  GTECH_AND2 C427 ( .A(a1stg_dp_dblopa[2]), .B(a1stg_in2a[54]), .Z(N166) );
  GTECH_AND2 C428 ( .A(a1stg_dp_sngopa[2]), .B(a1stg_in2a[57]), .Z(N167) );
  GTECH_OR2 C429 ( .A(N168), .B(N169), .Z(a1stg_expadd2_in1[1]) );
  GTECH_AND2 C430 ( .A(a1stg_dp_dblopa[1]), .B(a1stg_in2a[53]), .Z(N168) );
  GTECH_AND2 C431 ( .A(a1stg_dp_sngopa[1]), .B(a1stg_in2a[56]), .Z(N169) );
  GTECH_OR2 C432 ( .A(N170), .B(N171), .Z(a1stg_expadd2_in1[0]) );
  GTECH_AND2 C433 ( .A(a1stg_dp_dblopa[0]), .B(a1stg_in2a[52]), .Z(N170) );
  GTECH_AND2 C434 ( .A(a1stg_dp_sngopa[0]), .B(a1stg_in2a[55]), .Z(N171) );
  GTECH_NOT I_45 ( .A(a1stg_expadd1[12]), .Z(N36) );
  GTECH_AND2 C436 ( .A(a1stg_fsdtoix), .B(1'b0), .Z(a2stg_exp_in[12]) );
  GTECH_AND2 C437 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[11]), .Z(
        a2stg_exp_in[11]) );
  GTECH_OR2 C438 ( .A(N178), .B(N179), .Z(a2stg_exp_in[10]) );
  GTECH_OR2 C439 ( .A(N176), .B(N177), .Z(N178) );
  GTECH_OR2 C440 ( .A(N173), .B(N175), .Z(N176) );
  GTECH_AND2 C441 ( .A(N172), .B(a1stg_in1a[62]), .Z(N173) );
  GTECH_AND2 C442 ( .A(a1stg_faddsubd), .B(N36), .Z(N172) );
  GTECH_AND2 C443 ( .A(N174), .B(a1stg_in2[62]), .Z(N175) );
  GTECH_AND2 C444 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N174) );
  GTECH_AND2 C445 ( .A(a1stg_fdtos), .B(a1stg_in2[62]), .Z(N177) );
  GTECH_AND2 C446 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[10]), .Z(N179) );
  GTECH_OR2 C447 ( .A(N186), .B(N187), .Z(a2stg_exp_in[9]) );
  GTECH_OR2 C448 ( .A(N184), .B(N185), .Z(N186) );
  GTECH_OR2 C449 ( .A(N181), .B(N183), .Z(N184) );
  GTECH_AND2 C450 ( .A(N180), .B(a1stg_in1a[61]), .Z(N181) );
  GTECH_AND2 C451 ( .A(a1stg_faddsubd), .B(N36), .Z(N180) );
  GTECH_AND2 C452 ( .A(N182), .B(a1stg_in2[61]), .Z(N183) );
  GTECH_AND2 C453 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N182) );
  GTECH_AND2 C454 ( .A(a1stg_fdtos), .B(a1stg_in2[61]), .Z(N185) );
  GTECH_AND2 C455 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[9]), .Z(N187) );
  GTECH_OR2 C456 ( .A(N194), .B(N195), .Z(a2stg_exp_in[8]) );
  GTECH_OR2 C457 ( .A(N192), .B(N193), .Z(N194) );
  GTECH_OR2 C458 ( .A(N189), .B(N191), .Z(N192) );
  GTECH_AND2 C459 ( .A(N188), .B(a1stg_in1a[60]), .Z(N189) );
  GTECH_AND2 C460 ( .A(a1stg_faddsubd), .B(N36), .Z(N188) );
  GTECH_AND2 C461 ( .A(N190), .B(a1stg_in2[60]), .Z(N191) );
  GTECH_AND2 C462 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N190) );
  GTECH_AND2 C463 ( .A(a1stg_fdtos), .B(a1stg_in2[60]), .Z(N193) );
  GTECH_AND2 C464 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[8]), .Z(N195) );
  GTECH_OR2 C465 ( .A(N210), .B(N211), .Z(a2stg_exp_in[7]) );
  GTECH_OR2 C466 ( .A(N208), .B(N209), .Z(N210) );
  GTECH_OR2 C467 ( .A(N205), .B(N207), .Z(N208) );
  GTECH_OR2 C468 ( .A(N203), .B(N204), .Z(N205) );
  GTECH_OR2 C469 ( .A(N200), .B(N202), .Z(N203) );
  GTECH_OR2 C470 ( .A(N197), .B(N199), .Z(N200) );
  GTECH_AND2 C471 ( .A(N196), .B(a1stg_in1a[59]), .Z(N197) );
  GTECH_AND2 C472 ( .A(a1stg_faddsubd), .B(N36), .Z(N196) );
  GTECH_AND2 C473 ( .A(N198), .B(a1stg_in1a[62]), .Z(N199) );
  GTECH_AND2 C474 ( .A(a1stg_faddsubs), .B(N36), .Z(N198) );
  GTECH_AND2 C475 ( .A(N201), .B(a1stg_in2[59]), .Z(N202) );
  GTECH_AND2 C476 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N201) );
  GTECH_AND2 C477 ( .A(a1stg_fdtos), .B(a1stg_in2[59]), .Z(N204) );
  GTECH_AND2 C478 ( .A(N206), .B(a1stg_in2[62]), .Z(N207) );
  GTECH_AND2 C479 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N206) );
  GTECH_AND2 C480 ( .A(a1stg_fstod), .B(a1stg_in2[62]), .Z(N209) );
  GTECH_AND2 C481 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[7]), .Z(N211) );
  GTECH_OR2 C482 ( .A(N226), .B(N227), .Z(a2stg_exp_in[6]) );
  GTECH_OR2 C483 ( .A(N224), .B(N225), .Z(N226) );
  GTECH_OR2 C484 ( .A(N221), .B(N223), .Z(N224) );
  GTECH_OR2 C485 ( .A(N219), .B(N220), .Z(N221) );
  GTECH_OR2 C486 ( .A(N216), .B(N218), .Z(N219) );
  GTECH_OR2 C487 ( .A(N213), .B(N215), .Z(N216) );
  GTECH_AND2 C488 ( .A(N212), .B(a1stg_in1a[58]), .Z(N213) );
  GTECH_AND2 C489 ( .A(a1stg_faddsubd), .B(N36), .Z(N212) );
  GTECH_AND2 C490 ( .A(N214), .B(a1stg_in1a[61]), .Z(N215) );
  GTECH_AND2 C491 ( .A(a1stg_faddsubs), .B(N36), .Z(N214) );
  GTECH_AND2 C492 ( .A(N217), .B(a1stg_in2[58]), .Z(N218) );
  GTECH_AND2 C493 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N217) );
  GTECH_AND2 C494 ( .A(a1stg_fdtos), .B(a1stg_in2[58]), .Z(N220) );
  GTECH_AND2 C495 ( .A(N222), .B(a1stg_in2[61]), .Z(N223) );
  GTECH_AND2 C496 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N222) );
  GTECH_AND2 C497 ( .A(a1stg_fstod), .B(a1stg_in2[61]), .Z(N225) );
  GTECH_AND2 C498 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2[6]), .Z(N227) );
  GTECH_OR2 C499 ( .A(N242), .B(N243), .Z(a2stg_exp_in[5]) );
  GTECH_OR2 C500 ( .A(N240), .B(N241), .Z(N242) );
  GTECH_OR2 C501 ( .A(N237), .B(N239), .Z(N240) );
  GTECH_OR2 C502 ( .A(N235), .B(N236), .Z(N237) );
  GTECH_OR2 C503 ( .A(N232), .B(N234), .Z(N235) );
  GTECH_OR2 C504 ( .A(N229), .B(N231), .Z(N232) );
  GTECH_AND2 C505 ( .A(N228), .B(a1stg_in1a[57]), .Z(N229) );
  GTECH_AND2 C506 ( .A(a1stg_faddsubd), .B(N36), .Z(N228) );
  GTECH_AND2 C507 ( .A(N230), .B(a1stg_in1a[60]), .Z(N231) );
  GTECH_AND2 C508 ( .A(a1stg_faddsubs), .B(N36), .Z(N230) );
  GTECH_AND2 C509 ( .A(N233), .B(a1stg_in2[57]), .Z(N234) );
  GTECH_AND2 C510 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N233) );
  GTECH_AND2 C511 ( .A(a1stg_fdtos), .B(a1stg_in2[57]), .Z(N236) );
  GTECH_AND2 C512 ( .A(N238), .B(a1stg_in2[60]), .Z(N239) );
  GTECH_AND2 C513 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N238) );
  GTECH_AND2 C514 ( .A(a1stg_fstod), .B(a1stg_in2[60]), .Z(N241) );
  GTECH_AND2 C515 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[5]), .Z(N243) );
  GTECH_OR2 C516 ( .A(N258), .B(N259), .Z(a2stg_exp_in[4]) );
  GTECH_OR2 C517 ( .A(N256), .B(N257), .Z(N258) );
  GTECH_OR2 C518 ( .A(N253), .B(N255), .Z(N256) );
  GTECH_OR2 C519 ( .A(N251), .B(N252), .Z(N253) );
  GTECH_OR2 C520 ( .A(N248), .B(N250), .Z(N251) );
  GTECH_OR2 C521 ( .A(N245), .B(N247), .Z(N248) );
  GTECH_AND2 C522 ( .A(N244), .B(a1stg_in1a[56]), .Z(N245) );
  GTECH_AND2 C523 ( .A(a1stg_faddsubd), .B(N36), .Z(N244) );
  GTECH_AND2 C524 ( .A(N246), .B(a1stg_in1a[59]), .Z(N247) );
  GTECH_AND2 C525 ( .A(a1stg_faddsubs), .B(N36), .Z(N246) );
  GTECH_AND2 C526 ( .A(N249), .B(a1stg_in2[56]), .Z(N250) );
  GTECH_AND2 C527 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N249) );
  GTECH_AND2 C528 ( .A(a1stg_fdtos), .B(a1stg_in2[56]), .Z(N252) );
  GTECH_AND2 C529 ( .A(N254), .B(a1stg_in2[59]), .Z(N255) );
  GTECH_AND2 C530 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N254) );
  GTECH_AND2 C531 ( .A(a1stg_fstod), .B(a1stg_in2[59]), .Z(N257) );
  GTECH_AND2 C532 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[4]), .Z(N259) );
  GTECH_OR2 C533 ( .A(N274), .B(N275), .Z(a2stg_exp_in[3]) );
  GTECH_OR2 C534 ( .A(N272), .B(N273), .Z(N274) );
  GTECH_OR2 C535 ( .A(N269), .B(N271), .Z(N272) );
  GTECH_OR2 C536 ( .A(N267), .B(N268), .Z(N269) );
  GTECH_OR2 C537 ( .A(N264), .B(N266), .Z(N267) );
  GTECH_OR2 C538 ( .A(N261), .B(N263), .Z(N264) );
  GTECH_AND2 C539 ( .A(N260), .B(a1stg_in1a[55]), .Z(N261) );
  GTECH_AND2 C540 ( .A(a1stg_faddsubd), .B(N36), .Z(N260) );
  GTECH_AND2 C541 ( .A(N262), .B(a1stg_in1a[58]), .Z(N263) );
  GTECH_AND2 C542 ( .A(a1stg_faddsubs), .B(N36), .Z(N262) );
  GTECH_AND2 C543 ( .A(N265), .B(a1stg_in2[55]), .Z(N266) );
  GTECH_AND2 C544 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N265) );
  GTECH_AND2 C545 ( .A(a1stg_fdtos), .B(a1stg_in2[55]), .Z(N268) );
  GTECH_AND2 C546 ( .A(N270), .B(a1stg_in2[58]), .Z(N271) );
  GTECH_AND2 C547 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N270) );
  GTECH_AND2 C548 ( .A(a1stg_fstod), .B(a1stg_in2[58]), .Z(N273) );
  GTECH_AND2 C549 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[3]), .Z(N275) );
  GTECH_OR2 C550 ( .A(N290), .B(N291), .Z(a2stg_exp_in[2]) );
  GTECH_OR2 C551 ( .A(N288), .B(N289), .Z(N290) );
  GTECH_OR2 C552 ( .A(N285), .B(N287), .Z(N288) );
  GTECH_OR2 C553 ( .A(N283), .B(N284), .Z(N285) );
  GTECH_OR2 C554 ( .A(N280), .B(N282), .Z(N283) );
  GTECH_OR2 C555 ( .A(N277), .B(N279), .Z(N280) );
  GTECH_AND2 C556 ( .A(N276), .B(a1stg_in1a[54]), .Z(N277) );
  GTECH_AND2 C557 ( .A(a1stg_faddsubd), .B(N36), .Z(N276) );
  GTECH_AND2 C558 ( .A(N278), .B(a1stg_in1a[57]), .Z(N279) );
  GTECH_AND2 C559 ( .A(a1stg_faddsubs), .B(N36), .Z(N278) );
  GTECH_AND2 C560 ( .A(N281), .B(a1stg_in2[54]), .Z(N282) );
  GTECH_AND2 C561 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N281) );
  GTECH_AND2 C562 ( .A(a1stg_fdtos), .B(a1stg_in2[54]), .Z(N284) );
  GTECH_AND2 C563 ( .A(N286), .B(a1stg_in2[57]), .Z(N287) );
  GTECH_AND2 C564 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N286) );
  GTECH_AND2 C565 ( .A(a1stg_fstod), .B(a1stg_in2[57]), .Z(N289) );
  GTECH_AND2 C566 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[2]), .Z(N291) );
  GTECH_OR2 C567 ( .A(N306), .B(N307), .Z(a2stg_exp_in[1]) );
  GTECH_OR2 C568 ( .A(N304), .B(N305), .Z(N306) );
  GTECH_OR2 C569 ( .A(N301), .B(N303), .Z(N304) );
  GTECH_OR2 C570 ( .A(N299), .B(N300), .Z(N301) );
  GTECH_OR2 C571 ( .A(N296), .B(N298), .Z(N299) );
  GTECH_OR2 C572 ( .A(N293), .B(N295), .Z(N296) );
  GTECH_AND2 C573 ( .A(N292), .B(a1stg_in1a[53]), .Z(N293) );
  GTECH_AND2 C574 ( .A(a1stg_faddsubd), .B(N36), .Z(N292) );
  GTECH_AND2 C575 ( .A(N294), .B(a1stg_in1a[56]), .Z(N295) );
  GTECH_AND2 C576 ( .A(a1stg_faddsubs), .B(N36), .Z(N294) );
  GTECH_AND2 C577 ( .A(N297), .B(a1stg_in2[53]), .Z(N298) );
  GTECH_AND2 C578 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N297) );
  GTECH_AND2 C579 ( .A(a1stg_fdtos), .B(a1stg_in2[53]), .Z(N300) );
  GTECH_AND2 C580 ( .A(N302), .B(a1stg_in2[56]), .Z(N303) );
  GTECH_AND2 C581 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N302) );
  GTECH_AND2 C582 ( .A(a1stg_fstod), .B(a1stg_in2[56]), .Z(N305) );
  GTECH_AND2 C583 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[1]), .Z(N307) );
  GTECH_OR2 C584 ( .A(N322), .B(N323), .Z(a2stg_exp_in[0]) );
  GTECH_OR2 C585 ( .A(N320), .B(N321), .Z(N322) );
  GTECH_OR2 C586 ( .A(N317), .B(N319), .Z(N320) );
  GTECH_OR2 C587 ( .A(N315), .B(N316), .Z(N317) );
  GTECH_OR2 C588 ( .A(N312), .B(N314), .Z(N315) );
  GTECH_OR2 C589 ( .A(N309), .B(N311), .Z(N312) );
  GTECH_AND2 C590 ( .A(N308), .B(a1stg_in1a[52]), .Z(N309) );
  GTECH_AND2 C591 ( .A(a1stg_faddsubd), .B(N36), .Z(N308) );
  GTECH_AND2 C592 ( .A(N310), .B(a1stg_in1a[55]), .Z(N311) );
  GTECH_AND2 C593 ( .A(a1stg_faddsubs), .B(N36), .Z(N310) );
  GTECH_AND2 C594 ( .A(N313), .B(a1stg_in2[52]), .Z(N314) );
  GTECH_AND2 C595 ( .A(a1stg_faddsubd), .B(a1stg_expadd1[12]), .Z(N313) );
  GTECH_AND2 C596 ( .A(a1stg_fdtos), .B(a1stg_in2[52]), .Z(N316) );
  GTECH_AND2 C597 ( .A(N318), .B(a1stg_in2[55]), .Z(N319) );
  GTECH_AND2 C598 ( .A(a1stg_faddsubs), .B(a1stg_expadd1[12]), .Z(N318) );
  GTECH_AND2 C599 ( .A(a1stg_fstod), .B(a1stg_in2[55]), .Z(N321) );
  GTECH_AND2 C600 ( .A(a1stg_fsdtoix), .B(a1stg_expadd2_5_0[0]), .Z(N323) );
  GTECH_OR2 C601 ( .A(N326), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[12]) );
  GTECH_OR2 C602 ( .A(N325), .B(a1stg_fdtoi), .Z(N326) );
  GTECH_OR2 C603 ( .A(N324), .B(a1stg_fstox), .Z(N325) );
  GTECH_OR2 C604 ( .A(a1stg_fdtos), .B(a1stg_fstoi), .Z(N324) );
  GTECH_OR2 C605 ( .A(N329), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[11]) );
  GTECH_OR2 C606 ( .A(N328), .B(a1stg_fdtoi), .Z(N329) );
  GTECH_OR2 C607 ( .A(N327), .B(a1stg_fstox), .Z(N328) );
  GTECH_OR2 C608 ( .A(a1stg_fdtos), .B(a1stg_fstoi), .Z(N327) );
  GTECH_OR2 C609 ( .A(N330), .B(a1stg_fstox), .Z(a2stg_expadd_in2_in[10]) );
  GTECH_OR2 C610 ( .A(a1stg_fdtos), .B(a1stg_fstoi), .Z(N330) );
  GTECH_OR2 C611 ( .A(N333), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[9]) );
  GTECH_OR2 C612 ( .A(N332), .B(a1stg_fdtoi), .Z(N333) );
  GTECH_OR2 C613 ( .A(N331), .B(a1stg_fstox), .Z(N332) );
  GTECH_OR2 C614 ( .A(a1stg_fstod), .B(a1stg_fstoi), .Z(N331) );
  GTECH_OR2 C615 ( .A(N336), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[8]) );
  GTECH_OR2 C616 ( .A(N335), .B(a1stg_fdtoi), .Z(N336) );
  GTECH_OR2 C617 ( .A(N334), .B(a1stg_fstox), .Z(N335) );
  GTECH_OR2 C618 ( .A(a1stg_fstod), .B(a1stg_fstoi), .Z(N334) );
  GTECH_OR2 C619 ( .A(N337), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[7]) );
  GTECH_OR2 C620 ( .A(a1stg_fstod), .B(a1stg_fdtoi), .Z(N337) );
  GTECH_OR2 C621 ( .A(N340), .B(a1stg_fdtox), .Z(a2stg_expadd_in2_in[6]) );
  GTECH_OR2 C622 ( .A(N339), .B(a1stg_fdtoi), .Z(N340) );
  GTECH_OR2 C623 ( .A(N338), .B(a1stg_fstox), .Z(N339) );
  GTECH_OR2 C624 ( .A(a1stg_fdtos), .B(a1stg_fstoi), .Z(N338) );
  GTECH_OR2 C625 ( .A(N341), .B(a1stg_fdtoi), .Z(a2stg_expadd_in2_in[5]) );
  GTECH_OR2 C626 ( .A(a1stg_fdtos), .B(a1stg_fstoi), .Z(N341) );
  GTECH_OR2 C627 ( .A(N342), .B(N345), .Z(a3stg_exp_in[12]) );
  GTECH_AND2 C628 ( .A(a2stg_faddsubop), .B(a2stg_expa[12]), .Z(N342) );
  GTECH_AND2 C629 ( .A(a3stg_exp_add), .B(N344), .Z(N345) );
  GTECH_AND2 C630 ( .A(a2stg_expadd[12]), .B(N343), .Z(N344) );
  GTECH_NOT I_46 ( .A(a2stg_expadd[11]), .Z(N343) );
  GTECH_OR2 C632 ( .A(N346), .B(N348), .Z(a3stg_exp_in[11]) );
  GTECH_AND2 C633 ( .A(a2stg_faddsubop), .B(a2stg_expa[11]), .Z(N346) );
  GTECH_AND2 C634 ( .A(a3stg_exp_add), .B(N347), .Z(N348) );
  GTECH_AND2 C635 ( .A(a2stg_expadd[11]), .B(N343), .Z(N347) );
  GTECH_OR2 C637 ( .A(N352), .B(N354), .Z(a3stg_exp_in[10]) );
  GTECH_OR2 C638 ( .A(N351), .B(a3stg_exp_7ff), .Z(N352) );
  GTECH_OR2 C639 ( .A(N350), .B(a2stg_fxtod), .Z(N351) );
  GTECH_OR2 C640 ( .A(N349), .B(a2stg_fitod), .Z(N350) );
  GTECH_AND2 C641 ( .A(a2stg_faddsubop), .B(a2stg_expa[10]), .Z(N349) );
  GTECH_AND2 C642 ( .A(a3stg_exp_add), .B(N353), .Z(N354) );
  GTECH_AND2 C643 ( .A(a2stg_expadd[10]), .B(N343), .Z(N353) );
  GTECH_OR2 C645 ( .A(N356), .B(N358), .Z(a3stg_exp_in[9]) );
  GTECH_OR2 C646 ( .A(N355), .B(a3stg_exp_7ff), .Z(N356) );
  GTECH_AND2 C647 ( .A(a2stg_faddsubop), .B(a2stg_expa[9]), .Z(N355) );
  GTECH_AND2 C648 ( .A(a3stg_exp_add), .B(N357), .Z(N358) );
  GTECH_AND2 C649 ( .A(a2stg_expadd[9]), .B(N343), .Z(N357) );
  GTECH_OR2 C651 ( .A(N360), .B(N362), .Z(a3stg_exp_in[8]) );
  GTECH_OR2 C652 ( .A(N359), .B(a3stg_exp_7ff), .Z(N360) );
  GTECH_AND2 C653 ( .A(a2stg_faddsubop), .B(a2stg_expa[8]), .Z(N359) );
  GTECH_AND2 C654 ( .A(a3stg_exp_add), .B(N361), .Z(N362) );
  GTECH_AND2 C655 ( .A(a2stg_expadd[8]), .B(N343), .Z(N361) );
  GTECH_OR2 C657 ( .A(N367), .B(N369), .Z(a3stg_exp_in[7]) );
  GTECH_OR2 C658 ( .A(N366), .B(a3stg_exp_ff), .Z(N367) );
  GTECH_OR2 C659 ( .A(N365), .B(a3stg_exp_7ff), .Z(N366) );
  GTECH_OR2 C660 ( .A(N364), .B(a2stg_fxtos), .Z(N365) );
  GTECH_OR2 C661 ( .A(N363), .B(a2stg_fitos), .Z(N364) );
  GTECH_AND2 C662 ( .A(a2stg_faddsubop), .B(a2stg_expa[7]), .Z(N363) );
  GTECH_AND2 C663 ( .A(a3stg_exp_add), .B(N368), .Z(N369) );
  GTECH_AND2 C664 ( .A(a2stg_expadd[7]), .B(N343), .Z(N368) );
  GTECH_OR2 C666 ( .A(N372), .B(N374), .Z(a3stg_exp_in[6]) );
  GTECH_OR2 C667 ( .A(N371), .B(a3stg_exp_ff), .Z(N372) );
  GTECH_OR2 C668 ( .A(N370), .B(a3stg_exp_7ff), .Z(N371) );
  GTECH_AND2 C669 ( .A(a2stg_faddsubop), .B(a2stg_expa[6]), .Z(N370) );
  GTECH_AND2 C670 ( .A(a3stg_exp_add), .B(N373), .Z(N374) );
  GTECH_AND2 C671 ( .A(a2stg_expadd[6]), .B(N343), .Z(N373) );
  GTECH_OR2 C673 ( .A(N379), .B(N381), .Z(a3stg_exp_in[5]) );
  GTECH_OR2 C674 ( .A(N378), .B(a3stg_exp_ff), .Z(N379) );
  GTECH_OR2 C675 ( .A(N377), .B(a3stg_exp_7ff), .Z(N378) );
  GTECH_OR2 C676 ( .A(N376), .B(a2stg_fxtod), .Z(N377) );
  GTECH_OR2 C677 ( .A(N375), .B(a2stg_fxtos), .Z(N376) );
  GTECH_AND2 C678 ( .A(a2stg_faddsubop), .B(a2stg_expa[5]), .Z(N375) );
  GTECH_AND2 C679 ( .A(a3stg_exp_add), .B(N380), .Z(N381) );
  GTECH_AND2 C680 ( .A(a2stg_expadd[5]), .B(N343), .Z(N380) );
  GTECH_OR2 C682 ( .A(N388), .B(N390), .Z(a3stg_exp_in[4]) );
  GTECH_OR2 C683 ( .A(N387), .B(a3stg_exp_ff), .Z(N388) );
  GTECH_OR2 C684 ( .A(N386), .B(a3stg_exp_7ff), .Z(N387) );
  GTECH_OR2 C685 ( .A(N385), .B(a2stg_fxtod), .Z(N386) );
  GTECH_OR2 C686 ( .A(N384), .B(a2stg_fxtos), .Z(N385) );
  GTECH_OR2 C687 ( .A(N383), .B(a2stg_fitod), .Z(N384) );
  GTECH_OR2 C688 ( .A(N382), .B(a2stg_fitos), .Z(N383) );
  GTECH_AND2 C689 ( .A(a2stg_faddsubop), .B(a2stg_expa[4]), .Z(N382) );
  GTECH_AND2 C690 ( .A(a3stg_exp_add), .B(N389), .Z(N390) );
  GTECH_AND2 C691 ( .A(a2stg_expadd[4]), .B(N343), .Z(N389) );
  GTECH_OR2 C693 ( .A(N397), .B(N399), .Z(a3stg_exp_in[3]) );
  GTECH_OR2 C694 ( .A(N396), .B(a3stg_exp_ff), .Z(N397) );
  GTECH_OR2 C695 ( .A(N395), .B(a3stg_exp_7ff), .Z(N396) );
  GTECH_OR2 C696 ( .A(N394), .B(a2stg_fxtod), .Z(N395) );
  GTECH_OR2 C697 ( .A(N393), .B(a2stg_fxtos), .Z(N394) );
  GTECH_OR2 C698 ( .A(N392), .B(a2stg_fitod), .Z(N393) );
  GTECH_OR2 C699 ( .A(N391), .B(a2stg_fitos), .Z(N392) );
  GTECH_AND2 C700 ( .A(a2stg_faddsubop), .B(a2stg_expa[3]), .Z(N391) );
  GTECH_AND2 C701 ( .A(a3stg_exp_add), .B(N398), .Z(N399) );
  GTECH_AND2 C702 ( .A(a2stg_expadd[3]), .B(N343), .Z(N398) );
  GTECH_OR2 C704 ( .A(N406), .B(N408), .Z(a3stg_exp_in[2]) );
  GTECH_OR2 C705 ( .A(N405), .B(a3stg_exp_ff), .Z(N406) );
  GTECH_OR2 C706 ( .A(N404), .B(a3stg_exp_7ff), .Z(N405) );
  GTECH_OR2 C707 ( .A(N403), .B(a2stg_fxtod), .Z(N404) );
  GTECH_OR2 C708 ( .A(N402), .B(a2stg_fxtos), .Z(N403) );
  GTECH_OR2 C709 ( .A(N401), .B(a2stg_fitod), .Z(N402) );
  GTECH_OR2 C710 ( .A(N400), .B(a2stg_fitos), .Z(N401) );
  GTECH_AND2 C711 ( .A(a2stg_faddsubop), .B(a2stg_expa[2]), .Z(N400) );
  GTECH_AND2 C712 ( .A(a3stg_exp_add), .B(N407), .Z(N408) );
  GTECH_AND2 C713 ( .A(a2stg_expadd[2]), .B(N343), .Z(N407) );
  GTECH_OR2 C715 ( .A(N415), .B(N417), .Z(a3stg_exp_in[1]) );
  GTECH_OR2 C716 ( .A(N414), .B(a3stg_exp_ff), .Z(N415) );
  GTECH_OR2 C717 ( .A(N413), .B(a3stg_exp_7ff), .Z(N414) );
  GTECH_OR2 C718 ( .A(N412), .B(a2stg_fxtod), .Z(N413) );
  GTECH_OR2 C719 ( .A(N411), .B(a2stg_fxtos), .Z(N412) );
  GTECH_OR2 C720 ( .A(N410), .B(a2stg_fitod), .Z(N411) );
  GTECH_OR2 C721 ( .A(N409), .B(a2stg_fitos), .Z(N410) );
  GTECH_AND2 C722 ( .A(a2stg_faddsubop), .B(a2stg_expa[1]), .Z(N409) );
  GTECH_AND2 C723 ( .A(a3stg_exp_add), .B(N416), .Z(N417) );
  GTECH_AND2 C724 ( .A(a2stg_expadd[1]), .B(N343), .Z(N416) );
  GTECH_OR2 C726 ( .A(N420), .B(N422), .Z(a3stg_exp_in[0]) );
  GTECH_OR2 C727 ( .A(N419), .B(a3stg_exp_ff), .Z(N420) );
  GTECH_OR2 C728 ( .A(N418), .B(a3stg_exp_7ff), .Z(N419) );
  GTECH_AND2 C729 ( .A(a2stg_faddsubop), .B(a2stg_expa[0]), .Z(N418) );
  GTECH_AND2 C730 ( .A(a3stg_exp_add), .B(N421), .Z(N422) );
  GTECH_AND2 C731 ( .A(a2stg_expadd[0]), .B(N343), .Z(N421) );
  GTECH_AND2 C733 ( .A(N425), .B(a3stg_exp_plus1[12]), .Z(
        a4stg_exp_pre1_in[12]) );
  GTECH_AND2 C734 ( .A(N423), .B(N424), .Z(N425) );
  GTECH_AND2 C735 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N423) );
  GTECH_NOT I_47 ( .A(a3stg_inc_exp_inv), .Z(N424) );
  GTECH_AND2 C737 ( .A(N427), .B(a3stg_exp_plus1[11]), .Z(
        a4stg_exp_pre1_in[11]) );
  GTECH_AND2 C738 ( .A(N426), .B(N424), .Z(N427) );
  GTECH_AND2 C739 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N426) );
  GTECH_AND2 C741 ( .A(N429), .B(a3stg_exp_plus1[10]), .Z(
        a4stg_exp_pre1_in[10]) );
  GTECH_AND2 C742 ( .A(N428), .B(N424), .Z(N429) );
  GTECH_AND2 C743 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N428) );
  GTECH_AND2 C745 ( .A(N431), .B(a3stg_exp_plus1[9]), .Z(a4stg_exp_pre1_in[9])
         );
  GTECH_AND2 C746 ( .A(N430), .B(N424), .Z(N431) );
  GTECH_AND2 C747 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N430) );
  GTECH_AND2 C749 ( .A(N433), .B(a3stg_exp_plus1[8]), .Z(a4stg_exp_pre1_in[8])
         );
  GTECH_AND2 C750 ( .A(N432), .B(N424), .Z(N433) );
  GTECH_AND2 C751 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N432) );
  GTECH_AND2 C753 ( .A(N435), .B(a3stg_exp_plus1[7]), .Z(a4stg_exp_pre1_in[7])
         );
  GTECH_AND2 C754 ( .A(N434), .B(N424), .Z(N435) );
  GTECH_AND2 C755 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N434) );
  GTECH_AND2 C757 ( .A(N437), .B(a3stg_exp_plus1[6]), .Z(a4stg_exp_pre1_in[6])
         );
  GTECH_AND2 C758 ( .A(N436), .B(N424), .Z(N437) );
  GTECH_AND2 C759 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N436) );
  GTECH_AND2 C761 ( .A(N439), .B(a3stg_exp_plus1[5]), .Z(a4stg_exp_pre1_in[5])
         );
  GTECH_AND2 C762 ( .A(N438), .B(N424), .Z(N439) );
  GTECH_AND2 C763 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N438) );
  GTECH_AND2 C765 ( .A(N441), .B(a3stg_exp_plus1[4]), .Z(a4stg_exp_pre1_in[4])
         );
  GTECH_AND2 C766 ( .A(N440), .B(N424), .Z(N441) );
  GTECH_AND2 C767 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N440) );
  GTECH_AND2 C769 ( .A(N443), .B(a3stg_exp_plus1[3]), .Z(a4stg_exp_pre1_in[3])
         );
  GTECH_AND2 C770 ( .A(N442), .B(N424), .Z(N443) );
  GTECH_AND2 C771 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N442) );
  GTECH_AND2 C773 ( .A(N445), .B(a3stg_exp_plus1[2]), .Z(a4stg_exp_pre1_in[2])
         );
  GTECH_AND2 C774 ( .A(N444), .B(N424), .Z(N445) );
  GTECH_AND2 C775 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N444) );
  GTECH_AND2 C777 ( .A(N447), .B(a3stg_exp_plus1[1]), .Z(a4stg_exp_pre1_in[1])
         );
  GTECH_AND2 C778 ( .A(N446), .B(N424), .Z(N447) );
  GTECH_AND2 C779 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N446) );
  GTECH_AND2 C781 ( .A(N449), .B(a3stg_exp_plus1[0]), .Z(a4stg_exp_pre1_in[0])
         );
  GTECH_AND2 C782 ( .A(N448), .B(N424), .Z(N449) );
  GTECH_AND2 C783 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N448) );
  GTECH_AND2 C785 ( .A(N452), .B(a3stg_exp_minus1[12]), .Z(
        a4stg_exp_pre3_in[12]) );
  GTECH_AND2 C786 ( .A(N450), .B(N451), .Z(N452) );
  GTECH_AND2 C787 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N450) );
  GTECH_NOT I_48 ( .A(a3stg_dec_exp_inv), .Z(N451) );
  GTECH_AND2 C789 ( .A(N454), .B(a3stg_exp_minus1[11]), .Z(
        a4stg_exp_pre3_in[11]) );
  GTECH_AND2 C790 ( .A(N453), .B(N451), .Z(N454) );
  GTECH_AND2 C791 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N453) );
  GTECH_AND2 C793 ( .A(N456), .B(a3stg_exp_minus1[10]), .Z(
        a4stg_exp_pre3_in[10]) );
  GTECH_AND2 C794 ( .A(N455), .B(N451), .Z(N456) );
  GTECH_AND2 C795 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N455) );
  GTECH_AND2 C797 ( .A(N458), .B(a3stg_exp_minus1[9]), .Z(a4stg_exp_pre3_in[9]) );
  GTECH_AND2 C798 ( .A(N457), .B(N451), .Z(N458) );
  GTECH_AND2 C799 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N457) );
  GTECH_AND2 C801 ( .A(N460), .B(a3stg_exp_minus1[8]), .Z(a4stg_exp_pre3_in[8]) );
  GTECH_AND2 C802 ( .A(N459), .B(N451), .Z(N460) );
  GTECH_AND2 C803 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N459) );
  GTECH_AND2 C805 ( .A(N462), .B(a3stg_exp_minus1[7]), .Z(a4stg_exp_pre3_in[7]) );
  GTECH_AND2 C806 ( .A(N461), .B(N451), .Z(N462) );
  GTECH_AND2 C807 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N461) );
  GTECH_AND2 C809 ( .A(N464), .B(a3stg_exp_minus1[6]), .Z(a4stg_exp_pre3_in[6]) );
  GTECH_AND2 C810 ( .A(N463), .B(N451), .Z(N464) );
  GTECH_AND2 C811 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N463) );
  GTECH_AND2 C813 ( .A(N466), .B(a3stg_exp_minus1[5]), .Z(a4stg_exp_pre3_in[5]) );
  GTECH_AND2 C814 ( .A(N465), .B(N451), .Z(N466) );
  GTECH_AND2 C815 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N465) );
  GTECH_AND2 C817 ( .A(N468), .B(a3stg_exp_minus1[4]), .Z(a4stg_exp_pre3_in[4]) );
  GTECH_AND2 C818 ( .A(N467), .B(N451), .Z(N468) );
  GTECH_AND2 C819 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N467) );
  GTECH_AND2 C821 ( .A(N470), .B(a3stg_exp_minus1[3]), .Z(a4stg_exp_pre3_in[3]) );
  GTECH_AND2 C822 ( .A(N469), .B(N451), .Z(N470) );
  GTECH_AND2 C823 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N469) );
  GTECH_AND2 C825 ( .A(N472), .B(a3stg_exp_minus1[2]), .Z(a4stg_exp_pre3_in[2]) );
  GTECH_AND2 C826 ( .A(N471), .B(N451), .Z(N472) );
  GTECH_AND2 C827 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N471) );
  GTECH_AND2 C829 ( .A(N474), .B(a3stg_exp_minus1[1]), .Z(a4stg_exp_pre3_in[1]) );
  GTECH_AND2 C830 ( .A(N473), .B(N451), .Z(N474) );
  GTECH_AND2 C831 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N473) );
  GTECH_AND2 C833 ( .A(N476), .B(a3stg_exp_minus1[0]), .Z(a4stg_exp_pre3_in[0]) );
  GTECH_AND2 C834 ( .A(N475), .B(N451), .Z(N476) );
  GTECH_AND2 C835 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N475) );
  GTECH_OR2 C837 ( .A(N483), .B(N485), .Z(a4stg_exp_pre2_in[12]) );
  GTECH_OR2 C838 ( .A(N479), .B(N482), .Z(N483) );
  GTECH_AND2 C839 ( .A(N478), .B(a3stg_exp[12]), .Z(N479) );
  GTECH_AND2 C840 ( .A(N477), .B(a6stg_step), .Z(N478) );
  GTECH_NOT I_49 ( .A(a3stg_fdtos_inv), .Z(N477) );
  GTECH_AND2 C842 ( .A(N481), .B(a4stg_expshl[12]), .Z(N482) );
  GTECH_AND2 C843 ( .A(N480), .B(a6stg_step), .Z(N481) );
  GTECH_NOT I_50 ( .A(a4stg_fixtos_fxtod_inv), .Z(N480) );
  GTECH_AND2 C845 ( .A(N484), .B(a4stg_exp[12]), .Z(N485) );
  GTECH_NOT I_51 ( .A(a6stg_step), .Z(N484) );
  GTECH_OR2 C847 ( .A(N490), .B(N492), .Z(a4stg_exp_pre2_in[11]) );
  GTECH_OR2 C848 ( .A(N487), .B(N489), .Z(N490) );
  GTECH_AND2 C849 ( .A(N486), .B(a3stg_exp[11]), .Z(N487) );
  GTECH_AND2 C850 ( .A(N477), .B(a6stg_step), .Z(N486) );
  GTECH_AND2 C852 ( .A(N488), .B(a4stg_expshl[11]), .Z(N489) );
  GTECH_AND2 C853 ( .A(N480), .B(a6stg_step), .Z(N488) );
  GTECH_AND2 C855 ( .A(N491), .B(a4stg_exp_11_0[11]), .Z(N492) );
  GTECH_NOT I_52 ( .A(a6stg_step), .Z(N491) );
  GTECH_OR2 C857 ( .A(N497), .B(N499), .Z(a4stg_exp_pre2_in[10]) );
  GTECH_OR2 C858 ( .A(N494), .B(N496), .Z(N497) );
  GTECH_AND2 C859 ( .A(N493), .B(a3stg_exp_10_0[10]), .Z(N494) );
  GTECH_AND2 C860 ( .A(N477), .B(a6stg_step), .Z(N493) );
  GTECH_AND2 C862 ( .A(N495), .B(a4stg_expshl[10]), .Z(N496) );
  GTECH_AND2 C863 ( .A(N480), .B(a6stg_step), .Z(N495) );
  GTECH_AND2 C865 ( .A(N498), .B(a4stg_exp_11_0[10]), .Z(N499) );
  GTECH_NOT I_53 ( .A(a6stg_step), .Z(N498) );
  GTECH_OR2 C867 ( .A(N504), .B(N506), .Z(a4stg_exp_pre2_in[9]) );
  GTECH_OR2 C868 ( .A(N501), .B(N503), .Z(N504) );
  GTECH_AND2 C869 ( .A(N500), .B(a3stg_exp_10_0[9]), .Z(N501) );
  GTECH_AND2 C870 ( .A(N477), .B(a6stg_step), .Z(N500) );
  GTECH_AND2 C872 ( .A(N502), .B(a4stg_expshl[9]), .Z(N503) );
  GTECH_AND2 C873 ( .A(N480), .B(a6stg_step), .Z(N502) );
  GTECH_AND2 C875 ( .A(N505), .B(a4stg_exp_11_0[9]), .Z(N506) );
  GTECH_NOT I_54 ( .A(a6stg_step), .Z(N505) );
  GTECH_OR2 C877 ( .A(N511), .B(N513), .Z(a4stg_exp_pre2_in[8]) );
  GTECH_OR2 C878 ( .A(N508), .B(N510), .Z(N511) );
  GTECH_AND2 C879 ( .A(N507), .B(a3stg_exp_10_0[8]), .Z(N508) );
  GTECH_AND2 C880 ( .A(N477), .B(a6stg_step), .Z(N507) );
  GTECH_AND2 C882 ( .A(N509), .B(a4stg_expshl[8]), .Z(N510) );
  GTECH_AND2 C883 ( .A(N480), .B(a6stg_step), .Z(N509) );
  GTECH_AND2 C885 ( .A(N512), .B(a4stg_exp_11_0[8]), .Z(N513) );
  GTECH_NOT I_55 ( .A(a6stg_step), .Z(N512) );
  GTECH_OR2 C887 ( .A(N518), .B(N520), .Z(a4stg_exp_pre2_in[7]) );
  GTECH_OR2 C888 ( .A(N515), .B(N517), .Z(N518) );
  GTECH_AND2 C889 ( .A(N514), .B(a3stg_exp_10_0[7]), .Z(N515) );
  GTECH_AND2 C890 ( .A(N477), .B(a6stg_step), .Z(N514) );
  GTECH_AND2 C892 ( .A(N516), .B(a4stg_expshl[7]), .Z(N517) );
  GTECH_AND2 C893 ( .A(N480), .B(a6stg_step), .Z(N516) );
  GTECH_AND2 C895 ( .A(N519), .B(a4stg_exp_11_0[7]), .Z(N520) );
  GTECH_NOT I_56 ( .A(a6stg_step), .Z(N519) );
  GTECH_OR2 C897 ( .A(N525), .B(N527), .Z(a4stg_exp_pre2_in[6]) );
  GTECH_OR2 C898 ( .A(N522), .B(N524), .Z(N525) );
  GTECH_AND2 C899 ( .A(N521), .B(a3stg_exp_10_0[6]), .Z(N522) );
  GTECH_AND2 C900 ( .A(N477), .B(a6stg_step), .Z(N521) );
  GTECH_AND2 C902 ( .A(N523), .B(a4stg_expshl[6]), .Z(N524) );
  GTECH_AND2 C903 ( .A(N480), .B(a6stg_step), .Z(N523) );
  GTECH_AND2 C905 ( .A(N526), .B(a4stg_exp_11_0[6]), .Z(N527) );
  GTECH_NOT I_57 ( .A(a6stg_step), .Z(N526) );
  GTECH_OR2 C907 ( .A(N532), .B(N534), .Z(a4stg_exp_pre2_in[5]) );
  GTECH_OR2 C908 ( .A(N529), .B(N531), .Z(N532) );
  GTECH_AND2 C909 ( .A(N528), .B(a3stg_exp_10_0[5]), .Z(N529) );
  GTECH_AND2 C910 ( .A(N477), .B(a6stg_step), .Z(N528) );
  GTECH_AND2 C912 ( .A(N530), .B(a4stg_expshl[5]), .Z(N531) );
  GTECH_AND2 C913 ( .A(N480), .B(a6stg_step), .Z(N530) );
  GTECH_AND2 C915 ( .A(N533), .B(a4stg_exp_11_0[5]), .Z(N534) );
  GTECH_NOT I_58 ( .A(a6stg_step), .Z(N533) );
  GTECH_OR2 C917 ( .A(N539), .B(N541), .Z(a4stg_exp_pre2_in[4]) );
  GTECH_OR2 C918 ( .A(N536), .B(N538), .Z(N539) );
  GTECH_AND2 C919 ( .A(N535), .B(a3stg_exp_10_0[4]), .Z(N536) );
  GTECH_AND2 C920 ( .A(N477), .B(a6stg_step), .Z(N535) );
  GTECH_AND2 C922 ( .A(N537), .B(a4stg_expshl[4]), .Z(N538) );
  GTECH_AND2 C923 ( .A(N480), .B(a6stg_step), .Z(N537) );
  GTECH_AND2 C925 ( .A(N540), .B(a4stg_exp_11_0[4]), .Z(N541) );
  GTECH_NOT I_59 ( .A(a6stg_step), .Z(N540) );
  GTECH_OR2 C927 ( .A(N546), .B(N548), .Z(a4stg_exp_pre2_in[3]) );
  GTECH_OR2 C928 ( .A(N543), .B(N545), .Z(N546) );
  GTECH_AND2 C929 ( .A(N542), .B(a3stg_exp_10_0[3]), .Z(N543) );
  GTECH_AND2 C930 ( .A(N477), .B(a6stg_step), .Z(N542) );
  GTECH_AND2 C932 ( .A(N544), .B(a4stg_expshl[3]), .Z(N545) );
  GTECH_AND2 C933 ( .A(N480), .B(a6stg_step), .Z(N544) );
  GTECH_AND2 C935 ( .A(N547), .B(a4stg_exp_11_0[3]), .Z(N548) );
  GTECH_NOT I_60 ( .A(a6stg_step), .Z(N547) );
  GTECH_OR2 C937 ( .A(N553), .B(N555), .Z(a4stg_exp_pre2_in[2]) );
  GTECH_OR2 C938 ( .A(N550), .B(N552), .Z(N553) );
  GTECH_AND2 C939 ( .A(N549), .B(a3stg_exp_10_0[2]), .Z(N550) );
  GTECH_AND2 C940 ( .A(N477), .B(a6stg_step), .Z(N549) );
  GTECH_AND2 C942 ( .A(N551), .B(a4stg_expshl[2]), .Z(N552) );
  GTECH_AND2 C943 ( .A(N480), .B(a6stg_step), .Z(N551) );
  GTECH_AND2 C945 ( .A(N554), .B(a4stg_exp_11_0[2]), .Z(N555) );
  GTECH_NOT I_61 ( .A(a6stg_step), .Z(N554) );
  GTECH_OR2 C947 ( .A(N560), .B(N562), .Z(a4stg_exp_pre2_in[1]) );
  GTECH_OR2 C948 ( .A(N557), .B(N559), .Z(N560) );
  GTECH_AND2 C949 ( .A(N556), .B(a3stg_exp_10_0[1]), .Z(N557) );
  GTECH_AND2 C950 ( .A(N477), .B(a6stg_step), .Z(N556) );
  GTECH_AND2 C952 ( .A(N558), .B(a4stg_expshl[1]), .Z(N559) );
  GTECH_AND2 C953 ( .A(N480), .B(a6stg_step), .Z(N558) );
  GTECH_AND2 C955 ( .A(N561), .B(a4stg_exp_11_0[1]), .Z(N562) );
  GTECH_NOT I_62 ( .A(a6stg_step), .Z(N561) );
  GTECH_OR2 C957 ( .A(N567), .B(N569), .Z(a4stg_exp_pre2_in[0]) );
  GTECH_OR2 C958 ( .A(N564), .B(N566), .Z(N567) );
  GTECH_AND2 C959 ( .A(N563), .B(a3stg_exp_10_0[0]), .Z(N564) );
  GTECH_AND2 C960 ( .A(N477), .B(a6stg_step), .Z(N563) );
  GTECH_AND2 C962 ( .A(N565), .B(a4stg_expshl[0]), .Z(N566) );
  GTECH_AND2 C963 ( .A(N480), .B(a6stg_step), .Z(N565) );
  GTECH_AND2 C965 ( .A(N568), .B(a4stg_exp_11_0[0]), .Z(N569) );
  GTECH_NOT I_63 ( .A(a6stg_step), .Z(N568) );
  GTECH_AND2 C967 ( .A(N572), .B(a3stg_exp[12]), .Z(a4stg_exp_pre4_in[12]) );
  GTECH_AND2 C968 ( .A(N570), .B(N571), .Z(N572) );
  GTECH_AND2 C969 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N570) );
  GTECH_NOT I_64 ( .A(a3stg_same_exp_inv), .Z(N571) );
  GTECH_AND2 C971 ( .A(N574), .B(a3stg_exp[11]), .Z(a4stg_exp_pre4_in[11]) );
  GTECH_AND2 C972 ( .A(N573), .B(N571), .Z(N574) );
  GTECH_AND2 C973 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N573) );
  GTECH_AND2 C975 ( .A(N576), .B(a3stg_exp_10_0[10]), .Z(a4stg_exp_pre4_in[10]) );
  GTECH_AND2 C976 ( .A(N575), .B(N571), .Z(N576) );
  GTECH_AND2 C977 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N575) );
  GTECH_AND2 C979 ( .A(N578), .B(a3stg_exp_10_0[9]), .Z(a4stg_exp_pre4_in[9])
         );
  GTECH_AND2 C980 ( .A(N577), .B(N571), .Z(N578) );
  GTECH_AND2 C981 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N577) );
  GTECH_AND2 C983 ( .A(N580), .B(a3stg_exp_10_0[8]), .Z(a4stg_exp_pre4_in[8])
         );
  GTECH_AND2 C984 ( .A(N579), .B(N571), .Z(N580) );
  GTECH_AND2 C985 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N579) );
  GTECH_AND2 C987 ( .A(N582), .B(a3stg_exp_10_0[7]), .Z(a4stg_exp_pre4_in[7])
         );
  GTECH_AND2 C988 ( .A(N581), .B(N571), .Z(N582) );
  GTECH_AND2 C989 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N581) );
  GTECH_AND2 C991 ( .A(N584), .B(a3stg_exp_10_0[6]), .Z(a4stg_exp_pre4_in[6])
         );
  GTECH_AND2 C992 ( .A(N583), .B(N571), .Z(N584) );
  GTECH_AND2 C993 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N583) );
  GTECH_AND2 C995 ( .A(N586), .B(a3stg_exp_10_0[5]), .Z(a4stg_exp_pre4_in[5])
         );
  GTECH_AND2 C996 ( .A(N585), .B(N571), .Z(N586) );
  GTECH_AND2 C997 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N585) );
  GTECH_AND2 C999 ( .A(N588), .B(a3stg_exp_10_0[4]), .Z(a4stg_exp_pre4_in[4])
         );
  GTECH_AND2 C1000 ( .A(N587), .B(N571), .Z(N588) );
  GTECH_AND2 C1001 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N587) );
  GTECH_AND2 C1003 ( .A(N590), .B(a3stg_exp_10_0[3]), .Z(a4stg_exp_pre4_in[3])
         );
  GTECH_AND2 C1004 ( .A(N589), .B(N571), .Z(N590) );
  GTECH_AND2 C1005 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N589) );
  GTECH_AND2 C1007 ( .A(N592), .B(a3stg_exp_10_0[2]), .Z(a4stg_exp_pre4_in[2])
         );
  GTECH_AND2 C1008 ( .A(N591), .B(N571), .Z(N592) );
  GTECH_AND2 C1009 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N591) );
  GTECH_AND2 C1011 ( .A(N594), .B(a3stg_exp_10_0[1]), .Z(a4stg_exp_pre4_in[1])
         );
  GTECH_AND2 C1012 ( .A(N593), .B(N571), .Z(N594) );
  GTECH_AND2 C1013 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N593) );
  GTECH_AND2 C1015 ( .A(N596), .B(a3stg_exp_10_0[0]), .Z(a4stg_exp_pre4_in[0])
         );
  GTECH_AND2 C1016 ( .A(N595), .B(N571), .Z(N596) );
  GTECH_AND2 C1017 ( .A(a3stg_faddsubop), .B(a6stg_step), .Z(N595) );
  GTECH_OR2 C1019 ( .A(N598), .B(a4stg_exp_pre4[12]), .Z(a4stg_exp[12]) );
  GTECH_OR2 C1020 ( .A(N597), .B(a4stg_exp_pre3[12]), .Z(N598) );
  GTECH_OR2 C1021 ( .A(a4stg_exp_pre1[12]), .B(a4stg_exp_pre2[12]), .Z(N597)
         );
  GTECH_OR2 C1022 ( .A(N600), .B(a4stg_exp_pre4[11]), .Z(a4stg_exp_11_0[11])
         );
  GTECH_OR2 C1023 ( .A(N599), .B(a4stg_exp_pre3[11]), .Z(N600) );
  GTECH_OR2 C1024 ( .A(a4stg_exp_pre1[11]), .B(a4stg_exp_pre2[11]), .Z(N599)
         );
  GTECH_OR2 C1025 ( .A(N602), .B(a4stg_exp_pre4[10]), .Z(a4stg_exp_11_0[10])
         );
  GTECH_OR2 C1026 ( .A(N601), .B(a4stg_exp_pre3[10]), .Z(N602) );
  GTECH_OR2 C1027 ( .A(a4stg_exp_pre1[10]), .B(a4stg_exp_pre2[10]), .Z(N601)
         );
  GTECH_OR2 C1028 ( .A(N604), .B(a4stg_exp_pre4[9]), .Z(a4stg_exp_11_0[9]) );
  GTECH_OR2 C1029 ( .A(N603), .B(a4stg_exp_pre3[9]), .Z(N604) );
  GTECH_OR2 C1030 ( .A(a4stg_exp_pre1[9]), .B(a4stg_exp_pre2[9]), .Z(N603) );
  GTECH_OR2 C1031 ( .A(N606), .B(a4stg_exp_pre4[8]), .Z(a4stg_exp_11_0[8]) );
  GTECH_OR2 C1032 ( .A(N605), .B(a4stg_exp_pre3[8]), .Z(N606) );
  GTECH_OR2 C1033 ( .A(a4stg_exp_pre1[8]), .B(a4stg_exp_pre2[8]), .Z(N605) );
  GTECH_OR2 C1034 ( .A(N608), .B(a4stg_exp_pre4[7]), .Z(a4stg_exp_11_0[7]) );
  GTECH_OR2 C1035 ( .A(N607), .B(a4stg_exp_pre3[7]), .Z(N608) );
  GTECH_OR2 C1036 ( .A(a4stg_exp_pre1[7]), .B(a4stg_exp_pre2[7]), .Z(N607) );
  GTECH_OR2 C1037 ( .A(N610), .B(a4stg_exp_pre4[6]), .Z(a4stg_exp_11_0[6]) );
  GTECH_OR2 C1038 ( .A(N609), .B(a4stg_exp_pre3[6]), .Z(N610) );
  GTECH_OR2 C1039 ( .A(a4stg_exp_pre1[6]), .B(a4stg_exp_pre2[6]), .Z(N609) );
  GTECH_OR2 C1040 ( .A(N612), .B(a4stg_exp_pre4[5]), .Z(a4stg_exp_11_0[5]) );
  GTECH_OR2 C1041 ( .A(N611), .B(a4stg_exp_pre3[5]), .Z(N612) );
  GTECH_OR2 C1042 ( .A(a4stg_exp_pre1[5]), .B(a4stg_exp_pre2[5]), .Z(N611) );
  GTECH_OR2 C1043 ( .A(N614), .B(a4stg_exp_pre4[4]), .Z(a4stg_exp_11_0[4]) );
  GTECH_OR2 C1044 ( .A(N613), .B(a4stg_exp_pre3[4]), .Z(N614) );
  GTECH_OR2 C1045 ( .A(a4stg_exp_pre1[4]), .B(a4stg_exp_pre2[4]), .Z(N613) );
  GTECH_OR2 C1046 ( .A(N616), .B(a4stg_exp_pre4[3]), .Z(a4stg_exp_11_0[3]) );
  GTECH_OR2 C1047 ( .A(N615), .B(a4stg_exp_pre3[3]), .Z(N616) );
  GTECH_OR2 C1048 ( .A(a4stg_exp_pre1[3]), .B(a4stg_exp_pre2[3]), .Z(N615) );
  GTECH_OR2 C1049 ( .A(N618), .B(a4stg_exp_pre4[2]), .Z(a4stg_exp_11_0[2]) );
  GTECH_OR2 C1050 ( .A(N617), .B(a4stg_exp_pre3[2]), .Z(N618) );
  GTECH_OR2 C1051 ( .A(a4stg_exp_pre1[2]), .B(a4stg_exp_pre2[2]), .Z(N617) );
  GTECH_OR2 C1052 ( .A(N620), .B(a4stg_exp_pre4[1]), .Z(a4stg_exp_11_0[1]) );
  GTECH_OR2 C1053 ( .A(N619), .B(a4stg_exp_pre3[1]), .Z(N620) );
  GTECH_OR2 C1054 ( .A(a4stg_exp_pre1[1]), .B(a4stg_exp_pre2[1]), .Z(N619) );
  GTECH_OR2 C1055 ( .A(N622), .B(a4stg_exp_pre4[0]), .Z(a4stg_exp_11_0[0]) );
  GTECH_OR2 C1056 ( .A(N621), .B(a4stg_exp_pre3[0]), .Z(N622) );
  GTECH_OR2 C1057 ( .A(a4stg_exp_pre1[0]), .B(a4stg_exp_pre2[0]), .Z(N621) );
  GTECH_NOT I_65 ( .A(a4stg_shl_cnt[5]), .Z(a4stg_expadd_in2[5]) );
  GTECH_NOT I_66 ( .A(a4stg_shl_cnt[4]), .Z(a4stg_expadd_in2[4]) );
  GTECH_NOT I_67 ( .A(a4stg_shl_cnt[3]), .Z(a4stg_expadd_in2[3]) );
  GTECH_NOT I_68 ( .A(a4stg_shl_cnt[2]), .Z(a4stg_expadd_in2[2]) );
  GTECH_NOT I_69 ( .A(a4stg_shl_cnt[1]), .Z(a4stg_expadd_in2[1]) );
  GTECH_NOT I_70 ( .A(a4stg_shl_cnt[0]), .Z(a4stg_expadd_in2[0]) );
  GTECH_AND2 C1064 ( .A(a4stg_expadd[12]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[12]) );
  GTECH_AND2 C1065 ( .A(a4stg_expadd[11]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[11]) );
  GTECH_AND2 C1066 ( .A(a4stg_expadd[10]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[10]) );
  GTECH_AND2 C1067 ( .A(a4stg_expadd[9]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[9]) );
  GTECH_AND2 C1068 ( .A(a4stg_expadd[8]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[8]) );
  GTECH_AND2 C1069 ( .A(a4stg_expadd[7]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[7]) );
  GTECH_AND2 C1070 ( .A(a4stg_expadd[6]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[6]) );
  GTECH_AND2 C1071 ( .A(a4stg_expadd[5]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[5]) );
  GTECH_AND2 C1072 ( .A(a4stg_expadd[4]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[4]) );
  GTECH_AND2 C1073 ( .A(a4stg_expadd[3]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[3]) );
  GTECH_AND2 C1074 ( .A(a4stg_expadd[2]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[2]) );
  GTECH_AND2 C1075 ( .A(a4stg_expadd[1]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[1]) );
  GTECH_AND2 C1076 ( .A(a4stg_expadd[0]), .B(a4stg_denorm_inv), .Z(
        a4stg_expshl[0]) );
  GTECH_NOT I_71 ( .A(N627), .Z(add_exp_out_in1[10]) );
  GTECH_OR2 C1078 ( .A(N625), .B(N626), .Z(N627) );
  GTECH_OR2 C1079 ( .A(N623), .B(N624), .Z(N625) );
  GTECH_AND2 C1080 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[10]), .Z(N623) );
  GTECH_AND2 C1081 ( .A(a4stg_in_of), .B(a4stg_dblop), .Z(N624) );
  GTECH_AND2 C1082 ( .A(add_exp_out_expadd), .B(a4stg_expshl[10]), .Z(N626) );
  GTECH_NOT I_72 ( .A(N632), .Z(add_exp_out_in1[9]) );
  GTECH_OR2 C1084 ( .A(N630), .B(N631), .Z(N632) );
  GTECH_OR2 C1085 ( .A(N628), .B(N629), .Z(N630) );
  GTECH_AND2 C1086 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[9]), .Z(N628) );
  GTECH_AND2 C1087 ( .A(a4stg_in_of), .B(a4stg_dblop), .Z(N629) );
  GTECH_AND2 C1088 ( .A(add_exp_out_expadd), .B(a4stg_expshl[9]), .Z(N631) );
  GTECH_NOT I_73 ( .A(N637), .Z(add_exp_out_in1[8]) );
  GTECH_OR2 C1090 ( .A(N635), .B(N636), .Z(N637) );
  GTECH_OR2 C1091 ( .A(N633), .B(N634), .Z(N635) );
  GTECH_AND2 C1092 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[8]), .Z(N633) );
  GTECH_AND2 C1093 ( .A(a4stg_in_of), .B(a4stg_dblop), .Z(N634) );
  GTECH_AND2 C1094 ( .A(add_exp_out_expadd), .B(a4stg_expshl[8]), .Z(N636) );
  GTECH_NOT I_74 ( .A(N641), .Z(add_exp_out_in1[7]) );
  GTECH_OR2 C1096 ( .A(N639), .B(N640), .Z(N641) );
  GTECH_OR2 C1097 ( .A(N638), .B(a4stg_in_of), .Z(N639) );
  GTECH_AND2 C1098 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[7]), .Z(N638) );
  GTECH_AND2 C1099 ( .A(add_exp_out_expadd), .B(a4stg_expshl[7]), .Z(N640) );
  GTECH_NOT I_75 ( .A(N645), .Z(add_exp_out_in1[6]) );
  GTECH_OR2 C1101 ( .A(N643), .B(N644), .Z(N645) );
  GTECH_OR2 C1102 ( .A(N642), .B(a4stg_in_of), .Z(N643) );
  GTECH_AND2 C1103 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[6]), .Z(N642) );
  GTECH_AND2 C1104 ( .A(add_exp_out_expadd), .B(a4stg_expshl[6]), .Z(N644) );
  GTECH_NOT I_76 ( .A(N649), .Z(add_exp_out_in1[5]) );
  GTECH_OR2 C1106 ( .A(N647), .B(N648), .Z(N649) );
  GTECH_OR2 C1107 ( .A(N646), .B(a4stg_in_of), .Z(N647) );
  GTECH_AND2 C1108 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[5]), .Z(N646) );
  GTECH_AND2 C1109 ( .A(add_exp_out_expadd), .B(a4stg_expshl[5]), .Z(N648) );
  GTECH_NOT I_77 ( .A(N653), .Z(add_exp_out_in1[4]) );
  GTECH_OR2 C1111 ( .A(N651), .B(N652), .Z(N653) );
  GTECH_OR2 C1112 ( .A(N650), .B(a4stg_in_of), .Z(N651) );
  GTECH_AND2 C1113 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[4]), .Z(N650) );
  GTECH_AND2 C1114 ( .A(add_exp_out_expadd), .B(a4stg_expshl[4]), .Z(N652) );
  GTECH_NOT I_78 ( .A(N657), .Z(add_exp_out_in1[3]) );
  GTECH_OR2 C1116 ( .A(N655), .B(N656), .Z(N657) );
  GTECH_OR2 C1117 ( .A(N654), .B(a4stg_in_of), .Z(N655) );
  GTECH_AND2 C1118 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[3]), .Z(N654) );
  GTECH_AND2 C1119 ( .A(add_exp_out_expadd), .B(a4stg_expshl[3]), .Z(N656) );
  GTECH_NOT I_79 ( .A(N661), .Z(add_exp_out_in1[2]) );
  GTECH_OR2 C1121 ( .A(N659), .B(N660), .Z(N661) );
  GTECH_OR2 C1122 ( .A(N658), .B(a4stg_in_of), .Z(N659) );
  GTECH_AND2 C1123 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[2]), .Z(N658) );
  GTECH_AND2 C1124 ( .A(add_exp_out_expadd), .B(a4stg_expshl[2]), .Z(N660) );
  GTECH_NOT I_80 ( .A(N665), .Z(add_exp_out_in1[1]) );
  GTECH_OR2 C1126 ( .A(N663), .B(N664), .Z(N665) );
  GTECH_OR2 C1127 ( .A(N662), .B(a4stg_in_of), .Z(N663) );
  GTECH_AND2 C1128 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[1]), .Z(N662) );
  GTECH_AND2 C1129 ( .A(add_exp_out_expadd), .B(a4stg_expshl[1]), .Z(N664) );
  GTECH_NOT I_81 ( .A(N670), .Z(add_exp_out_in1[0]) );
  GTECH_OR2 C1131 ( .A(N668), .B(N669), .Z(N670) );
  GTECH_OR2 C1132 ( .A(N666), .B(N667), .Z(N668) );
  GTECH_AND2 C1133 ( .A(add_exp_out_exp1), .B(a4stg_exp_11_0[0]), .Z(N666) );
  GTECH_AND2 C1134 ( .A(a4stg_in_of), .B(a4stg_to_0_inv), .Z(N667) );
  GTECH_AND2 C1135 ( .A(add_exp_out_expadd), .B(a4stg_expshl[0]), .Z(N669) );
  GTECH_NOT I_82 ( .A(N672), .Z(add_exp_out_in2[10]) );
  GTECH_AND2 C1137 ( .A(N671), .B(a4stg_expinc[10]), .Z(N672) );
  GTECH_AND2 C1138 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N671)
         );
  GTECH_NOT I_83 ( .A(N674), .Z(add_exp_out_in2[9]) );
  GTECH_AND2 C1140 ( .A(N673), .B(a4stg_expinc[9]), .Z(N674) );
  GTECH_AND2 C1141 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N673)
         );
  GTECH_NOT I_84 ( .A(N676), .Z(add_exp_out_in2[8]) );
  GTECH_AND2 C1143 ( .A(N675), .B(a4stg_expinc[8]), .Z(N676) );
  GTECH_AND2 C1144 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N675)
         );
  GTECH_NOT I_85 ( .A(N678), .Z(add_exp_out_in2[7]) );
  GTECH_AND2 C1146 ( .A(N677), .B(a4stg_expinc[7]), .Z(N678) );
  GTECH_AND2 C1147 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N677)
         );
  GTECH_NOT I_86 ( .A(N680), .Z(add_exp_out_in2[6]) );
  GTECH_AND2 C1149 ( .A(N679), .B(a4stg_expinc[6]), .Z(N680) );
  GTECH_AND2 C1150 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N679)
         );
  GTECH_NOT I_87 ( .A(N682), .Z(add_exp_out_in2[5]) );
  GTECH_AND2 C1152 ( .A(N681), .B(a4stg_expinc[5]), .Z(N682) );
  GTECH_AND2 C1153 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N681)
         );
  GTECH_NOT I_88 ( .A(N684), .Z(add_exp_out_in2[4]) );
  GTECH_AND2 C1155 ( .A(N683), .B(a4stg_expinc[4]), .Z(N684) );
  GTECH_AND2 C1156 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N683)
         );
  GTECH_NOT I_89 ( .A(N686), .Z(add_exp_out_in2[3]) );
  GTECH_AND2 C1158 ( .A(N685), .B(a4stg_expinc[3]), .Z(N686) );
  GTECH_AND2 C1159 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N685)
         );
  GTECH_NOT I_90 ( .A(N688), .Z(add_exp_out_in2[2]) );
  GTECH_AND2 C1161 ( .A(N687), .B(a4stg_expinc[2]), .Z(N688) );
  GTECH_AND2 C1162 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N687)
         );
  GTECH_NOT I_91 ( .A(N690), .Z(add_exp_out_in2[1]) );
  GTECH_AND2 C1164 ( .A(N689), .B(a4stg_expinc[1]), .Z(N690) );
  GTECH_AND2 C1165 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N689)
         );
  GTECH_NOT I_92 ( .A(N692), .Z(add_exp_out_in2[0]) );
  GTECH_AND2 C1167 ( .A(N691), .B(a4stg_expinc[0]), .Z(N692) );
  GTECH_AND2 C1168 ( .A(add_exp_out_expinc), .B(a4stg_rndadd_cout), .Z(N691)
         );
  GTECH_NOT I_93 ( .A(N693), .Z(add_exp_out_in3[10]) );
  GTECH_AND2 C1170 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[10]), .Z(N693) );
  GTECH_NOT I_94 ( .A(N694), .Z(add_exp_out_in3[9]) );
  GTECH_AND2 C1172 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[9]), .Z(N694) );
  GTECH_NOT I_95 ( .A(N695), .Z(add_exp_out_in3[8]) );
  GTECH_AND2 C1174 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[8]), .Z(N695) );
  GTECH_NOT I_96 ( .A(N696), .Z(add_exp_out_in3[7]) );
  GTECH_AND2 C1176 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[7]), .Z(N696) );
  GTECH_NOT I_97 ( .A(N697), .Z(add_exp_out_in3[6]) );
  GTECH_AND2 C1178 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[6]), .Z(N697) );
  GTECH_NOT I_98 ( .A(N698), .Z(add_exp_out_in3[5]) );
  GTECH_AND2 C1180 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[5]), .Z(N698) );
  GTECH_NOT I_99 ( .A(N699), .Z(add_exp_out_in3[4]) );
  GTECH_AND2 C1182 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[4]), .Z(N699) );
  GTECH_NOT I_100 ( .A(N700), .Z(add_exp_out_in3[3]) );
  GTECH_AND2 C1184 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[3]), .Z(N700) );
  GTECH_NOT I_101 ( .A(N701), .Z(add_exp_out_in3[2]) );
  GTECH_AND2 C1186 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[2]), .Z(N701) );
  GTECH_NOT I_102 ( .A(N702), .Z(add_exp_out_in3[1]) );
  GTECH_AND2 C1188 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[1]), .Z(N702) );
  GTECH_NOT I_103 ( .A(N703), .Z(add_exp_out_in3[0]) );
  GTECH_AND2 C1190 ( .A(add_exp_out_exp), .B(a4stg_exp_11_0[0]), .Z(N703) );
  GTECH_NOT I_104 ( .A(N706), .Z(add_exp_out[10]) );
  GTECH_AND2 C1192 ( .A(N704), .B(N705), .Z(N706) );
  GTECH_AND2 C1193 ( .A(add_exp_out1[10]), .B(add_exp_out2[10]), .Z(N704) );
  GTECH_OR2 C1194 ( .A(add_exp_out3[10]), .B(add_exp_out4[10]), .Z(N705) );
  GTECH_NOT I_105 ( .A(N709), .Z(add_exp_out[9]) );
  GTECH_AND2 C1196 ( .A(N707), .B(N708), .Z(N709) );
  GTECH_AND2 C1197 ( .A(add_exp_out1[9]), .B(add_exp_out2[9]), .Z(N707) );
  GTECH_OR2 C1198 ( .A(add_exp_out3[9]), .B(add_exp_out4[9]), .Z(N708) );
  GTECH_NOT I_106 ( .A(N712), .Z(add_exp_out[8]) );
  GTECH_AND2 C1200 ( .A(N710), .B(N711), .Z(N712) );
  GTECH_AND2 C1201 ( .A(add_exp_out1[8]), .B(add_exp_out2[8]), .Z(N710) );
  GTECH_OR2 C1202 ( .A(add_exp_out3[8]), .B(add_exp_out4[8]), .Z(N711) );
  GTECH_NOT I_107 ( .A(N715), .Z(add_exp_out[7]) );
  GTECH_AND2 C1204 ( .A(N713), .B(N714), .Z(N715) );
  GTECH_AND2 C1205 ( .A(add_exp_out1[7]), .B(add_exp_out2[7]), .Z(N713) );
  GTECH_OR2 C1206 ( .A(add_exp_out3[7]), .B(add_exp_out4[7]), .Z(N714) );
  GTECH_NOT I_108 ( .A(N718), .Z(add_exp_out[6]) );
  GTECH_AND2 C1208 ( .A(N716), .B(N717), .Z(N718) );
  GTECH_AND2 C1209 ( .A(add_exp_out1[6]), .B(add_exp_out2[6]), .Z(N716) );
  GTECH_OR2 C1210 ( .A(add_exp_out3[6]), .B(add_exp_out4[6]), .Z(N717) );
  GTECH_NOT I_109 ( .A(N721), .Z(add_exp_out[5]) );
  GTECH_AND2 C1212 ( .A(N719), .B(N720), .Z(N721) );
  GTECH_AND2 C1213 ( .A(add_exp_out1[5]), .B(add_exp_out2[5]), .Z(N719) );
  GTECH_OR2 C1214 ( .A(add_exp_out3[5]), .B(add_exp_out4[5]), .Z(N720) );
  GTECH_NOT I_110 ( .A(N724), .Z(add_exp_out[4]) );
  GTECH_AND2 C1216 ( .A(N722), .B(N723), .Z(N724) );
  GTECH_AND2 C1217 ( .A(add_exp_out1[4]), .B(add_exp_out2[4]), .Z(N722) );
  GTECH_OR2 C1218 ( .A(add_exp_out3[4]), .B(add_exp_out4[4]), .Z(N723) );
  GTECH_NOT I_111 ( .A(N727), .Z(add_exp_out[3]) );
  GTECH_AND2 C1220 ( .A(N725), .B(N726), .Z(N727) );
  GTECH_AND2 C1221 ( .A(add_exp_out1[3]), .B(add_exp_out2[3]), .Z(N725) );
  GTECH_OR2 C1222 ( .A(add_exp_out3[3]), .B(add_exp_out4[3]), .Z(N726) );
  GTECH_NOT I_112 ( .A(N730), .Z(add_exp_out[2]) );
  GTECH_AND2 C1224 ( .A(N728), .B(N729), .Z(N730) );
  GTECH_AND2 C1225 ( .A(add_exp_out1[2]), .B(add_exp_out2[2]), .Z(N728) );
  GTECH_OR2 C1226 ( .A(add_exp_out3[2]), .B(add_exp_out4[2]), .Z(N729) );
  GTECH_NOT I_113 ( .A(N733), .Z(add_exp_out[1]) );
  GTECH_AND2 C1228 ( .A(N731), .B(N732), .Z(N733) );
  GTECH_AND2 C1229 ( .A(add_exp_out1[1]), .B(add_exp_out2[1]), .Z(N731) );
  GTECH_OR2 C1230 ( .A(add_exp_out3[1]), .B(add_exp_out4[1]), .Z(N732) );
  GTECH_NOT I_114 ( .A(N736), .Z(add_exp_out[0]) );
  GTECH_AND2 C1232 ( .A(N734), .B(N735), .Z(N736) );
  GTECH_AND2 C1233 ( .A(add_exp_out1[0]), .B(add_exp_out2[0]), .Z(N734) );
  GTECH_OR2 C1234 ( .A(add_exp_out3[0]), .B(add_exp_out4[0]), .Z(N735) );
endmodule


module dffe_SIZE63 ( din, en, clk, q, se, si, so );
  input [62:0] din;
  output [62:0] q;
  input [62:0] si;
  output [62:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68;
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N68) );
  SELECT_OP C267 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C275 ( .A(N3), .B(N2), .Z(N67) );
  GTECH_NOT I_2 ( .A(N67), .Z(N68) );
endmodule


module dffe_SIZE55 ( din, en, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60;
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N60) );
  SELECT_OP C235 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C243 ( .A(N3), .B(N2), .Z(N59) );
  GTECH_NOT I_2 ( .A(N59), .Z(N60) );
endmodule


module dffe_SIZE64 ( din, en, clk, q, se, si, so );
  input [63:0] din;
  output [63:0] q;
  input [63:0] si;
  output [63:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69;
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N69) );
  SELECT_OP C271 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C279 ( .A(N3), .B(N2), .Z(N68) );
  GTECH_NOT I_2 ( .A(N68), .Z(N69) );
endmodule


module fpu_in2_gt_in1_3b ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [2:0] din1;
  input [2:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14;
  wire   [2:0] din2_eq_din1;

  GTECH_NOT I_0 ( .A(N0), .Z(din2_eq_din1[2]) );
  GTECH_XOR2 C12 ( .A(din1[2]), .B(din2[2]), .Z(N0) );
  GTECH_NOT I_1 ( .A(N1), .Z(din2_eq_din1[1]) );
  GTECH_XOR2 C14 ( .A(din1[1]), .B(din2[1]), .Z(N1) );
  GTECH_NOT I_2 ( .A(N2), .Z(din2_eq_din1[0]) );
  GTECH_XOR2 C16 ( .A(din1[0]), .B(din2[0]), .Z(N2) );
  GTECH_NOT I_3 ( .A(N4), .Z(din2_neq_din1) );
  GTECH_AND2 C18 ( .A(N3), .B(din2_eq_din1[0]), .Z(N4) );
  GTECH_AND2 C19 ( .A(din2_eq_din1[2]), .B(din2_eq_din1[1]), .Z(N3) );
  GTECH_OR2 C20 ( .A(N10), .B(N14), .Z(din2_gt_din1) );
  GTECH_OR2 C21 ( .A(N6), .B(N9), .Z(N10) );
  GTECH_AND2 C22 ( .A(N5), .B(din2[2]), .Z(N6) );
  GTECH_NOT I_4 ( .A(din1[2]), .Z(N5) );
  GTECH_AND2 C24 ( .A(N8), .B(din2[1]), .Z(N9) );
  GTECH_AND2 C25 ( .A(din2_eq_din1[2]), .B(N7), .Z(N8) );
  GTECH_NOT I_5 ( .A(din1[1]), .Z(N7) );
  GTECH_AND2 C27 ( .A(N13), .B(din2[0]), .Z(N14) );
  GTECH_AND2 C28 ( .A(N11), .B(N12), .Z(N13) );
  GTECH_AND2 C29 ( .A(din2_eq_din1[2]), .B(din2_eq_din1[1]), .Z(N11) );
  GTECH_NOT I_6 ( .A(din1[0]), .Z(N12) );
endmodule


module fpu_in2_gt_in1_2b ( din1, din2, din2_neq_din1, din2_gt_din1 );
  input [1:0] din1;
  input [1:0] din2;
  output din2_neq_din1, din2_gt_din1;
  wire   N0, N1, N2, N3, N4, N5, N6, N7;
  wire   [1:0] din2_eq_din1;

  GTECH_NOT I_0 ( .A(N0), .Z(din2_eq_din1[1]) );
  GTECH_XOR2 C11 ( .A(din1[1]), .B(din2[1]), .Z(N0) );
  GTECH_NOT I_1 ( .A(N1), .Z(din2_eq_din1[0]) );
  GTECH_XOR2 C13 ( .A(din1[0]), .B(din2[0]), .Z(N1) );
  GTECH_NOT I_2 ( .A(N2), .Z(din2_neq_din1) );
  GTECH_AND2 C15 ( .A(din2_eq_din1[1]), .B(din2_eq_din1[0]), .Z(N2) );
  GTECH_OR2 C16 ( .A(N4), .B(N7), .Z(din2_gt_din1) );
  GTECH_AND2 C17 ( .A(N3), .B(din2[1]), .Z(N4) );
  GTECH_NOT I_3 ( .A(din1[1]), .Z(N3) );
  GTECH_AND2 C19 ( .A(N6), .B(din2[0]), .Z(N7) );
  GTECH_AND2 C20 ( .A(din2_eq_din1[1]), .B(N5), .Z(N6) );
  GTECH_NOT I_4 ( .A(din1[0]), .Z(N5) );
endmodule


module fpu_in2_gt_in1_3to1 ( din2_neq_din1_hi, din2_gt_din1_hi, 
        din2_neq_din1_mid, din2_gt_din1_mid, din2_neq_din1_lo, din2_gt_din1_lo, 
        din2_neq_din1, din2_gt_din1 );
  input din2_neq_din1_hi, din2_gt_din1_hi, din2_neq_din1_mid, din2_gt_din1_mid,
         din2_neq_din1_lo, din2_gt_din1_lo;
  output din2_neq_din1, din2_gt_din1;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8;

  GTECH_OR2 C9 ( .A(N1), .B(din2_neq_din1_lo), .Z(din2_neq_din1) );
  GTECH_OR2 C10 ( .A(din2_neq_din1_hi), .B(din2_neq_din1_mid), .Z(N1) );
  GTECH_NOT I_0 ( .A(din2_neq_din1_hi), .Z(N0) );
  GTECH_OR2 C12 ( .A(N5), .B(N8), .Z(din2_gt_din1) );
  GTECH_OR2 C13 ( .A(N2), .B(N4), .Z(N5) );
  GTECH_AND2 C14 ( .A(din2_neq_din1_hi), .B(din2_gt_din1_hi), .Z(N2) );
  GTECH_AND2 C15 ( .A(N3), .B(din2_gt_din1_mid), .Z(N4) );
  GTECH_AND2 C16 ( .A(N0), .B(din2_neq_din1_mid), .Z(N3) );
  GTECH_AND2 C17 ( .A(N7), .B(din2_gt_din1_lo), .Z(N8) );
  GTECH_AND2 C18 ( .A(N0), .B(N6), .Z(N7) );
  GTECH_NOT I_1 ( .A(din2_neq_din1_mid), .Z(N6) );
endmodule


module fpu_in2_gt_in1_frac ( din1, din2, sngop, expadd11, expeq, din2_neq_din1, 
        din2_gt_din1, din2_gt1_din1 );
  input [54:0] din1;
  input [54:0] din2;
  input sngop, expadd11, expeq;
  output din2_neq_din1, din2_gt_din1, din2_gt1_din1;
  wire   din2_neq_din1_54_52, din2_gt_din1_54_52, din2_neq_din1_51_50,
         din2_gt_din1_51_50, din2_neq_din1_49_48, din2_gt_din1_49_48,
         din2_neq_din1_47_45, din2_gt_din1_47_45, din2_neq_din1_44_42,
         din2_gt_din1_44_42, din2_neq_din1_41_39, din2_gt_din1_41_39,
         din2_neq_din1_38_36, din2_gt_din1_38_36, din2_neq_din1_35_33,
         din2_gt_din1_35_33, din2_neq_din1_32_30, din2_gt_din1_32_30,
         din2_neq_din1_29_27, din2_gt_din1_29_27, din2_neq_din1_26_24,
         din2_gt_din1_26_24, din2_neq_din1_23_21, din2_gt_din1_23_21,
         din2_neq_din1_20_18, din2_gt_din1_20_18, din2_neq_din1_17_15,
         din2_gt_din1_17_15, din2_neq_din1_14_12, din2_gt_din1_14_12,
         din2_neq_din1_11_9, din2_gt_din1_11_9, din2_neq_din1_8_6,
         din2_gt_din1_8_6, din2_neq_din1_5_3, din2_gt_din1_5_3,
         din2_neq_din1_2_0, din2_gt_din1_2_0, din2_neq_din1_51_45,
         din2_gt_din1_51_45, din2_neq_din1_44_36, din2_gt_din1_44_36,
         din2_neq_din1_35_27, din2_gt_din1_35_27, din2_neq_din1_26_18,
         din2_gt_din1_26_18, din2_neq_din1_17_9, din2_gt_din1_17_9,
         din2_neq_din1_8_0, din2_gt_din1_8_0, din2_neq_din1_51_27,
         din2_gt_din1_51_27, din2_neq_din1_26_0, din2_gt_din1_26_0, N0, N1, N2,
         N3, N4, N5, N6, N7, N8, N9, N10, N11, N12;

  fpu_in2_gt_in1_3b fpu_in2_gt_in1_54_52 ( .din1(din1[54:52]), .din2(
        din2[54:52]), .din2_neq_din1(din2_neq_din1_54_52), .din2_gt_din1(
        din2_gt_din1_54_52) );
  fpu_in2_gt_in1_2b fpu_in2_gt_in1_51_50 ( .din1(din1[51:50]), .din2(
        din2[51:50]), .din2_neq_din1(din2_neq_din1_51_50), .din2_gt_din1(
        din2_gt_din1_51_50) );
  fpu_in2_gt_in1_2b fpu_in2_gt_in1_49_48 ( .din1(din1[49:48]), .din2(
        din2[49:48]), .din2_neq_din1(din2_neq_din1_49_48), .din2_gt_din1(
        din2_gt_din1_49_48) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_47_45 ( .din1(din1[47:45]), .din2(
        din2[47:45]), .din2_neq_din1(din2_neq_din1_47_45), .din2_gt_din1(
        din2_gt_din1_47_45) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_44_42 ( .din1(din1[44:42]), .din2(
        din2[44:42]), .din2_neq_din1(din2_neq_din1_44_42), .din2_gt_din1(
        din2_gt_din1_44_42) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_41_39 ( .din1(din1[41:39]), .din2(
        din2[41:39]), .din2_neq_din1(din2_neq_din1_41_39), .din2_gt_din1(
        din2_gt_din1_41_39) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_38_36 ( .din1(din1[38:36]), .din2(
        din2[38:36]), .din2_neq_din1(din2_neq_din1_38_36), .din2_gt_din1(
        din2_gt_din1_38_36) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_35_33 ( .din1(din1[35:33]), .din2(
        din2[35:33]), .din2_neq_din1(din2_neq_din1_35_33), .din2_gt_din1(
        din2_gt_din1_35_33) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_32_30 ( .din1(din1[32:30]), .din2(
        din2[32:30]), .din2_neq_din1(din2_neq_din1_32_30), .din2_gt_din1(
        din2_gt_din1_32_30) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_29_27 ( .din1(din1[29:27]), .din2(
        din2[29:27]), .din2_neq_din1(din2_neq_din1_29_27), .din2_gt_din1(
        din2_gt_din1_29_27) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_26_24 ( .din1(din1[26:24]), .din2(
        din2[26:24]), .din2_neq_din1(din2_neq_din1_26_24), .din2_gt_din1(
        din2_gt_din1_26_24) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_23_21 ( .din1(din1[23:21]), .din2(
        din2[23:21]), .din2_neq_din1(din2_neq_din1_23_21), .din2_gt_din1(
        din2_gt_din1_23_21) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_20_18 ( .din1(din1[20:18]), .din2(
        din2[20:18]), .din2_neq_din1(din2_neq_din1_20_18), .din2_gt_din1(
        din2_gt_din1_20_18) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_17_15 ( .din1(din1[17:15]), .din2(
        din2[17:15]), .din2_neq_din1(din2_neq_din1_17_15), .din2_gt_din1(
        din2_gt_din1_17_15) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_14_12 ( .din1(din1[14:12]), .din2(
        din2[14:12]), .din2_neq_din1(din2_neq_din1_14_12), .din2_gt_din1(
        din2_gt_din1_14_12) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_11_9 ( .din1(din1[11:9]), .din2(din2[11:9]), 
        .din2_neq_din1(din2_neq_din1_11_9), .din2_gt_din1(din2_gt_din1_11_9)
         );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_8_6 ( .din1(din1[8:6]), .din2(din2[8:6]), 
        .din2_neq_din1(din2_neq_din1_8_6), .din2_gt_din1(din2_gt_din1_8_6) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_5_3 ( .din1(din1[5:3]), .din2(din2[5:3]), 
        .din2_neq_din1(din2_neq_din1_5_3), .din2_gt_din1(din2_gt_din1_5_3) );
  fpu_in2_gt_in1_3b fpu_in2_gt_in1_2_0 ( .din1(din1[2:0]), .din2(din2[2:0]), 
        .din2_neq_din1(din2_neq_din1_2_0), .din2_gt_din1(din2_gt_din1_2_0) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_51_45 ( .din2_neq_din1_hi(
        din2_neq_din1_51_50), .din2_gt_din1_hi(din2_gt_din1_51_50), 
        .din2_neq_din1_mid(din2_neq_din1_49_48), .din2_gt_din1_mid(
        din2_gt_din1_49_48), .din2_neq_din1_lo(din2_neq_din1_47_45), 
        .din2_gt_din1_lo(din2_gt_din1_47_45), .din2_neq_din1(
        din2_neq_din1_51_45), .din2_gt_din1(din2_gt_din1_51_45) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_44_36 ( .din2_neq_din1_hi(
        din2_neq_din1_44_42), .din2_gt_din1_hi(din2_gt_din1_44_42), 
        .din2_neq_din1_mid(din2_neq_din1_41_39), .din2_gt_din1_mid(
        din2_gt_din1_41_39), .din2_neq_din1_lo(din2_neq_din1_38_36), 
        .din2_gt_din1_lo(din2_gt_din1_38_36), .din2_neq_din1(
        din2_neq_din1_44_36), .din2_gt_din1(din2_gt_din1_44_36) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_35_27 ( .din2_neq_din1_hi(
        din2_neq_din1_35_33), .din2_gt_din1_hi(din2_gt_din1_35_33), 
        .din2_neq_din1_mid(din2_neq_din1_32_30), .din2_gt_din1_mid(
        din2_gt_din1_32_30), .din2_neq_din1_lo(din2_neq_din1_29_27), 
        .din2_gt_din1_lo(din2_gt_din1_29_27), .din2_neq_din1(
        din2_neq_din1_35_27), .din2_gt_din1(din2_gt_din1_35_27) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_26_18 ( .din2_neq_din1_hi(
        din2_neq_din1_26_24), .din2_gt_din1_hi(din2_gt_din1_26_24), 
        .din2_neq_din1_mid(din2_neq_din1_23_21), .din2_gt_din1_mid(
        din2_gt_din1_23_21), .din2_neq_din1_lo(din2_neq_din1_20_18), 
        .din2_gt_din1_lo(din2_gt_din1_20_18), .din2_neq_din1(
        din2_neq_din1_26_18), .din2_gt_din1(din2_gt_din1_26_18) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_17_9 ( .din2_neq_din1_hi(
        din2_neq_din1_17_15), .din2_gt_din1_hi(din2_gt_din1_17_15), 
        .din2_neq_din1_mid(din2_neq_din1_14_12), .din2_gt_din1_mid(
        din2_gt_din1_14_12), .din2_neq_din1_lo(din2_neq_din1_11_9), 
        .din2_gt_din1_lo(din2_gt_din1_11_9), .din2_neq_din1(din2_neq_din1_17_9), .din2_gt_din1(din2_gt_din1_17_9) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_8_0 ( .din2_neq_din1_hi(din2_neq_din1_8_6), .din2_gt_din1_hi(din2_gt_din1_8_6), .din2_neq_din1_mid(din2_neq_din1_5_3), 
        .din2_gt_din1_mid(din2_gt_din1_5_3), .din2_neq_din1_lo(
        din2_neq_din1_2_0), .din2_gt_din1_lo(din2_gt_din1_2_0), 
        .din2_neq_din1(din2_neq_din1_8_0), .din2_gt_din1(din2_gt_din1_8_0) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_51_27 ( .din2_neq_din1_hi(
        din2_neq_din1_51_45), .din2_gt_din1_hi(din2_gt_din1_51_45), 
        .din2_neq_din1_mid(din2_neq_din1_44_36), .din2_gt_din1_mid(
        din2_gt_din1_44_36), .din2_neq_din1_lo(din2_neq_din1_35_27), 
        .din2_gt_din1_lo(din2_gt_din1_35_27), .din2_neq_din1(
        din2_neq_din1_51_27), .din2_gt_din1(din2_gt_din1_51_27) );
  fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_26_0 ( .din2_neq_din1_hi(
        din2_neq_din1_26_18), .din2_gt_din1_hi(din2_gt_din1_26_18), 
        .din2_neq_din1_mid(din2_neq_din1_17_9), .din2_gt_din1_mid(
        din2_gt_din1_17_9), .din2_neq_din1_lo(din2_neq_din1_8_0), 
        .din2_gt_din1_lo(din2_gt_din1_8_0), .din2_neq_din1(din2_neq_din1_26_0), 
        .din2_gt_din1(din2_gt_din1_26_0) );
  GTECH_OR2 C10 ( .A(N1), .B(N2), .Z(din2_neq_din1) );
  GTECH_OR2 C11 ( .A(din2_neq_din1_51_27), .B(din2_neq_din1_26_0), .Z(N1) );
  GTECH_AND2 C12 ( .A(din2_neq_din1_54_52), .B(sngop), .Z(N2) );
  GTECH_NOT I_0 ( .A(N3), .Z(N0) );
  GTECH_AND2 C14 ( .A(din2_neq_din1_54_52), .B(sngop), .Z(N3) );
  GTECH_OR2 C15 ( .A(N8), .B(N11), .Z(din2_gt_din1) );
  GTECH_OR2 C16 ( .A(N5), .B(N7), .Z(N8) );
  GTECH_AND2 C17 ( .A(N4), .B(sngop), .Z(N5) );
  GTECH_AND2 C18 ( .A(din2_neq_din1_54_52), .B(din2_gt_din1_54_52), .Z(N4) );
  GTECH_AND2 C19 ( .A(N6), .B(din2_gt_din1_51_27), .Z(N7) );
  GTECH_AND2 C20 ( .A(N0), .B(din2_neq_din1_51_27), .Z(N6) );
  GTECH_AND2 C21 ( .A(N10), .B(din2_gt_din1_26_0), .Z(N11) );
  GTECH_AND2 C22 ( .A(N0), .B(N9), .Z(N10) );
  GTECH_NOT I_1 ( .A(din2_neq_din1_51_27), .Z(N9) );
  GTECH_OR2 C24 ( .A(expadd11), .B(N12), .Z(din2_gt1_din1) );
  GTECH_AND2 C25 ( .A(din2_gt_din1), .B(expeq), .Z(N12) );
endmodule


module dffe_SIZE54 ( din, en, clk, q, se, si, so );
  input [53:0] din;
  output [53:0] q;
  input [53:0] si;
  output [53:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59;
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N59) );
  SELECT_OP C231 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C239 ( .A(N3), .B(N2), .Z(N58) );
  GTECH_NOT I_2 ( .A(N58), .Z(N59) );
endmodule


module fpu_denorm_3b ( din1, din2, din2_din1_nz, din2_din1_denorm );
  input [2:0] din1;
  input [2:0] din2;
  output din2_din1_nz, din2_din1_denorm;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8;
  wire   [2:0] din2_din1_zero;

  GTECH_NOT I_0 ( .A(N0), .Z(din2_din1_zero[2]) );
  GTECH_OR2 C12 ( .A(din1[2]), .B(din2[2]), .Z(N0) );
  GTECH_NOT I_1 ( .A(N1), .Z(din2_din1_zero[1]) );
  GTECH_OR2 C14 ( .A(din1[1]), .B(din2[1]), .Z(N1) );
  GTECH_NOT I_2 ( .A(N2), .Z(din2_din1_zero[0]) );
  GTECH_OR2 C16 ( .A(din1[0]), .B(din2[0]), .Z(N2) );
  GTECH_NOT I_3 ( .A(N4), .Z(din2_din1_nz) );
  GTECH_AND2 C18 ( .A(N3), .B(din2_din1_zero[0]), .Z(N4) );
  GTECH_AND2 C19 ( .A(din2_din1_zero[2]), .B(din2_din1_zero[1]), .Z(N3) );
  GTECH_OR2 C20 ( .A(N6), .B(N8), .Z(din2_din1_denorm) );
  GTECH_OR2 C21 ( .A(din2[2]), .B(N5), .Z(N6) );
  GTECH_AND2 C22 ( .A(din2_din1_zero[2]), .B(din2[1]), .Z(N5) );
  GTECH_AND2 C23 ( .A(N7), .B(din2[0]), .Z(N8) );
  GTECH_AND2 C24 ( .A(din2_din1_zero[2]), .B(din2_din1_zero[1]), .Z(N7) );
endmodule


module fpu_denorm_3to1 ( din2_din1_nz_hi, din2_din1_denorm_hi, 
        din2_din1_nz_mid, din2_din1_denorm_mid, din2_din1_nz_lo, 
        din2_din1_denorm_lo, din2_din1_nz, din2_din1_denorm );
  input din2_din1_nz_hi, din2_din1_denorm_hi, din2_din1_nz_mid,
         din2_din1_denorm_mid, din2_din1_nz_lo, din2_din1_denorm_lo;
  output din2_din1_nz, din2_din1_denorm;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8;

  GTECH_OR2 C9 ( .A(N1), .B(din2_din1_nz_lo), .Z(din2_din1_nz) );
  GTECH_OR2 C10 ( .A(din2_din1_nz_hi), .B(din2_din1_nz_mid), .Z(N1) );
  GTECH_NOT I_0 ( .A(din2_din1_nz_hi), .Z(N0) );
  GTECH_OR2 C12 ( .A(N5), .B(N8), .Z(din2_din1_denorm) );
  GTECH_OR2 C13 ( .A(N2), .B(N4), .Z(N5) );
  GTECH_AND2 C14 ( .A(din2_din1_nz_hi), .B(din2_din1_denorm_hi), .Z(N2) );
  GTECH_AND2 C15 ( .A(N3), .B(din2_din1_denorm_mid), .Z(N4) );
  GTECH_AND2 C16 ( .A(N0), .B(din2_din1_nz_mid), .Z(N3) );
  GTECH_AND2 C17 ( .A(N7), .B(din2_din1_denorm_lo), .Z(N8) );
  GTECH_AND2 C18 ( .A(N0), .B(N6), .Z(N7) );
  GTECH_NOT I_1 ( .A(din2_din1_nz_mid), .Z(N6) );
endmodule


module fpu_denorm_frac ( din1, din2, din2_din1_denorm, din2_din1_denorm_inv, 
        din2_din1_denorma, din2_din1_denorm_inva );
  input [53:0] din1;
  input [53:0] din2;
  output din2_din1_denorm, din2_din1_denorm_inv, din2_din1_denorma,
         din2_din1_denorm_inva;
  wire   din2_din1_denorm, din2_din1_denorm_inv, din2_din1_nz_53_51,
         din2_din1_denorm_53_51, din2_din1_nz_50_48, din2_din1_denorm_50_48,
         din2_din1_nz_47_45, din2_din1_denorm_47_45, din2_din1_nz_44_42,
         din2_din1_denorm_44_42, din2_din1_nz_41_39, din2_din1_denorm_41_39,
         din2_din1_nz_38_36, din2_din1_denorm_38_36, din2_din1_nz_35_33,
         din2_din1_denorm_35_33, din2_din1_nz_32_30, din2_din1_denorm_32_30,
         din2_din1_nz_29_27, din2_din1_denorm_29_27, din2_din1_nz_26_24,
         din2_din1_denorm_26_24, din2_din1_nz_23_21, din2_din1_denorm_23_21,
         din2_din1_nz_20_18, din2_din1_denorm_20_18, din2_din1_nz_17_15,
         din2_din1_denorm_17_15, din2_din1_nz_14_12, din2_din1_denorm_14_12,
         din2_din1_nz_11_9, din2_din1_denorm_11_9, din2_din1_nz_8_6,
         din2_din1_denorm_8_6, din2_din1_nz_5_3, din2_din1_denorm_5_3,
         din2_din1_nz_2_0, din2_din1_denorm_2_0, din2_din1_nz_53_45,
         din2_din1_denorm_53_45, din2_din1_nz_44_36, din2_din1_denorm_44_36,
         din2_din1_nz_35_27, din2_din1_denorm_35_27, din2_din1_nz_26_18,
         din2_din1_denorm_26_18, din2_din1_nz_17_9, din2_din1_denorm_17_9,
         din2_din1_nz_8_0, din2_din1_denorm_8_0, din2_din1_nz_53_27,
         din2_din1_denorm_53_27, din2_din1_nz_26_0, din2_din1_denorm_26_0, N0,
         N1, N2, N3, N4, N5;
  assign din2_din1_denorma = din2_din1_denorm;
  assign din2_din1_denorm_inva = din2_din1_denorm_inv;

  fpu_denorm_3b i_fpu_denorm_53_51 ( .din1(din1[53:51]), .din2(din2[53:51]), 
        .din2_din1_nz(din2_din1_nz_53_51), .din2_din1_denorm(
        din2_din1_denorm_53_51) );
  fpu_denorm_3b i_fpu_denorm_50_48 ( .din1(din1[50:48]), .din2(din2[50:48]), 
        .din2_din1_nz(din2_din1_nz_50_48), .din2_din1_denorm(
        din2_din1_denorm_50_48) );
  fpu_denorm_3b i_fpu_denorm_47_45 ( .din1(din1[47:45]), .din2(din2[47:45]), 
        .din2_din1_nz(din2_din1_nz_47_45), .din2_din1_denorm(
        din2_din1_denorm_47_45) );
  fpu_denorm_3b i_fpu_denorm_44_42 ( .din1(din1[44:42]), .din2(din2[44:42]), 
        .din2_din1_nz(din2_din1_nz_44_42), .din2_din1_denorm(
        din2_din1_denorm_44_42) );
  fpu_denorm_3b i_fpu_denorm_41_39 ( .din1(din1[41:39]), .din2(din2[41:39]), 
        .din2_din1_nz(din2_din1_nz_41_39), .din2_din1_denorm(
        din2_din1_denorm_41_39) );
  fpu_denorm_3b i_fpu_denorm_38_36 ( .din1(din1[38:36]), .din2(din2[38:36]), 
        .din2_din1_nz(din2_din1_nz_38_36), .din2_din1_denorm(
        din2_din1_denorm_38_36) );
  fpu_denorm_3b i_fpu_denorm_35_33 ( .din1(din1[35:33]), .din2(din2[35:33]), 
        .din2_din1_nz(din2_din1_nz_35_33), .din2_din1_denorm(
        din2_din1_denorm_35_33) );
  fpu_denorm_3b i_fpu_denorm_32_30 ( .din1(din1[32:30]), .din2(din2[32:30]), 
        .din2_din1_nz(din2_din1_nz_32_30), .din2_din1_denorm(
        din2_din1_denorm_32_30) );
  fpu_denorm_3b i_fpu_denorm_29_27 ( .din1(din1[29:27]), .din2(din2[29:27]), 
        .din2_din1_nz(din2_din1_nz_29_27), .din2_din1_denorm(
        din2_din1_denorm_29_27) );
  fpu_denorm_3b i_fpu_denorm_26_24 ( .din1(din1[26:24]), .din2(din2[26:24]), 
        .din2_din1_nz(din2_din1_nz_26_24), .din2_din1_denorm(
        din2_din1_denorm_26_24) );
  fpu_denorm_3b i_fpu_denorm_23_21 ( .din1(din1[23:21]), .din2(din2[23:21]), 
        .din2_din1_nz(din2_din1_nz_23_21), .din2_din1_denorm(
        din2_din1_denorm_23_21) );
  fpu_denorm_3b i_fpu_denorm_20_18 ( .din1(din1[20:18]), .din2(din2[20:18]), 
        .din2_din1_nz(din2_din1_nz_20_18), .din2_din1_denorm(
        din2_din1_denorm_20_18) );
  fpu_denorm_3b i_fpu_denorm_17_15 ( .din1(din1[17:15]), .din2(din2[17:15]), 
        .din2_din1_nz(din2_din1_nz_17_15), .din2_din1_denorm(
        din2_din1_denorm_17_15) );
  fpu_denorm_3b i_fpu_denorm_14_12 ( .din1(din1[14:12]), .din2(din2[14:12]), 
        .din2_din1_nz(din2_din1_nz_14_12), .din2_din1_denorm(
        din2_din1_denorm_14_12) );
  fpu_denorm_3b i_fpu_denorm_11_9 ( .din1(din1[11:9]), .din2(din2[11:9]), 
        .din2_din1_nz(din2_din1_nz_11_9), .din2_din1_denorm(
        din2_din1_denorm_11_9) );
  fpu_denorm_3b i_fpu_denorm_8_6 ( .din1(din1[8:6]), .din2(din2[8:6]), 
        .din2_din1_nz(din2_din1_nz_8_6), .din2_din1_denorm(
        din2_din1_denorm_8_6) );
  fpu_denorm_3b i_fpu_denorm_5_3 ( .din1(din1[5:3]), .din2(din2[5:3]), 
        .din2_din1_nz(din2_din1_nz_5_3), .din2_din1_denorm(
        din2_din1_denorm_5_3) );
  fpu_denorm_3b i_fpu_denorm_2_0 ( .din1(din1[2:0]), .din2(din2[2:0]), 
        .din2_din1_nz(din2_din1_nz_2_0), .din2_din1_denorm(
        din2_din1_denorm_2_0) );
  fpu_denorm_3to1 i_fpu_denorm_53_45 ( .din2_din1_nz_hi(din2_din1_nz_53_51), 
        .din2_din1_denorm_hi(din2_din1_denorm_53_51), .din2_din1_nz_mid(
        din2_din1_nz_50_48), .din2_din1_denorm_mid(din2_din1_denorm_50_48), 
        .din2_din1_nz_lo(din2_din1_nz_47_45), .din2_din1_denorm_lo(
        din2_din1_denorm_47_45), .din2_din1_nz(din2_din1_nz_53_45), 
        .din2_din1_denorm(din2_din1_denorm_53_45) );
  fpu_denorm_3to1 i_fpu_denorm_44_36 ( .din2_din1_nz_hi(din2_din1_nz_44_42), 
        .din2_din1_denorm_hi(din2_din1_denorm_44_42), .din2_din1_nz_mid(
        din2_din1_nz_41_39), .din2_din1_denorm_mid(din2_din1_denorm_41_39), 
        .din2_din1_nz_lo(din2_din1_nz_38_36), .din2_din1_denorm_lo(
        din2_din1_denorm_38_36), .din2_din1_nz(din2_din1_nz_44_36), 
        .din2_din1_denorm(din2_din1_denorm_44_36) );
  fpu_denorm_3to1 i_fpu_denorm_35_27 ( .din2_din1_nz_hi(din2_din1_nz_35_33), 
        .din2_din1_denorm_hi(din2_din1_denorm_35_33), .din2_din1_nz_mid(
        din2_din1_nz_32_30), .din2_din1_denorm_mid(din2_din1_denorm_32_30), 
        .din2_din1_nz_lo(din2_din1_nz_29_27), .din2_din1_denorm_lo(
        din2_din1_denorm_29_27), .din2_din1_nz(din2_din1_nz_35_27), 
        .din2_din1_denorm(din2_din1_denorm_35_27) );
  fpu_denorm_3to1 i_fpu_denorm_26_18 ( .din2_din1_nz_hi(din2_din1_nz_26_24), 
        .din2_din1_denorm_hi(din2_din1_denorm_26_24), .din2_din1_nz_mid(
        din2_din1_nz_23_21), .din2_din1_denorm_mid(din2_din1_denorm_23_21), 
        .din2_din1_nz_lo(din2_din1_nz_20_18), .din2_din1_denorm_lo(
        din2_din1_denorm_20_18), .din2_din1_nz(din2_din1_nz_26_18), 
        .din2_din1_denorm(din2_din1_denorm_26_18) );
  fpu_denorm_3to1 i_fpu_denorm_17_9 ( .din2_din1_nz_hi(din2_din1_nz_17_15), 
        .din2_din1_denorm_hi(din2_din1_denorm_17_15), .din2_din1_nz_mid(
        din2_din1_nz_14_12), .din2_din1_denorm_mid(din2_din1_denorm_14_12), 
        .din2_din1_nz_lo(din2_din1_nz_11_9), .din2_din1_denorm_lo(
        din2_din1_denorm_11_9), .din2_din1_nz(din2_din1_nz_17_9), 
        .din2_din1_denorm(din2_din1_denorm_17_9) );
  fpu_denorm_3to1 i_fpu_denorm_8_0 ( .din2_din1_nz_hi(din2_din1_nz_8_6), 
        .din2_din1_denorm_hi(din2_din1_denorm_8_6), .din2_din1_nz_mid(
        din2_din1_nz_5_3), .din2_din1_denorm_mid(din2_din1_denorm_5_3), 
        .din2_din1_nz_lo(din2_din1_nz_2_0), .din2_din1_denorm_lo(
        din2_din1_denorm_2_0), .din2_din1_nz(din2_din1_nz_8_0), 
        .din2_din1_denorm(din2_din1_denorm_8_0) );
  fpu_denorm_3to1 i_fpu_denorm_53_27 ( .din2_din1_nz_hi(din2_din1_nz_53_45), 
        .din2_din1_denorm_hi(din2_din1_denorm_53_45), .din2_din1_nz_mid(
        din2_din1_nz_44_36), .din2_din1_denorm_mid(din2_din1_denorm_44_36), 
        .din2_din1_nz_lo(din2_din1_nz_35_27), .din2_din1_denorm_lo(
        din2_din1_denorm_35_27), .din2_din1_nz(din2_din1_nz_53_27), 
        .din2_din1_denorm(din2_din1_denorm_53_27) );
  fpu_denorm_3to1 i_fpu_denorm_26_0 ( .din2_din1_nz_hi(din2_din1_nz_26_18), 
        .din2_din1_denorm_hi(din2_din1_denorm_26_18), .din2_din1_nz_mid(
        din2_din1_nz_17_9), .din2_din1_denorm_mid(din2_din1_denorm_17_9), 
        .din2_din1_nz_lo(din2_din1_nz_8_0), .din2_din1_denorm_lo(
        din2_din1_denorm_8_0), .din2_din1_nz(din2_din1_nz_26_0), 
        .din2_din1_denorm(din2_din1_denorm_26_0) );
  GTECH_NOT I_0 ( .A(din2_din1_nz_53_27), .Z(N0) );
  GTECH_OR2 C10 ( .A(N4), .B(N5), .Z(din2_din1_denorm) );
  GTECH_OR2 C11 ( .A(N1), .B(N3), .Z(N4) );
  GTECH_AND2 C12 ( .A(din2_din1_nz_53_27), .B(din2_din1_denorm_53_27), .Z(N1)
         );
  GTECH_AND2 C13 ( .A(N0), .B(N2), .Z(N3) );
  GTECH_NOT I_1 ( .A(din2_din1_nz_26_0), .Z(N2) );
  GTECH_AND2 C15 ( .A(N0), .B(din2_din1_denorm_26_0), .Z(N5) );
  GTECH_NOT I_2 ( .A(din2_din1_denorm), .Z(din2_din1_denorm_inv) );
endmodule


module fpu_cnt_lead0_lvl1 ( din, din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0 );
  input [3:0] din;
  output din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8;

  GTECH_NOT I_0 ( .A(N2), .Z(din_3_0_eq_0) );
  GTECH_OR2 C10 ( .A(N1), .B(din[0]), .Z(N2) );
  GTECH_OR2 C11 ( .A(N0), .B(din[1]), .Z(N1) );
  GTECH_OR2 C12 ( .A(din[3]), .B(din[2]), .Z(N0) );
  GTECH_NOT I_1 ( .A(N3), .Z(din_3_2_eq_0) );
  GTECH_OR2 C14 ( .A(din[3]), .B(din[2]), .Z(N3) );
  GTECH_OR2 C15 ( .A(N6), .B(N8), .Z(lead0_4b_0) );
  GTECH_AND2 C16 ( .A(N4), .B(N5), .Z(N6) );
  GTECH_NOT I_2 ( .A(din_3_2_eq_0), .Z(N4) );
  GTECH_NOT I_3 ( .A(din[3]), .Z(N5) );
  GTECH_AND2 C19 ( .A(din_3_2_eq_0), .B(N7), .Z(N8) );
  GTECH_NOT I_4 ( .A(din[1]), .Z(N7) );
endmodule


module fpu_cnt_lead0_lvl2 ( din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, 
        din_3_0_eq_0, din_3_2_eq_0, lead0_4b_0_lo, din_7_0_eq_0, lead0_8b_1, 
        lead0_8b_0 );
  input din_7_4_eq_0, din_7_6_eq_0, lead0_4b_0_hi, din_3_0_eq_0, din_3_2_eq_0,
         lead0_4b_0_lo;
  output din_7_0_eq_0, lead0_8b_1, lead0_8b_0;
  wire   N0, N1, N2, N3, N4;

  GTECH_AND2 C9 ( .A(din_3_0_eq_0), .B(din_7_4_eq_0), .Z(din_7_0_eq_0) );
  GTECH_OR2 C10 ( .A(N1), .B(N2), .Z(lead0_8b_1) );
  GTECH_AND2 C11 ( .A(N0), .B(din_7_6_eq_0), .Z(N1) );
  GTECH_NOT I_0 ( .A(din_7_4_eq_0), .Z(N0) );
  GTECH_AND2 C13 ( .A(din_7_4_eq_0), .B(din_3_2_eq_0), .Z(N2) );
  GTECH_OR2 C14 ( .A(N3), .B(N4), .Z(lead0_8b_0) );
  GTECH_AND2 C15 ( .A(N0), .B(lead0_4b_0_hi), .Z(N3) );
  GTECH_AND2 C17 ( .A(din_7_4_eq_0), .B(lead0_4b_0_lo), .Z(N4) );
endmodule


module fpu_cnt_lead0_lvl3 ( din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, 
        lead0_8b_0_hi, din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, 
        lead0_8b_0_lo, din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0 );
  input din_15_8_eq_0, din_15_12_eq_0, lead0_8b_1_hi, lead0_8b_0_hi,
         din_7_0_eq_0, din_7_4_eq_0, lead0_8b_1_lo, lead0_8b_0_lo;
  output din_15_0_eq_0, lead0_16b_2, lead0_16b_1, lead0_16b_0;
  wire   N0, N1, N2, N3, N4, N5, N6;

  GTECH_AND2 C10 ( .A(din_7_0_eq_0), .B(din_15_8_eq_0), .Z(din_15_0_eq_0) );
  GTECH_OR2 C11 ( .A(N1), .B(N2), .Z(lead0_16b_2) );
  GTECH_AND2 C12 ( .A(N0), .B(din_15_12_eq_0), .Z(N1) );
  GTECH_NOT I_0 ( .A(din_15_8_eq_0), .Z(N0) );
  GTECH_AND2 C14 ( .A(din_15_8_eq_0), .B(din_7_4_eq_0), .Z(N2) );
  GTECH_OR2 C15 ( .A(N3), .B(N4), .Z(lead0_16b_1) );
  GTECH_AND2 C16 ( .A(N0), .B(lead0_8b_1_hi), .Z(N3) );
  GTECH_AND2 C18 ( .A(din_15_8_eq_0), .B(lead0_8b_1_lo), .Z(N4) );
  GTECH_OR2 C19 ( .A(N5), .B(N6), .Z(lead0_16b_0) );
  GTECH_AND2 C20 ( .A(N0), .B(lead0_8b_0_hi), .Z(N5) );
  GTECH_AND2 C22 ( .A(din_15_8_eq_0), .B(lead0_8b_0_lo), .Z(N6) );
endmodule


module fpu_cnt_lead0_lvl4 ( din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, 
        lead0_16b_1_hi, lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, 
        lead0_16b_2_lo, lead0_16b_1_lo, lead0_16b_0_lo, din_31_0_eq_0, 
        lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0 );
  input din_31_16_eq_0, din_31_24_eq_0, lead0_16b_2_hi, lead0_16b_1_hi,
         lead0_16b_0_hi, din_15_0_eq_0, din_15_8_eq_0, lead0_16b_2_lo,
         lead0_16b_1_lo, lead0_16b_0_lo;
  output din_31_0_eq_0, lead0_32b_3, lead0_32b_2, lead0_32b_1, lead0_32b_0;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8;

  GTECH_AND2 C11 ( .A(din_15_0_eq_0), .B(din_31_16_eq_0), .Z(din_31_0_eq_0) );
  GTECH_OR2 C12 ( .A(N1), .B(N2), .Z(lead0_32b_3) );
  GTECH_AND2 C13 ( .A(N0), .B(din_31_24_eq_0), .Z(N1) );
  GTECH_NOT I_0 ( .A(din_31_16_eq_0), .Z(N0) );
  GTECH_AND2 C15 ( .A(din_31_16_eq_0), .B(din_15_8_eq_0), .Z(N2) );
  GTECH_OR2 C16 ( .A(N3), .B(N4), .Z(lead0_32b_2) );
  GTECH_AND2 C17 ( .A(N0), .B(lead0_16b_2_hi), .Z(N3) );
  GTECH_AND2 C19 ( .A(din_31_16_eq_0), .B(lead0_16b_2_lo), .Z(N4) );
  GTECH_OR2 C20 ( .A(N5), .B(N6), .Z(lead0_32b_1) );
  GTECH_AND2 C21 ( .A(N0), .B(lead0_16b_1_hi), .Z(N5) );
  GTECH_AND2 C23 ( .A(din_31_16_eq_0), .B(lead0_16b_1_lo), .Z(N6) );
  GTECH_OR2 C24 ( .A(N7), .B(N8), .Z(lead0_32b_0) );
  GTECH_AND2 C25 ( .A(N0), .B(lead0_16b_0_hi), .Z(N7) );
  GTECH_AND2 C27 ( .A(din_31_16_eq_0), .B(lead0_16b_0_lo), .Z(N8) );
endmodule


module fpu_cnt_lead0_64b ( din, lead0 );
  input [63:0] din;
  output [5:0] lead0;
  wire   din_63_60_eq_0, din_63_62_eq_0, lead0_63_60_0, din_59_56_eq_0,
         din_59_58_eq_0, lead0_59_56_0, din_55_52_eq_0, din_55_54_eq_0,
         lead0_55_52_0, din_51_48_eq_0, din_51_50_eq_0, lead0_51_48_0,
         din_47_44_eq_0, din_47_46_eq_0, lead0_47_44_0, din_43_40_eq_0,
         din_43_42_eq_0, lead0_43_40_0, din_39_36_eq_0, din_39_38_eq_0,
         lead0_39_36_0, din_35_32_eq_0, din_35_34_eq_0, lead0_35_32_0,
         din_31_28_eq_0, din_31_30_eq_0, lead0_31_28_0, din_27_24_eq_0,
         din_27_26_eq_0, lead0_27_24_0, din_23_20_eq_0, din_23_22_eq_0,
         lead0_23_20_0, din_19_16_eq_0, din_19_18_eq_0, lead0_19_16_0,
         din_15_12_eq_0, din_15_14_eq_0, lead0_15_12_0, din_11_8_eq_0,
         din_11_10_eq_0, lead0_11_8_0, din_7_4_eq_0, din_7_6_eq_0, lead0_7_4_0,
         din_3_0_eq_0, din_3_2_eq_0, lead0_3_0_0, din_63_56_eq_0,
         lead0_63_56_1, lead0_63_56_0, din_55_48_eq_0, lead0_55_48_1,
         lead0_55_48_0, din_47_40_eq_0, lead0_47_40_1, lead0_47_40_0,
         din_39_32_eq_0, lead0_39_32_1, lead0_39_32_0, din_31_24_eq_0,
         lead0_31_24_1, lead0_31_24_0, din_23_16_eq_0, lead0_23_16_1,
         lead0_23_16_0, din_15_8_eq_0, lead0_15_8_1, lead0_15_8_0,
         din_7_0_eq_0, lead0_7_0_1, lead0_7_0_0, din_63_48_eq_0, lead0_63_48_2,
         lead0_63_48_1, lead0_63_48_0, din_47_32_eq_0, lead0_47_32_2,
         lead0_47_32_1, lead0_47_32_0, din_31_16_eq_0, lead0_31_16_2,
         lead0_31_16_1, lead0_31_16_0, din_15_0_eq_0, lead0_15_0_2,
         lead0_15_0_1, lead0_15_0_0, din_63_32_eq_0, lead0_63_32_3,
         lead0_63_32_2, lead0_63_32_1, lead0_63_32_0, din_31_0_eq_0,
         lead0_31_0_3, lead0_31_0_2, lead0_31_0_1, lead0_31_0_0, lead0_6, N0,
         N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16
;

  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_63_60 ( .din(din[63:60]), 
        .din_3_0_eq_0(din_63_60_eq_0), .din_3_2_eq_0(din_63_62_eq_0), 
        .lead0_4b_0(lead0_63_60_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_59_56 ( .din(din[59:56]), 
        .din_3_0_eq_0(din_59_56_eq_0), .din_3_2_eq_0(din_59_58_eq_0), 
        .lead0_4b_0(lead0_59_56_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_55_52 ( .din(din[55:52]), 
        .din_3_0_eq_0(din_55_52_eq_0), .din_3_2_eq_0(din_55_54_eq_0), 
        .lead0_4b_0(lead0_55_52_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_51_48 ( .din(din[51:48]), 
        .din_3_0_eq_0(din_51_48_eq_0), .din_3_2_eq_0(din_51_50_eq_0), 
        .lead0_4b_0(lead0_51_48_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_47_44 ( .din(din[47:44]), 
        .din_3_0_eq_0(din_47_44_eq_0), .din_3_2_eq_0(din_47_46_eq_0), 
        .lead0_4b_0(lead0_47_44_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_43_40 ( .din(din[43:40]), 
        .din_3_0_eq_0(din_43_40_eq_0), .din_3_2_eq_0(din_43_42_eq_0), 
        .lead0_4b_0(lead0_43_40_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_39_36 ( .din(din[39:36]), 
        .din_3_0_eq_0(din_39_36_eq_0), .din_3_2_eq_0(din_39_38_eq_0), 
        .lead0_4b_0(lead0_39_36_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_35_32 ( .din(din[35:32]), 
        .din_3_0_eq_0(din_35_32_eq_0), .din_3_2_eq_0(din_35_34_eq_0), 
        .lead0_4b_0(lead0_35_32_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_31_28 ( .din(din[31:28]), 
        .din_3_0_eq_0(din_31_28_eq_0), .din_3_2_eq_0(din_31_30_eq_0), 
        .lead0_4b_0(lead0_31_28_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_27_24 ( .din(din[27:24]), 
        .din_3_0_eq_0(din_27_24_eq_0), .din_3_2_eq_0(din_27_26_eq_0), 
        .lead0_4b_0(lead0_27_24_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_23_20 ( .din(din[23:20]), 
        .din_3_0_eq_0(din_23_20_eq_0), .din_3_2_eq_0(din_23_22_eq_0), 
        .lead0_4b_0(lead0_23_20_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_19_16 ( .din(din[19:16]), 
        .din_3_0_eq_0(din_19_16_eq_0), .din_3_2_eq_0(din_19_18_eq_0), 
        .lead0_4b_0(lead0_19_16_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_15_12 ( .din(din[15:12]), 
        .din_3_0_eq_0(din_15_12_eq_0), .din_3_2_eq_0(din_15_14_eq_0), 
        .lead0_4b_0(lead0_15_12_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_11_8 ( .din(din[11:8]), 
        .din_3_0_eq_0(din_11_8_eq_0), .din_3_2_eq_0(din_11_10_eq_0), 
        .lead0_4b_0(lead0_11_8_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_7_4 ( .din(din[7:4]), .din_3_0_eq_0(
        din_7_4_eq_0), .din_3_2_eq_0(din_7_6_eq_0), .lead0_4b_0(lead0_7_4_0)
         );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_3_0 ( .din(din[3:0]), .din_3_0_eq_0(
        din_3_0_eq_0), .din_3_2_eq_0(din_3_2_eq_0), .lead0_4b_0(lead0_3_0_0)
         );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_63_56 ( .din_7_4_eq_0(din_63_60_eq_0), .din_7_6_eq_0(din_63_62_eq_0), .lead0_4b_0_hi(lead0_63_60_0), .din_3_0_eq_0(
        din_59_56_eq_0), .din_3_2_eq_0(din_59_58_eq_0), .lead0_4b_0_lo(
        lead0_59_56_0), .din_7_0_eq_0(din_63_56_eq_0), .lead0_8b_1(
        lead0_63_56_1), .lead0_8b_0(lead0_63_56_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_55_48 ( .din_7_4_eq_0(din_55_52_eq_0), .din_7_6_eq_0(din_55_54_eq_0), .lead0_4b_0_hi(lead0_55_52_0), .din_3_0_eq_0(
        din_51_48_eq_0), .din_3_2_eq_0(din_51_50_eq_0), .lead0_4b_0_lo(
        lead0_51_48_0), .din_7_0_eq_0(din_55_48_eq_0), .lead0_8b_1(
        lead0_55_48_1), .lead0_8b_0(lead0_55_48_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_47_40 ( .din_7_4_eq_0(din_47_44_eq_0), .din_7_6_eq_0(din_47_46_eq_0), .lead0_4b_0_hi(lead0_47_44_0), .din_3_0_eq_0(
        din_43_40_eq_0), .din_3_2_eq_0(din_43_42_eq_0), .lead0_4b_0_lo(
        lead0_43_40_0), .din_7_0_eq_0(din_47_40_eq_0), .lead0_8b_1(
        lead0_47_40_1), .lead0_8b_0(lead0_47_40_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_39_32 ( .din_7_4_eq_0(din_39_36_eq_0), .din_7_6_eq_0(din_39_38_eq_0), .lead0_4b_0_hi(lead0_39_36_0), .din_3_0_eq_0(
        din_35_32_eq_0), .din_3_2_eq_0(din_35_34_eq_0), .lead0_4b_0_lo(
        lead0_35_32_0), .din_7_0_eq_0(din_39_32_eq_0), .lead0_8b_1(
        lead0_39_32_1), .lead0_8b_0(lead0_39_32_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_31_24 ( .din_7_4_eq_0(din_31_28_eq_0), .din_7_6_eq_0(din_31_30_eq_0), .lead0_4b_0_hi(lead0_31_28_0), .din_3_0_eq_0(
        din_27_24_eq_0), .din_3_2_eq_0(din_27_26_eq_0), .lead0_4b_0_lo(
        lead0_27_24_0), .din_7_0_eq_0(din_31_24_eq_0), .lead0_8b_1(
        lead0_31_24_1), .lead0_8b_0(lead0_31_24_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_23_16 ( .din_7_4_eq_0(din_23_20_eq_0), .din_7_6_eq_0(din_23_22_eq_0), .lead0_4b_0_hi(lead0_23_20_0), .din_3_0_eq_0(
        din_19_16_eq_0), .din_3_2_eq_0(din_19_18_eq_0), .lead0_4b_0_lo(
        lead0_19_16_0), .din_7_0_eq_0(din_23_16_eq_0), .lead0_8b_1(
        lead0_23_16_1), .lead0_8b_0(lead0_23_16_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_15_8 ( .din_7_4_eq_0(din_15_12_eq_0), 
        .din_7_6_eq_0(din_15_14_eq_0), .lead0_4b_0_hi(lead0_15_12_0), 
        .din_3_0_eq_0(din_11_8_eq_0), .din_3_2_eq_0(din_11_10_eq_0), 
        .lead0_4b_0_lo(lead0_11_8_0), .din_7_0_eq_0(din_15_8_eq_0), 
        .lead0_8b_1(lead0_15_8_1), .lead0_8b_0(lead0_15_8_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_7_0 ( .din_7_4_eq_0(din_7_4_eq_0), 
        .din_7_6_eq_0(din_7_6_eq_0), .lead0_4b_0_hi(lead0_7_4_0), 
        .din_3_0_eq_0(din_3_0_eq_0), .din_3_2_eq_0(din_3_2_eq_0), 
        .lead0_4b_0_lo(lead0_3_0_0), .din_7_0_eq_0(din_7_0_eq_0), .lead0_8b_1(
        lead0_7_0_1), .lead0_8b_0(lead0_7_0_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_63_48 ( .din_15_8_eq_0(
        din_63_56_eq_0), .din_15_12_eq_0(din_63_60_eq_0), .lead0_8b_1_hi(
        lead0_63_56_1), .lead0_8b_0_hi(lead0_63_56_0), .din_7_0_eq_0(
        din_55_48_eq_0), .din_7_4_eq_0(din_55_52_eq_0), .lead0_8b_1_lo(
        lead0_55_48_1), .lead0_8b_0_lo(lead0_55_48_0), .din_15_0_eq_0(
        din_63_48_eq_0), .lead0_16b_2(lead0_63_48_2), .lead0_16b_1(
        lead0_63_48_1), .lead0_16b_0(lead0_63_48_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_47_32 ( .din_15_8_eq_0(
        din_47_40_eq_0), .din_15_12_eq_0(din_47_44_eq_0), .lead0_8b_1_hi(
        lead0_47_40_1), .lead0_8b_0_hi(lead0_47_40_0), .din_7_0_eq_0(
        din_39_32_eq_0), .din_7_4_eq_0(din_39_36_eq_0), .lead0_8b_1_lo(
        lead0_39_32_1), .lead0_8b_0_lo(lead0_39_32_0), .din_15_0_eq_0(
        din_47_32_eq_0), .lead0_16b_2(lead0_47_32_2), .lead0_16b_1(
        lead0_47_32_1), .lead0_16b_0(lead0_47_32_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_31_16 ( .din_15_8_eq_0(
        din_31_24_eq_0), .din_15_12_eq_0(din_31_28_eq_0), .lead0_8b_1_hi(
        lead0_31_24_1), .lead0_8b_0_hi(lead0_31_24_0), .din_7_0_eq_0(
        din_23_16_eq_0), .din_7_4_eq_0(din_23_20_eq_0), .lead0_8b_1_lo(
        lead0_23_16_1), .lead0_8b_0_lo(lead0_23_16_0), .din_15_0_eq_0(
        din_31_16_eq_0), .lead0_16b_2(lead0_31_16_2), .lead0_16b_1(
        lead0_31_16_1), .lead0_16b_0(lead0_31_16_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_15_0 ( .din_15_8_eq_0(din_15_8_eq_0), 
        .din_15_12_eq_0(din_15_12_eq_0), .lead0_8b_1_hi(lead0_15_8_1), 
        .lead0_8b_0_hi(lead0_15_8_0), .din_7_0_eq_0(din_7_0_eq_0), 
        .din_7_4_eq_0(din_7_4_eq_0), .lead0_8b_1_lo(lead0_7_0_1), 
        .lead0_8b_0_lo(lead0_7_0_0), .din_15_0_eq_0(din_15_0_eq_0), 
        .lead0_16b_2(lead0_15_0_2), .lead0_16b_1(lead0_15_0_1), .lead0_16b_0(
        lead0_15_0_0) );
  fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_63_32 ( .din_31_16_eq_0(
        din_63_48_eq_0), .din_31_24_eq_0(din_63_56_eq_0), .lead0_16b_2_hi(
        lead0_63_48_2), .lead0_16b_1_hi(lead0_63_48_1), .lead0_16b_0_hi(
        lead0_63_48_0), .din_15_0_eq_0(din_47_32_eq_0), .din_15_8_eq_0(
        din_47_40_eq_0), .lead0_16b_2_lo(lead0_47_32_2), .lead0_16b_1_lo(
        lead0_47_32_1), .lead0_16b_0_lo(lead0_47_32_0), .din_31_0_eq_0(
        din_63_32_eq_0), .lead0_32b_3(lead0_63_32_3), .lead0_32b_2(
        lead0_63_32_2), .lead0_32b_1(lead0_63_32_1), .lead0_32b_0(
        lead0_63_32_0) );
  fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_31_0 ( .din_31_16_eq_0(
        din_31_16_eq_0), .din_31_24_eq_0(din_31_24_eq_0), .lead0_16b_2_hi(
        lead0_31_16_2), .lead0_16b_1_hi(lead0_31_16_1), .lead0_16b_0_hi(
        lead0_31_16_0), .din_15_0_eq_0(din_15_0_eq_0), .din_15_8_eq_0(
        din_15_8_eq_0), .lead0_16b_2_lo(lead0_15_0_2), .lead0_16b_1_lo(
        lead0_15_0_1), .lead0_16b_0_lo(lead0_15_0_0), .din_31_0_eq_0(
        din_31_0_eq_0), .lead0_32b_3(lead0_31_0_3), .lead0_32b_2(lead0_31_0_2), 
        .lead0_32b_1(lead0_31_0_1), .lead0_32b_0(lead0_31_0_0) );
  GTECH_AND2 C13 ( .A(din_63_32_eq_0), .B(din_31_0_eq_0), .Z(lead0_6) );
  GTECH_AND2 C14 ( .A(N0), .B(din_63_32_eq_0), .Z(lead0[5]) );
  GTECH_NOT I_0 ( .A(lead0_6), .Z(N0) );
  GTECH_OR2 C16 ( .A(N2), .B(N4), .Z(lead0[4]) );
  GTECH_AND2 C17 ( .A(N1), .B(din_63_48_eq_0), .Z(N2) );
  GTECH_NOT I_1 ( .A(din_63_32_eq_0), .Z(N1) );
  GTECH_AND2 C19 ( .A(N3), .B(N0), .Z(N4) );
  GTECH_AND2 C20 ( .A(din_63_32_eq_0), .B(din_31_16_eq_0), .Z(N3) );
  GTECH_OR2 C22 ( .A(N5), .B(N7), .Z(lead0[3]) );
  GTECH_AND2 C23 ( .A(N1), .B(lead0_63_32_3), .Z(N5) );
  GTECH_AND2 C25 ( .A(N6), .B(N0), .Z(N7) );
  GTECH_AND2 C26 ( .A(din_63_32_eq_0), .B(lead0_31_0_3), .Z(N6) );
  GTECH_OR2 C28 ( .A(N8), .B(N10), .Z(lead0[2]) );
  GTECH_AND2 C29 ( .A(N1), .B(lead0_63_32_2), .Z(N8) );
  GTECH_AND2 C31 ( .A(N9), .B(N0), .Z(N10) );
  GTECH_AND2 C32 ( .A(din_63_32_eq_0), .B(lead0_31_0_2), .Z(N9) );
  GTECH_OR2 C34 ( .A(N11), .B(N13), .Z(lead0[1]) );
  GTECH_AND2 C35 ( .A(N1), .B(lead0_63_32_1), .Z(N11) );
  GTECH_AND2 C37 ( .A(N12), .B(N0), .Z(N13) );
  GTECH_AND2 C38 ( .A(din_63_32_eq_0), .B(lead0_31_0_1), .Z(N12) );
  GTECH_OR2 C40 ( .A(N14), .B(N16), .Z(lead0[0]) );
  GTECH_AND2 C41 ( .A(N1), .B(lead0_63_32_0), .Z(N14) );
  GTECH_AND2 C43 ( .A(N15), .B(N0), .Z(N16) );
  GTECH_AND2 C44 ( .A(din_63_32_eq_0), .B(lead0_31_0_0), .Z(N15) );
endmodule


module dffe_SIZE58 ( din, en, clk, q, se, si, so );
  input [57:0] din;
  output [57:0] q;
  input [57:0] si;
  output [57:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63;
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N63) );
  SELECT_OP C247 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C255 ( .A(N3), .B(N2), .Z(N62) );
  GTECH_NOT I_2 ( .A(N62), .Z(N63) );
endmodule


module fpu_add_frac_dp ( inq_in1, inq_in2, a1stg_step, a1stg_sngop, 
        a1stg_expadd3_11, a1stg_norm_dbl_in1, a1stg_denorm_dbl_in1, 
        a1stg_norm_sng_in1, a1stg_denorm_sng_in1, a1stg_norm_dbl_in2, 
        a1stg_denorm_dbl_in2, a1stg_norm_sng_in2, a1stg_denorm_sng_in2, 
        a1stg_intlngop, a2stg_frac1_in_frac1, a2stg_frac1_in_frac2, 
        a1stg_2nan_in_inv, a1stg_faddsubop_inv, a2stg_frac1_in_qnan, 
        a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, a6stg_step, 
        a2stg_frac2_in_frac1, a2stg_frac2_in_qnan, a2stg_shr_cnt_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int, 
        a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max, 
        a2stg_expadd_11, a2stg_sub_step, a2stg_fracadd_frac2_inv_in, 
        a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2, 
        a2stg_fracadd_cin_in, a2stg_exp, a2stg_expdec_neq_0, a3stg_faddsubopa, 
        a3stg_sub_in, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, a3stg_exp_0, 
        a4stg_rnd_frac_add_inv, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, 
        a4stg_rnd_sng, a4stg_rnd_dbl, a4stg_shl_cnt_in, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0, 
        fadd_clken_l, rclk, a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, 
        a1stg_in2_eq_in1_exp, a2stg_frac2_63, a2stg_frac2hi_neq_0, 
        a2stg_frac2lo_neq_0, a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a3stg_denorm, 
        a3stg_denorm_inv, a3stg_lead0, a4stg_round, a4stg_shl_cnt, 
        a4stg_denorm_inv, a3stg_inc_exp_inv, a3stg_same_exp_inv, 
        a3stg_dec_exp_inv, a4stg_rnd_frac_40, a4stg_rnd_frac_39, 
        a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_rndadd_cout, 
        a4stg_frac_9_0_nx, a4stg_frac_dbl_nx, a4stg_frac_38_0_nx, 
        a4stg_frac_sng_nx, a4stg_frac_neq_0, a4stg_shl_data_neq_0, 
        add_of_out_cout, add_frac_out, se, si, so );
  input [62:0] inq_in1;
  input [63:0] inq_in2;
  input [5:0] a2stg_shr_cnt_in;
  input [5:0] a2stg_exp;
  input [1:0] a3stg_faddsubopa;
  input [9:0] a4stg_shl_cnt_in;
  output [5:0] a3stg_lead0;
  output [5:0] a4stg_shl_cnt;
  output [63:0] add_frac_out;
  input a1stg_step, a1stg_sngop, a1stg_expadd3_11, a1stg_norm_dbl_in1,
         a1stg_denorm_dbl_in1, a1stg_norm_sng_in1, a1stg_denorm_sng_in1,
         a1stg_norm_dbl_in2, a1stg_denorm_dbl_in2, a1stg_norm_sng_in2,
         a1stg_denorm_sng_in2, a1stg_intlngop, a2stg_frac1_in_frac1,
         a2stg_frac1_in_frac2, a1stg_2nan_in_inv, a1stg_faddsubop_inv,
         a2stg_frac1_in_qnan, a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl,
         a6stg_step, a2stg_frac2_in_frac1, a2stg_frac2_in_qnan,
         a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_expadd_11, a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a2stg_expdec_neq_0, a3stg_sub_in,
         a3stg_exp10_0_eq0, a3stg_exp10_1_eq0, a3stg_exp_0,
         a4stg_rnd_frac_add_inv, a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0,
         fadd_clken_l, rclk, se, si;
  output a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, a1stg_in2_eq_in1_exp,
         a2stg_frac2_63, a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0,
         a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, a3stg_denorm, a3stg_denorm_inv,
         a4stg_round, a4stg_denorm_inv, a3stg_inc_exp_inv, a3stg_same_exp_inv,
         a3stg_dec_exp_inv, a4stg_rnd_frac_40, a4stg_rnd_frac_39,
         a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_rndadd_cout,
         a4stg_frac_9_0_nx, a4stg_frac_dbl_nx, a4stg_frac_38_0_nx,
         a4stg_frac_sng_nx, a4stg_frac_neq_0, a4stg_shl_data_neq_0,
         add_of_out_cout, so;
  wire   se_l, clk, a1stg_in2_gt_in1, N0, N1, a2stg_fsdtoi_nx,
         a2stg_nx_neq0_84_tmp_4_54, a2stg_nx_neq0_84_tmp_4_53,
         a2stg_nx_neq0_84_tmp_4_52, a2stg_nx_neq0_84_tmp_4_51,
         a2stg_nx_neq0_84_tmp_4_50, a2stg_nx_neq0_84_tmp_4_49,
         a2stg_nx_neq0_84_tmp_4_48, a2stg_nx_neq0_84_tmp_5_52,
         a2stg_nx_neq0_84_tmp_5_51, a2stg_nx_neq0_84_tmp_5_50,
         a2stg_nx_neq0_84_tmp_6_51, a2stg_fsdtoix_nx, a2stg_shr_60_0_neq_0,
         a2stg_fracadd_frac2_inv, a2stg_fracadd_frac2_inv_shr1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, a2stg_fracadd_cin, a3stg_ld0_dnrm_10, a3stg_denorma,
         a3stg_denorm_inva, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, a3stg_suba, a3stg_sub, a4stg_round_in,
         N130, a3stg_inc_exp_inva, a3stg_fsame_exp_inv, a3stg_fdec_exp_inv,
         a4stg_rnd_frac_63, a4stg_rnd_frac_62, a4stg_rnd_frac_61,
         a4stg_rnd_frac_60, a4stg_rnd_frac_59, a4stg_rnd_frac_58,
         a4stg_rnd_frac_57, a4stg_rnd_frac_56, a4stg_rnd_frac_55,
         a4stg_rnd_frac_54, a4stg_rnd_frac_53, a4stg_rnd_frac_52,
         a4stg_rnd_frac_51, a4stg_rnd_frac_50, a4stg_rnd_frac_49,
         a4stg_rnd_frac_48, a4stg_rnd_frac_47, a4stg_rnd_frac_46,
         a4stg_rnd_frac_45, a4stg_rnd_frac_44, a4stg_rnd_frac_43,
         a4stg_rnd_frac_42, a4stg_rnd_frac_41, a4stg_rnd_frac_9,
         a4stg_rnd_frac_8, a4stg_rnd_frac_7, a4stg_rnd_frac_6,
         a4stg_rnd_frac_5, a4stg_rnd_frac_4, a4stg_rnd_frac_3,
         a4stg_rnd_frac_2, a4stg_rnd_frac_1, a4stg_rnd_frac_0,
         a5stg_frac_out_rndadd, a5stg_frac_out_rnd_frac, a5stg_in_of,
         a5stg_frac_out_shl, a5stg_to_0, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279,
         N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290,
         N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301,
         N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312,
         N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323,
         N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367,
         N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378,
         N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422,
         N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433,
         N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444,
         N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455,
         N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477,
         N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510,
         N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521,
         N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532,
         N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543,
         N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554,
         N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565,
         N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576,
         N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587,
         N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598,
         N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609,
         N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620,
         N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631,
         N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697,
         N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752,
         N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763,
         N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034,
         N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074,
         N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084,
         N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094,
         N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104,
         N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114,
         N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124,
         N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134,
         N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144,
         N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154,
         N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164,
         N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174,
         N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184,
         N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194,
         N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204,
         N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214,
         N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224,
         N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234,
         N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244,
         N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254,
         N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264,
         N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274,
         N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284,
         N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294,
         N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304,
         N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314,
         N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324,
         N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334,
         N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344,
         N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354,
         N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364,
         N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374,
         N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394,
         N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404,
         N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414,
         N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424,
         N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434,
         N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444,
         N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454,
         N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464,
         N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474,
         N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484,
         N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494,
         N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504,
         N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514,
         N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524,
         N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534,
         N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544,
         N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554,
         N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564,
         N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574,
         N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584,
         N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594,
         N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604,
         N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614,
         N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624,
         N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634,
         N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644,
         N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654,
         N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664,
         N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674,
         N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684,
         N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694,
         N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704,
         N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714,
         N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724,
         N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734,
         N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744,
         N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754,
         N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764,
         N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774,
         N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784,
         N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794,
         N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804,
         N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814,
         N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824,
         N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834,
         N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844,
         N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854,
         N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864,
         N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874,
         N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884,
         N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894,
         N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904,
         N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914,
         N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924,
         N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934,
         N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944,
         N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954,
         N1955, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964,
         N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974,
         N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984,
         N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992, N1993, N1994,
         N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, N2003, N2004,
         N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014,
         N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024,
         N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034,
         N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044,
         N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054,
         N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064,
         N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074,
         N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083, N2084,
         N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093, N2094,
         N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104,
         N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114,
         N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124,
         N2125, N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134,
         N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144,
         N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154,
         N2155, N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164,
         N2165, N2166, N2167, N2168, N2169, N2170, N2171, N2172, N2173, N2174,
         N2175, N2176, N2177, N2178, N2179, N2180, N2181, N2182, N2183, N2184,
         N2185, N2186, N2187, N2188, N2189, N2190, N2191, N2192, N2193, N2194,
         N2195, N2196, N2197, N2198, N2199, N2200, N2201, N2202, N2203, N2204,
         N2205, N2206, N2207, N2208, N2209, N2210, N2211, N2212, N2213, N2214,
         N2215, N2216, N2217, N2218, N2219, N2220, N2221, N2222, N2223, N2224,
         N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234,
         N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244,
         N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254,
         N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264,
         N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274,
         N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284,
         N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294,
         N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304,
         N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314,
         N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324,
         N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334,
         N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344,
         N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354,
         N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364,
         N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374,
         N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384,
         N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394,
         N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404,
         N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414,
         N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424,
         N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434,
         N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444,
         N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454,
         N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464,
         N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474,
         N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484,
         N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494,
         N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504,
         N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514,
         N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524,
         N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534,
         N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544,
         N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554,
         N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564,
         N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574,
         N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584,
         N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594,
         N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604,
         N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614,
         N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624,
         N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634,
         N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644,
         N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654,
         N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664,
         N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674,
         N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684,
         N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694,
         N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704,
         N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714,
         N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724,
         N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734,
         N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744,
         N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754,
         N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764,
         N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774,
         N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784,
         N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794,
         N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804,
         N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814,
         N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824,
         N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834,
         N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844,
         N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854,
         N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864,
         N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874,
         N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884,
         N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894,
         N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904,
         N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914,
         N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924,
         N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934,
         N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944,
         N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954,
         N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964,
         N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974,
         N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984,
         N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994,
         N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004,
         N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014,
         N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024,
         N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034,
         N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044,
         N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054,
         N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064,
         N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074,
         N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084,
         N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094,
         N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104,
         N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114,
         N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124,
         N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134,
         N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144,
         N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154,
         N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164,
         N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174,
         N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184,
         N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194,
         N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204,
         N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214,
         N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224,
         N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234,
         N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244,
         N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254,
         N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264,
         N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274,
         N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284,
         N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294,
         N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304,
         N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314,
         N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324,
         N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334,
         N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344,
         N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354,
         N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364,
         N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374,
         N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384,
         N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394,
         N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404,
         N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414,
         N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424,
         N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434,
         N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N3444,
         N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454,
         N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464,
         N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3474,
         N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484,
         N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494,
         N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504,
         N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514,
         N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524,
         N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534,
         N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544,
         N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554,
         N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564,
         N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574,
         N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584,
         N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594,
         N3595, N3596, N3597, N3598, N3599, N3600, N3601, N3602, N3603, N3604,
         N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614,
         N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624,
         N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634,
         N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644,
         N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654,
         N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664,
         N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674,
         N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684,
         N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694,
         N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704,
         N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714,
         N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724,
         N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734,
         N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744,
         N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754,
         N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764,
         N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774,
         N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784,
         N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794,
         N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804,
         N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814,
         N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824,
         N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834,
         N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3843, N3844,
         N3845, N3846, N3847, N3848, N3849, N3850, N3851, N3852, N3853, N3854,
         N3855, N3856, N3857, N3858, N3859, N3860, N3861, N3862, N3863, N3864,
         N3865, N3866, N3867, N3868, N3869, N3870, N3871, N3872, N3873, N3874,
         N3875, N3876, N3877, N3878, N3879, N3880, N3881, N3882, N3883, N3884,
         N3885, N3886, N3887, N3888, N3889, N3890, N3891, N3892, N3893, N3894,
         N3895, N3896, N3897, N3898, N3899, N3900, N3901, N3902, N3903, N3904,
         N3905, N3906, N3907, N3908, N3909, N3910, N3911, N3912, N3913, N3914,
         N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3922, N3923, N3924,
         N3925, N3926, N3927, N3928, N3929, N3930, N3931, N3932, N3933, N3934,
         N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944,
         N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954,
         N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964,
         N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974,
         N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984,
         N3985, N3986, N3987, N3988, N3989, N3990, N3991, N3992, N3993, N3994,
         N3995, N3996, N3997, N3998, N3999, N4000, N4001, N4002, N4003, N4004,
         N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014,
         N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4022, N4023, N4024,
         N4025, N4026, N4027, N4028, N4029, N4030, N4031, N4032, N4033, N4034,
         N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4043, N4044,
         N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054,
         N4055, N4056, N4057, N4058, N4059, N4060, N4061, N4062, N4063, N4064,
         N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073, N4074,
         N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083, N4084,
         N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093, N4094,
         N4095, N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104,
         N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114,
         N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124,
         N4125, N4126, N4127, N4128, N4129, N4130, N4131, N4132, N4133, N4134,
         N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143, N4144,
         N4145, N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154,
         N4155, N4156, N4157, N4158, N4159, N4160, N4161, N4162, N4163, N4164,
         N4165, N4166, N4167, N4168, N4169, N4170, N4171, N4172, N4173, N4174,
         N4175, N4176, N4177, N4178, N4179, N4180, N4181, N4182, N4183, N4184,
         N4185, N4186, N4187, N4188, N4189, N4190, N4191, N4192, N4193, N4194,
         N4195, N4196, N4197, N4198, N4199, N4200, N4201, N4202, N4203, N4204,
         N4205, N4206, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214,
         N4215, N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224,
         N4225, N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234,
         N4235, N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244,
         N4245, N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254,
         N4255, N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264,
         N4265, N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274,
         N4275, N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284,
         N4285, N4286, N4287, N4288, N4289, N4290, N4291, N4292, N4293, N4294,
         N4295, N4296, N4297, N4298, N4299, N4300, N4301, N4302, N4303, N4304,
         N4305, N4306, N4307, N4308, N4309, N4310, N4311, N4312, N4313, N4314,
         N4315, N4316, N4317, N4318, N4319, N4320, N4321, N4322, N4323, N4324,
         N4325, N4326, N4327, N4328, N4329, N4330, N4331, N4332, N4333, N4334,
         N4335, N4336, N4337, N4338, N4339, N4340, N4341, N4342, N4343, N4344,
         N4345, N4346, N4347, N4348, N4349, N4350, N4351, N4352, N4353, N4354,
         N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364,
         N4365, N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374,
         N4375, N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4383, N4384,
         N4385, N4386, N4387, N4388, N4389, N4390, N4391, N4392, N4393, N4394,
         N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402, N4403, N4404,
         N4405, N4406, N4407, N4408, N4409, N4410, N4411, N4412, N4413, N4414,
         N4415, N4416, N4417, N4418, N4419, N4420, N4421, N4422, N4423, N4424,
         N4425, N4426, N4427, N4428, N4429, N4430, N4431, N4432, N4433, N4434,
         N4435, N4436, N4437, N4438, N4439, N4440, N4441, N4442, N4443, N4444,
         N4445, N4446, N4447, N4448, N4449, N4450, N4451, N4452, N4453, N4454,
         N4455, N4456, N4457, N4458, N4459, N4460, N4461, N4462, N4463, N4464,
         N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4474,
         N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483, N4484,
         N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493, N4494,
         N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504,
         N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514,
         N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524,
         N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534,
         N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544,
         N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554,
         N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564,
         N4565, N4566, N4567, N4568, N4569, N4570, N4571, N4572, N4573, N4574,
         N4575, N4576, N4577, N4578, N4579, N4580, N4581, N4582, N4583, N4584,
         N4585, N4586, N4587, N4588, N4589, N4590, N4591, N4592, N4593, N4594,
         N4595, N4596, N4597, N4598, N4599, N4600, N4601, N4602, N4603, N4604,
         N4605, N4606, N4607, N4608, N4609, N4610, N4611, N4612, N4613, N4614,
         N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624,
         N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634,
         N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644,
         N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4654,
         N4655, N4656, N4657, N4658, N4659, N4660, N4661, N4662, N4663, N4664,
         N4665, N4666, N4667, N4668, N4669, N4670, N4671, N4672, N4673, N4674,
         N4675, N4676, N4677, N4678, N4679, N4680, N4681, N4682, N4683, N4684,
         N4685, N4686, N4687, N4688, N4689, N4690, N4691, N4692, N4693, N4694,
         N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4703, N4704,
         N4705, N4706, N4707, N4708, N4709, N4710, N4711, N4712, N4713, N4714,
         N4715, N4716, N4717, N4718, N4719, N4720, N4721, N4722, N4723, N4724,
         N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734,
         N4735, N4736, N4737, N4738, N4739, N4740, N4741, N4742, N4743, N4744,
         N4745, N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754,
         N4755, N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764,
         N4765, N4766, N4767, N4768, N4769, N4770, N4771, N4772, N4773, N4774,
         N4775, N4776, N4777, N4778, N4779, N4780, N4781, N4782, N4783, N4784,
         N4785, N4786, N4787, N4788, N4789, N4790, N4791, N4792, N4793, N4794,
         N4795, N4796, N4797, N4798, N4799, N4800, N4801, N4802, N4803, N4804,
         N4805, N4806, N4807, N4808, N4809, N4810, N4811, N4812, N4813, N4814,
         N4815, N4816, N4817, N4818, N4819, N4820, N4821, N4822, N4823, N4824,
         N4825, N4826, N4827, N4828, N4829, N4830, N4831, N4832, N4833, N4834,
         N4835, N4836, N4837, N4838, N4839, N4840, N4841, N4842, N4843, N4844,
         N4845, N4846, N4847, N4848, N4849, N4850, N4851, N4852, N4853, N4854,
         N4855, N4856, N4857, N4858, N4859, N4860, N4861, N4862, N4863, N4864,
         N4865, N4866, N4867, N4868, N4869, N4870, N4871, N4872, N4873, N4874,
         N4875, N4876, N4877, N4878, N4879, N4880, N4881, N4882, N4883, N4884,
         N4885, N4886, N4887, N4888, N4889, N4890, N4891, N4892, N4893, N4894,
         N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4902, N4903, N4904,
         N4905, N4906, N4907, N4908, N4909, N4910, N4911, N4912, N4913, N4914,
         N4915, N4916, N4917, N4918, N4919, N4920, N4921, N4922, N4923, N4924,
         N4925, N4926, N4927, N4928, N4929, N4930, N4931, N4932, N4933, N4934,
         N4935, N4936, N4937, N4938, N4939, N4940, N4941, N4942, N4943, N4944,
         N4945, N4946, N4947, N4948, N4949, N4950, N4951, N4952, N4953, N4954,
         N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4962, N4963, N4964,
         N4965, N4966, N4967, N4968, N4969, N4970, N4971, N4972, N4973, N4974,
         N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984,
         N4985, N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994,
         N4995, N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5003, N5004,
         N5005, N5006, N5007, N5008, N5009, N5010, N5011, N5012, N5013, N5014,
         N5015, N5016, N5017, N5018, N5019, N5020, N5021, N5022, N5023, N5024,
         N5025, N5026, N5027, N5028, N5029, N5030, N5031, N5032, N5033, N5034,
         N5035, N5036, N5037, N5038, N5039, N5040, N5041, N5042, N5043, N5044,
         N5045, N5046, N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054,
         N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5064,
         N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074,
         N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084,
         N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094,
         N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104,
         N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114,
         N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124,
         N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5134,
         N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144,
         N5145, N5146, N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154,
         N5155, N5156, N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164,
         N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174,
         N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184,
         N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5194,
         N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204,
         N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5214,
         N5215, N5216, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224,
         N5225, N5226, N5227, N5228, N5229, N5230, N5231, N5232, N5233, N5234,
         N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244,
         N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252, N5253, N5254,
         N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264,
         N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272, N5273, N5274,
         N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282, N5283, N5284,
         N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294,
         N5295, N5296, N5297, N5298, N5299, N5300, N5301, N5302, N5303, N5304,
         N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5313, N5314,
         N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324,
         N5325, N5326, N5327, N5328, N5329, N5330, N5331, N5332, N5333, N5334,
         N5335, N5336, N5337, N5338, N5339, N5340, N5341, N5342, N5343, N5344,
         N5345, N5346, N5347, N5348, N5349, N5350, N5351, N5352, N5353, N5354,
         N5355, N5356, N5357, N5358, N5359, N5360, N5361, N5362, N5363, N5364,
         N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5372, N5373, N5374,
         N5375, N5376, N5377, N5378, N5379, N5380, N5381, N5382, N5383, N5384,
         N5385, N5386, N5387, N5388, N5389, N5390, N5391, N5392, N5393, N5394,
         N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402, N5403, N5404,
         N5405, N5406, N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414,
         N5415, N5416, N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424,
         N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5434,
         N5435, N5436, N5437, N5438, N5439, N5440, N5441, N5442, N5443, N5444,
         N5445, N5446, N5447, N5448, N5449, N5450, N5451, N5452, N5453, N5454,
         N5455, N5456, N5457, N5458, N5459, N5460, N5461, N5462, N5463, N5464,
         N5465, N5466, N5467, N5468, N5469, N5470, N5471, N5472, N5473, N5474,
         N5475, N5476, N5477, N5478, N5479, N5480, N5481, N5482, N5483, N5484,
         N5485, N5486, N5487, N5488, N5489, N5490, N5491, N5492, N5493, N5494,
         N5495, N5496, N5497, N5498, N5499, N5500, N5501, N5502, N5503, N5504,
         N5505, N5506, N5507, N5508, N5509, N5510, N5511, N5512, N5513, N5514,
         N5515, N5516, N5517, N5518, N5519, N5520, N5521, N5522, N5523, N5524,
         N5525, N5526, N5527, N5528, N5529, N5530, N5531, N5532, N5533, N5534,
         N5535, N5536, N5537, N5538, N5539, N5540, N5541, N5542, N5543, N5544,
         N5545, N5546, N5547, N5548, N5549, N5550, N5551, N5552, N5553, N5554,
         N5555, N5556, N5557, N5558, N5559, N5560, N5561, N5562, N5563, N5564,
         N5565, N5566, N5567, N5568, N5569, N5570, N5571, N5572, N5573, N5574,
         N5575, N5576, N5577, N5578, N5579, N5580, N5581, N5582, N5583, N5584,
         N5585, N5586, N5587, N5588, N5589, N5590, N5591, N5592, N5593, N5594,
         N5595, N5596, N5597, N5598, N5599, N5600, N5601, N5602, N5603, N5604,
         N5605, N5606, N5607, N5608, N5609, N5610, N5611, N5612, N5613, N5614,
         N5615, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5623, N5624,
         N5625, N5626, N5627, N5628, N5629, N5630, N5631, N5632, N5633, N5634,
         N5635, N5636, N5637, N5638, N5639, N5640, N5641, N5642, N5643, N5644,
         N5645, N5646, N5647, N5648, N5649, N5650, N5651, N5652, N5653, N5654,
         N5655, N5656, N5657, N5658, N5659, N5660, N5661, N5662, N5663, N5664,
         N5665, N5666, N5667, N5668, N5669, N5670, N5671, N5672, N5673, N5674,
         N5675, N5676, N5677, N5678, N5679, N5680, N5681, N5682, N5683, N5684,
         N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692, N5693, N5694,
         N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702, N5703, N5704,
         N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712, N5713, N5714,
         N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722, N5723, N5724,
         N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732, N5733, N5734,
         N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742, N5743, N5744,
         N5745, N5746, N5747, N5748, N5749, N5750, N5751, N5752, N5753, N5754,
         N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762, N5763, N5764,
         N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772, N5773, N5774,
         N5775, N5776, N5777, N5778, N5779, N5780, N5781, N5782, N5783, N5784,
         N5785, N5786, N5787, N5788, N5789, N5790, N5791, N5792, N5793, N5794,
         N5795, N5796, N5797, N5798, N5799, N5800, N5801, N5802, N5803, N5804,
         N5805, N5806, N5807, N5808, N5809, N5810, N5811, N5812, N5813, N5814,
         N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824,
         N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834,
         N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842, N5843, N5844,
         N5845, N5846, N5847, N5848, N5849, N5850, N5851, N5852, N5853, N5854,
         N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862, N5863, N5864,
         N5865, N5866, N5867, N5868, N5869, N5870, N5871, N5872, N5873, N5874,
         N5875, N5876, N5877, N5878, N5879, N5880, N5881, N5882, N5883, N5884,
         N5885, N5886, N5887, N5888, N5889, N5890, N5891, N5892, N5893, N5894,
         N5895, N5896, N5897, N5898, N5899, N5900, N5901, N5902, N5903, N5904,
         N5905, N5906, N5907, N5908, N5909, N5910, N5911, N5912, N5913, N5914,
         N5915, N5916, N5917, N5918, N5919, N5920, N5921, N5922, N5923, N5924,
         N5925, N5926, N5927, N5928, N5929, N5930, N5931, N5932, N5933, N5934,
         N5935, N5936, N5937, N5938, N5939, N5940, N5941, N5942, N5943, N5944,
         N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954,
         N5955, N5956, N5957, N5958, N5959, N5960, N5961, N5962, N5963, N5964,
         N5965, N5966, N5967, N5968, N5969, N5970, N5971, N5972, N5973, N5974,
         N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5982, N5983, N5984,
         N5985, N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994,
         N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003, N6004,
         N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012, N6013, N6014,
         N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022, N6023, N6024,
         N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034,
         N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6042, N6043, N6044,
         N6045, N6046, N6047, N6048, N6049, N6050, N6051, N6052, N6053, N6054,
         N6055, N6056, N6057, N6058, N6059, N6060, N6061, N6062, N6063, N6064,
         N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073, N6074,
         N6075, N6076, N6077, N6078, N6079, N6080, N6081, N6082, N6083, N6084,
         N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6092, N6093, N6094,
         N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104,
         N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114,
         N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124,
         N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134,
         N6135, N6136, N6137, N6138, N6139, N6140, N6141, N6142, N6143, N6144,
         N6145, N6146, N6147, N6148, N6149, N6150, N6151, N6152, N6153, N6154,
         N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163,
         net14641, net14642, net14643, net14644, net14645, net14646, net14647,
         net14648, net14649, net14650, net14651, net14652, net14653, net14654,
         net14655, net14656, net14657, net14658, net14659, net14660, net14661,
         net14662, net14663, net14664, net14665, net14666, net14667, net14668,
         net14669, net14670, net14671, net14672, net14673, net14674, net14675,
         net14676, net14677, net14678, net14679, net14680, net14681, net14682,
         net14683, net14684, net14685, net14686, net14687, net14688, net14689,
         net14690, net14691, net14692, net14693, net14694, net14695, net14696,
         net14697, net14698, net14699, net14700, net14701, net14702, net14703,
         net14704, net14705, net14706, net14707, net14708, net14709, net14710,
         net14711, net14712, net14713, net14714, net14715, net14716, net14717,
         net14718, net14719, net14720, net14721, net14722, net14723, net14724,
         net14725, net14726, net14727, net14728, net14729, net14730, net14731,
         net14732, net14733, net14734, net14735, net14736, net14737, net14738,
         net14739, net14740, net14741, net14742, net14743, net14744, net14745,
         net14746, net14747, net14748, net14749, net14750, net14751, net14752,
         net14753, net14754, net14755, net14756, net14757, net14758, net14759,
         net14760, net14761, net14762, net14763, net14764, net14765, net14766,
         net14767, net14768, net14769, net14770, net14771, net14772, net14773,
         net14774, net14775, net14776, net14777, net14778, net14779, net14780,
         net14781, net14782, net14783, net14784, net14785, net14786, net14787,
         net14788, net14789, net14790, net14791, net14792, net14793, net14794,
         net14795, net14796, net14797, net14798, net14799, net14800, net14801,
         net14802, net14803, net14804, net14805, net14806, net14807, net14808,
         net14809, net14810, net14811, net14812, net14813, net14814, net14815,
         net14816, net14817, net14818, net14819, net14820, net14821, net14822,
         net14823, net14824, net14825, net14826, net14827, net14828, net14829,
         net14830, net14831, net14832, net14833, net14834, net14835, net14836,
         net14837, net14838, net14839, net14840, net14841, net14842, net14843,
         net14844, net14845, net14846, net14847, net14848, net14849, net14850,
         net14851, net14852, net14853, net14854, net14855, net14856, net14857,
         net14858, net14859, net14860, net14861, net14862, net14863, net14864,
         net14865, net14866, net14867, net14868, net14869, net14870, net14871,
         net14872, net14873, net14874, net14875, net14876, net14877, net14878,
         net14879, net14880, net14881, net14882, net14883, net14884, net14885,
         net14886, net14887, net14888, net14889, net14890, net14891, net14892,
         net14893, net14894, net14895, net14896, net14897, net14898, net14899,
         net14900, net14901, net14902, net14903, net14904, net14905, net14906,
         net14907, net14908, net14909, net14910, net14911, net14912, net14913,
         net14914, net14915, net14916, net14917, net14918, net14919, net14920,
         net14921, net14922, net14923, net14924, net14925, net14926, net14927,
         net14928, net14929, net14930, net14931, net14932, net14933, net14934,
         net14935, net14936, net14937, net14938, net14939, net14940, net14941,
         net14942, net14943, net14944, net14945, net14946, net14947, net14948,
         net14949, net14950, net14951, net14952, net14953, net14954, net14955,
         net14956, net14957, net14958, net14959, net14960, net14961, net14962,
         net14963, net14964, net14965, net14966, net14967, net14968, net14969,
         net14970, net14971, net14972, net14973, net14974, net14975, net14976,
         net14977, net14978, net14979, net14980, net14981, net14982, net14983,
         net14984, net14985, net14986, net14987, net14988, net14989, net14990,
         net14991, net14992, net14993, net14994, net14995, net14996, net14997,
         net14998, net14999, net15000, net15001, net15002, net15003, net15004,
         net15005, net15006, net15007, net15008, net15009, net15010, net15011,
         net15012, net15013, net15014, net15015, net15016, net15017, net15018,
         net15019, net15020, net15021, net15022, net15023, net15024, net15025,
         net15026, net15027, net15028, net15029, net15030, net15031, net15032,
         net15033, net15034, net15035, net15036, net15037, net15038, net15039,
         net15040, net15041, net15042, net15043, net15044, net15045, net15046,
         net15047, net15048, net15049, net15050, net15051, net15052, net15053,
         net15054, net15055, net15056, net15057, net15058, net15059, net15060,
         net15061, net15062, net15063, net15064, net15065, net15066, net15067,
         net15068, net15069, net15070, net15071, net15072, net15073, net15074,
         net15075, net15076, net15077, net15078, net15079, net15080, net15081,
         net15082, net15083, net15084, net15085, net15086, net15087, net15088,
         net15089, net15090, net15091, net15092, net15093, net15094, net15095,
         net15096, net15097, net15098, net15099, net15100, net15101, net15102,
         net15103, net15104, net15105, net15106, net15107, net15108, net15109,
         net15110, net15111, net15112, net15113, net15114, net15115, net15116,
         net15117, net15118, net15119, net15120, net15121, net15122, net15123,
         net15124, net15125, net15126, net15127, net15128, net15129, net15130,
         net15131, net15132, net15133, net15134, net15135, net15136, net15137,
         net15138, net15139, net15140, net15141, net15142, net15143, net15144,
         net15145, net15146, net15147, net15148, net15149, net15150, net15151,
         net15152, net15153, net15154, net15155, net15156, net15157, net15158,
         net15159, net15160, net15161, net15162, net15163, net15164, net15165,
         net15166, net15167, net15168, net15169, net15170, net15171, net15172,
         net15173, net15174, net15175, net15176, net15177, net15178, net15179,
         net15180, net15181, net15182, net15183, net15184, net15185, net15186,
         net15187, net15188, net15189, net15190, net15191, net15192, net15193,
         net15194, net15195, net15196, net15197, net15198, net15199, net15200,
         net15201, net15202, net15203, net15204, net15205, net15206, net15207,
         net15208, net15209, net15210, net15211, net15212, net15213, net15214,
         net15215, net15216, net15217, net15218, net15219, net15220, net15221,
         net15222, net15223, net15224, net15225, net15226, net15227, net15228,
         net15229, net15230, net15231, net15232, net15233, net15234, net15235,
         net15236, net15237, net15238, net15239, net15240, net15241, net15242,
         net15243, net15244, net15245, net15246, net15247, net15248, net15249,
         net15250, net15251, net15252, net15253, net15254, net15255, net15256,
         net15257, net15258, net15259, net15260, net15261, net15262, net15263,
         net15264, net15265, net15266, net15267, net15268, net15269, net15270,
         net15271, net15272, net15273, net15274, net15275, net15276, net15277,
         net15278, net15279, net15280, net15281, net15282, net15283, net15284,
         net15285, net15286, net15287, net15288, net15289, net15290, net15291,
         net15292, net15293, net15294, net15295, net15296, net15297, net15298,
         net15299, net15300, net15301, net15302, net15303, net15304, net15305,
         net15306, net15307, net15308, net15309, net15310, net15311, net15312,
         net15313, net15314, net15315, net15316, net15317, net15318, net15319,
         net15320, net15321, net15322, net15323, net15324, net15325, net15326,
         net15327, net15328, net15329, net15330, net15331, net15332, net15333,
         net15334, net15335, net15336, net15337, net15338, net15339, net15340,
         net15341, net15342, net15343, net15344, net15345, net15346, net15347,
         net15348, net15349, net15350, net15351, net15352, net15353, net15354,
         net15355, net15356, net15357, net15358, net15359, net15360, net15361,
         net15362, net15363, net15364, net15365, net15366, net15367, net15368,
         net15369, net15370, net15371, net15372, net15373, net15374, net15375,
         net15376, net15377, net15378, net15379, net15380, net15381, net15382,
         net15383, net15384, net15385, net15386, net15387, net15388, net15389,
         net15390, net15391, net15392, net15393, net15394, net15395, net15396,
         net15397, net15398, net15399, net15400, net15401, net15402, net15403,
         net15404, net15405, net15406, net15407, net15408, net15409, net15410,
         net15411, net15412, net15413, net15414, net15415, net15416, net15417,
         net15418, net15419, net15420, net15421, net15422, net15423, net15424,
         net15425, net15426, net15427, net15428, net15429, net15430, net15431,
         net15432, net15433, net15434, net15435, net15436, net15437, net15438,
         net15439, net15440, net15441, net15442, net15443, net15444, net15445,
         net15446, net15447, net15448, net15449, net15450, net15451, net15452,
         net15453, net15454, net15455, net15456, net15457, net15458, net15459,
         net15460, net15461, net15462, net15463, net15464, net15465, net15466,
         net15467, net15468, net15469, net15470, net15471, net15472, net15473,
         net15474, net15475, net15476, net15477, net15478, net15479, net15480,
         net15481, net15482, net15483, net15484, net15485, net15486, net15487,
         net15488, net15489, net15490, net15491, net15492, net15493, net15494,
         net15495, net15496, net15497, net15498, net15499, net15500, net15501,
         net15502, net15503, net15504, net15505, net15506, net15507, net15508,
         net15509, net15510, net15511, net15512, net15513, net15514, net15515,
         net15516, net15517, net15518, net15519, net15520, net15521, net15522,
         net15523, net15524, net15525, net15526, net15527, net15528, net15529,
         net15530, net15531, net15532, net15533, net15534, net15535, net15536,
         net15537, net15538, net15539, net15540, net15541, net15542, net15543,
         net15544, net15545, net15546, net15547, net15548, net15549, net15550,
         net15551, net15552, net15553, net15554, net15555, net15556, net15557,
         net15558, net15559, net15560, net15561, net15562, net15563, net15564,
         net15565, net15566, net15567, net15568, net15569, net15570, net15571,
         net15572, net15573, net15574, net15575, net15576, net15577, net15578,
         net15579, net15580, net15581, net15582, net15583, net15584, net15585,
         net15586, net15587, net15588, net15589, net15590, net15591, net15592,
         net15593, net15594, net15595, net15596, net15597, net15598, net15599,
         net15600, net15601, net15602, net15603, net15604, net15605, net15606,
         net15607, net15608, net15609, net15610, net15611, net15612, net15613,
         net15614, net15615, net15616, net15617, net15618, net15619, net15620,
         net15621, net15622, net15623, net15624, net15625, net15626, net15627,
         net15628, net15629, net15630, net15631, net15632, net15633, net15634,
         net15635, net15636, net15637, net15638, net15639, net15640, net15641,
         net15642, net15643, net15644, net15645, net15646, net15647, net15648,
         net15649, net15650, net15651, net15652, net15653, net15654, net15655,
         net15656, net15657, net15658, net15659, net15660, net15661, net15662,
         net15663, net15664, net15665, net15666, net15667, net15668, net15669,
         net15670, net15671, net15672, net15673, net15674, net15675, net15676,
         net15677, net15678, net15679, net15680, net15681, net15682, net15683,
         net15684, net15685, net15686, net15687, net15688, net15689, net15690,
         net15691, net15692, net15693, net15694, net15695, net15696, net15697,
         net15698, net15699, net15700, net15701, net15702, net15703, net15704,
         net15705, net15706, net15707, net15708, net15709, net15710, net15711,
         net15712, net15713, net15714, net15715, net15716, net15717, net15718,
         net15719, net15720, net15721, net15722, net15723, net15724, net15725,
         net15726, net15727, net15728, net15729, net15730, net15731, net15732,
         net15733, net15734, net15735, net15736, net15737, net15738, net15739,
         net15740, net15741, net15742, net15743, net15744, net15745, net15746,
         net15747, net15748, net15749, net15750, net15751, net15752, net15753,
         net15754, net15755, net15756, net15757, net15758, net15759, net15760,
         net15761, net15762, net15763, net15764, net15765, net15766, net15767,
         net15768, net15769, net15770, net15771, net15772, net15773, net15774,
         net15775, net15776, net15777, net15778, net15779, net15780, net15781,
         net15782, net15783, net15784, net15785, net15786, net15787, net15788,
         net15789, net15790, net15791, net15792, net15793, net15794, net15795,
         net15796, net15797, net15798, net15799, net15800, net15801, net15802,
         net15803, net15804, net15805, net15806, net15807, net15808, net15809,
         net15810, net15811, net15812, net15813, net15814, net15815, net15816,
         net15817, net15818, net15819, net15820, net15821, net15822;
  wire   [62:0] a1stg_in1;
  wire   [54:0] a1stg_in1a;
  wire   [63:0] a1stg_in2;
  wire   [54:0] a1stg_in2a;
  wire   [63:11] a1stg_norm_frac1;
  wire   [63:0] a1stg_norm_frac2;
  wire   [63:0] a2stg_frac1_in;
  wire   [63:0] a2stg_frac1;
  wire   [63:0] a2stg_frac2_in;
  wire   [62:0] a2stg_frac2;
  wire   [63:0] a2stg_frac2a;
  wire   [3:0] a2stg_shr_cnt_5;
  wire   [3:0] a2stg_shr_cnt_5_inv;
  wire   [63:0] a2stg_shr_tmp2;
  wire   [4:0] a2stg_shr_cnt_4;
  wire   [63:0] a2stg_shr_tmp4;
  wire   [4:0] a2stg_shr_cnt_3;
  wire   [63:0] a2stg_shr_tmp6;
  wire   [1:0] a2stg_shr_cnt_2;
  wire   [63:0] a2stg_shr_tmp8;
  wire   [1:0] a2stg_shr_cnt_1;
  wire   [63:0] a2stg_shr_tmp10;
  wire   [1:0] a2stg_shr_cnt_0;
  wire   [115:52] a2stg_shr;
  wire   [27:12] a2stg_shr_tmp18;
  wire   [5:0] a2stg_shr_cnt;
  wire   [63:20] a2stg_nx_neq0_84_tmp_1;
  wire   [63:36] a2stg_nx_neq0_84_tmp_2;
  wire   [63:44] a2stg_nx_neq0_84_tmp_3;
  wire   [63:57] a2stg_nx_neq0_84_tmp_4;
  wire   [61:59] a2stg_nx_neq0_84_tmp_5;
  wire   [60:59] a2stg_nx_neq0_84_tmp_6;
  wire   [63:0] a3stg_frac2;
  wire   [63:0] a2stg_shr_frac2_inv;
  wire   [63:0] a3stg_frac2_in;
  wire   [63:0] a3stg_frac1;
  wire   [63:0] a2stg_fracadd_in2;
  wire   [63:0] a2stg_fracadd;
  wire   [63:0] a3stg_ld0_frac;
  wire   [53:0] a2stg_expdec_tmp;
  wire   [53:0] a2stg_expdec;
  wire   [53:0] a3stg_expdec;
  wire   [63:0] a3stg_fracadd;
  wire   [3:3] astg_xtra_regs;
  wire   [5:3] a2stg_shr_cnta;
  wire   [2:0] a4stg_shl_cnt_dec54_0;
  wire   [2:0] a4stg_shl_cnt_dec54_1;
  wire   [2:0] a4stg_shl_cnt_dec54_2;
  wire   [2:0] a4stg_shl_cnt_dec54_3;
  wire   [2:0] a2stg_shr_cnta_5;
  wire   [63:2] a4stg_rnd_frac_pre1_in;
  wire   [63:0] a4stg_rnd_frac_pre1;
  wire   [63:1] a4stg_rnd_frac_pre3_in;
  wire   [63:0] a4stg_rnd_frac_pre3;
  wire   [63:0] a4stg_shl;
  wire   [38:12] a4stg_rnd_frac;
  wire   [63:0] a4stg_rnd_frac_pre2_in;
  wire   [63:0] a4stg_rnd_frac_pre2;
  wire   [63:0] a4stg_shl_data_in;
  wire   [63:0] a4stg_shl_data;
  wire   [51:0] a4stg_rndadd_tmp;
  wire   [63:0] a4stg_shl_tmp4;
  wire   [51:0] a5stg_rndadd;
  wire   [63:0] a5stg_rnd_frac;
  wire   [63:0] a5stg_shl;

  clken_buf ckbuf_add_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fadd_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE63 i_a1stg_in1 ( .din(inq_in1), .en(a1stg_step), .clk(clk), .q(
        a1stg_in1), .se(se), .si({net15760, net15761, net15762, net15763, 
        net15764, net15765, net15766, net15767, net15768, net15769, net15770, 
        net15771, net15772, net15773, net15774, net15775, net15776, net15777, 
        net15778, net15779, net15780, net15781, net15782, net15783, net15784, 
        net15785, net15786, net15787, net15788, net15789, net15790, net15791, 
        net15792, net15793, net15794, net15795, net15796, net15797, net15798, 
        net15799, net15800, net15801, net15802, net15803, net15804, net15805, 
        net15806, net15807, net15808, net15809, net15810, net15811, net15812, 
        net15813, net15814, net15815, net15816, net15817, net15818, net15819, 
        net15820, net15821, net15822}) );
  dffe_SIZE55 i_a1stg_in1a ( .din(inq_in1[54:0]), .en(a1stg_step), .clk(clk), 
        .q(a1stg_in1a), .se(se), .si({net15705, net15706, net15707, net15708, 
        net15709, net15710, net15711, net15712, net15713, net15714, net15715, 
        net15716, net15717, net15718, net15719, net15720, net15721, net15722, 
        net15723, net15724, net15725, net15726, net15727, net15728, net15729, 
        net15730, net15731, net15732, net15733, net15734, net15735, net15736, 
        net15737, net15738, net15739, net15740, net15741, net15742, net15743, 
        net15744, net15745, net15746, net15747, net15748, net15749, net15750, 
        net15751, net15752, net15753, net15754, net15755, net15756, net15757, 
        net15758, net15759}) );
  dffe_SIZE64 i_a1stg_in2 ( .din(inq_in2), .en(a1stg_step), .clk(clk), .q(
        a1stg_in2), .se(se), .si({net15641, net15642, net15643, net15644, 
        net15645, net15646, net15647, net15648, net15649, net15650, net15651, 
        net15652, net15653, net15654, net15655, net15656, net15657, net15658, 
        net15659, net15660, net15661, net15662, net15663, net15664, net15665, 
        net15666, net15667, net15668, net15669, net15670, net15671, net15672, 
        net15673, net15674, net15675, net15676, net15677, net15678, net15679, 
        net15680, net15681, net15682, net15683, net15684, net15685, net15686, 
        net15687, net15688, net15689, net15690, net15691, net15692, net15693, 
        net15694, net15695, net15696, net15697, net15698, net15699, net15700, 
        net15701, net15702, net15703, net15704}) );
  dffe_SIZE55 i_a1stg_in2a ( .din(inq_in2[54:0]), .en(a1stg_step), .clk(clk), 
        .q(a1stg_in2a), .se(se), .si({net15586, net15587, net15588, net15589, 
        net15590, net15591, net15592, net15593, net15594, net15595, net15596, 
        net15597, net15598, net15599, net15600, net15601, net15602, net15603, 
        net15604, net15605, net15606, net15607, net15608, net15609, net15610, 
        net15611, net15612, net15613, net15614, net15615, net15616, net15617, 
        net15618, net15619, net15620, net15621, net15622, net15623, net15624, 
        net15625, net15626, net15627, net15628, net15629, net15630, net15631, 
        net15632, net15633, net15634, net15635, net15636, net15637, net15638, 
        net15639, net15640}) );
  fpu_in2_gt_in1_frac i_a1stg_in2_gt_in1_frac ( .din1(a1stg_in1a), .din2(
        a1stg_in2a), .sngop(a1stg_sngop), .expadd11(a1stg_expadd3_11), .expeq(
        a1stg_in2_eq_in1_exp), .din2_neq_din1(a1stg_in2_neq_in1_frac), 
        .din2_gt_din1(a1stg_in2_gt_in1_frac), .din2_gt1_din1(a1stg_in2_gt_in1)
         );
  dffe_SIZE64 i_a2stg_frac1 ( .din(a2stg_frac1_in), .en(a6stg_step), .clk(clk), 
        .q(a2stg_frac1), .se(se), .si({net15522, net15523, net15524, net15525, 
        net15526, net15527, net15528, net15529, net15530, net15531, net15532, 
        net15533, net15534, net15535, net15536, net15537, net15538, net15539, 
        net15540, net15541, net15542, net15543, net15544, net15545, net15546, 
        net15547, net15548, net15549, net15550, net15551, net15552, net15553, 
        net15554, net15555, net15556, net15557, net15558, net15559, net15560, 
        net15561, net15562, net15563, net15564, net15565, net15566, net15567, 
        net15568, net15569, net15570, net15571, net15572, net15573, net15574, 
        net15575, net15576, net15577, net15578, net15579, net15580, net15581, 
        net15582, net15583, net15584, net15585}) );
  dffe_SIZE64 i_a2stg_frac2 ( .din(a2stg_frac2_in), .en(a6stg_step), .clk(clk), 
        .q({a2stg_frac2_63, a2stg_frac2}), .se(se), .si({net15458, net15459, 
        net15460, net15461, net15462, net15463, net15464, net15465, net15466, 
        net15467, net15468, net15469, net15470, net15471, net15472, net15473, 
        net15474, net15475, net15476, net15477, net15478, net15479, net15480, 
        net15481, net15482, net15483, net15484, net15485, net15486, net15487, 
        net15488, net15489, net15490, net15491, net15492, net15493, net15494, 
        net15495, net15496, net15497, net15498, net15499, net15500, net15501, 
        net15502, net15503, net15504, net15505, net15506, net15507, net15508, 
        net15509, net15510, net15511, net15512, net15513, net15514, net15515, 
        net15516, net15517, net15518, net15519, net15520, net15521}) );
  dffe_SIZE64 i_a2stg_frac2a ( .din(a2stg_frac2_in), .en(a6stg_step), .clk(clk), .q(a2stg_frac2a), .se(se), .si({net15394, net15395, net15396, net15397, 
        net15398, net15399, net15400, net15401, net15402, net15403, net15404, 
        net15405, net15406, net15407, net15408, net15409, net15410, net15411, 
        net15412, net15413, net15414, net15415, net15416, net15417, net15418, 
        net15419, net15420, net15421, net15422, net15423, net15424, net15425, 
        net15426, net15427, net15428, net15429, net15430, net15431, net15432, 
        net15433, net15434, net15435, net15436, net15437, net15438, net15439, 
        net15440, net15441, net15442, net15443, net15444, net15445, net15446, 
        net15447, net15448, net15449, net15450, net15451, net15452, net15453, 
        net15454, net15455, net15456, net15457}) );
  dff_SIZE64 i_a3stg_frac2 ( .din(a3stg_frac2_in), .clk(clk), .q(a3stg_frac2), 
        .se(se), .si({net15330, net15331, net15332, net15333, net15334, 
        net15335, net15336, net15337, net15338, net15339, net15340, net15341, 
        net15342, net15343, net15344, net15345, net15346, net15347, net15348, 
        net15349, net15350, net15351, net15352, net15353, net15354, net15355, 
        net15356, net15357, net15358, net15359, net15360, net15361, net15362, 
        net15363, net15364, net15365, net15366, net15367, net15368, net15369, 
        net15370, net15371, net15372, net15373, net15374, net15375, net15376, 
        net15377, net15378, net15379, net15380, net15381, net15382, net15383, 
        net15384, net15385, net15386, net15387, net15388, net15389, net15390, 
        net15391, net15392, net15393}) );
  dffe_SIZE64 i_a3stg_frac1 ( .din({1'b0, a2stg_frac1[63:1]}), .en(a6stg_step), 
        .clk(clk), .q(a3stg_frac1), .se(se), .si({net15266, net15267, net15268, 
        net15269, net15270, net15271, net15272, net15273, net15274, net15275, 
        net15276, net15277, net15278, net15279, net15280, net15281, net15282, 
        net15283, net15284, net15285, net15286, net15287, net15288, net15289, 
        net15290, net15291, net15292, net15293, net15294, net15295, net15296, 
        net15297, net15298, net15299, net15300, net15301, net15302, net15303, 
        net15304, net15305, net15306, net15307, net15308, net15309, net15310, 
        net15311, net15312, net15313, net15314, net15315, net15316, net15317, 
        net15318, net15319, net15320, net15321, net15322, net15323, net15324, 
        net15325, net15326, net15327, net15328, net15329}) );
  dffe_SIZE64 i_a3stg_ld0_frac ( .din(a2stg_fracadd), .en(a6stg_step), .clk(
        clk), .q(a3stg_ld0_frac), .se(se), .si({net15202, net15203, net15204, 
        net15205, net15206, net15207, net15208, net15209, net15210, net15211, 
        net15212, net15213, net15214, net15215, net15216, net15217, net15218, 
        net15219, net15220, net15221, net15222, net15223, net15224, net15225, 
        net15226, net15227, net15228, net15229, net15230, net15231, net15232, 
        net15233, net15234, net15235, net15236, net15237, net15238, net15239, 
        net15240, net15241, net15242, net15243, net15244, net15245, net15246, 
        net15247, net15248, net15249, net15250, net15251, net15252, net15253, 
        net15254, net15255, net15256, net15257, net15258, net15259, net15260, 
        net15261, net15262, net15263, net15264, net15265}) );
  ASHR_UNS_UNS_OP srl_705 ( .A({1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SH(
        a2stg_exp), .Z(a2stg_expdec_tmp) );
  dffe_SIZE54 i_a3stg_expdec ( .din(a2stg_expdec), .en(a6stg_step), .clk(clk), 
        .q(a3stg_expdec), .se(se), .si({net15148, net15149, net15150, net15151, 
        net15152, net15153, net15154, net15155, net15156, net15157, net15158, 
        net15159, net15160, net15161, net15162, net15163, net15164, net15165, 
        net15166, net15167, net15168, net15169, net15170, net15171, net15172, 
        net15173, net15174, net15175, net15176, net15177, net15178, net15179, 
        net15180, net15181, net15182, net15183, net15184, net15185, net15186, 
        net15187, net15188, net15189, net15190, net15191, net15192, net15193, 
        net15194, net15195, net15196, net15197, net15198, net15199, net15200, 
        net15201}) );
  fpu_denorm_frac i_a3stg_denorm ( .din1({a3stg_ld0_frac[63:11], 
        a3stg_ld0_dnrm_10}), .din2(a3stg_expdec), .din2_din1_denorm(
        a3stg_denorm), .din2_din1_denorm_inv(a3stg_denorm_inv), 
        .din2_din1_denorma(a3stg_denorma), .din2_din1_denorm_inva(
        a3stg_denorm_inva) );
  fpu_cnt_lead0_64b i_a3stg_lead0 ( .din(a3stg_ld0_frac), .lead0(a3stg_lead0)
         );
  dffe_SIZE64 i_astg_xtra_regs ( .din({a2stg_shr_cnt_5_inv_in, 
        a2stg_shr_cnt_5_inv_in, a2stg_shr_cnt_5_inv_in, a2stg_shr_cnt_5_inv_in, 
        a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], 
        a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5:3], a2stg_shr_cnt_in[4], 
        a2stg_shr_cnt_in[4], a2stg_shr_cnt_in[4], a2stg_shr_cnt_in[4], 
        a2stg_shr_cnt_in[4:3], a2stg_shr_cnt_in[3], a2stg_shr_cnt_in[3], 
        a2stg_shr_cnt_in[3], a2stg_shr_cnt_in[3], a2stg_shr_cnt_in, 
        a4stg_round_in, a2stg_shr_cnt_in[2], a2stg_shr_cnt_in[2:1], 
        a2stg_shr_cnt_in[1:0], a2stg_shr_cnt_in[0], a4stg_shl_cnt_in[6], 
        a4stg_shl_cnt_in[6], a4stg_shl_cnt_in[6], a4stg_shl_cnt_in[7], 
        a4stg_shl_cnt_in[7], a4stg_shl_cnt_in[7], a4stg_shl_cnt_in[8], 
        a4stg_shl_cnt_in[8], a4stg_shl_cnt_in[8], a4stg_shl_cnt_in[9], 
        a4stg_shl_cnt_in[9], a4stg_shl_cnt_in[9], a4stg_shl_cnt_in[5:0], 
        a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], a2stg_shr_cnt_in[5], 
        a2stg_fracadd_frac2_inv_in, a2stg_fracadd_frac2_inv_shr1_in, 
        a3stg_denorm_inva, a2stg_fsdtoix_nx, a2stg_fsdtoi_nx, 1'b0, 
        a2stg_fracadd_cin_in, a3stg_sub_in, a3stg_sub_in}), .en(a6stg_step), 
        .clk(clk), .q({a2stg_shr_cnt_5_inv, a2stg_shr_cnt_5, a2stg_shr_cnta, 
        a2stg_shr_cnt_4, a2stg_shr_cnt_3, a2stg_shr_cnt, a4stg_round, 
        a2stg_shr_cnt_2, a2stg_shr_cnt_1, a2stg_shr_cnt_0, 
        a4stg_shl_cnt_dec54_0, a4stg_shl_cnt_dec54_1, a4stg_shl_cnt_dec54_2, 
        a4stg_shl_cnt_dec54_3, a4stg_shl_cnt, a2stg_shr_cnta_5, 
        a2stg_fracadd_frac2_inv, a2stg_fracadd_frac2_inv_shr1, 
        a4stg_denorm_inv, a3stg_fsdtoix_nx, a3stg_fsdtoi_nx, astg_xtra_regs[3], 
        a2stg_fracadd_cin, a3stg_sub, a3stg_suba}), .se(se), .si({net15084, 
        net15085, net15086, net15087, net15088, net15089, net15090, net15091, 
        net15092, net15093, net15094, net15095, net15096, net15097, net15098, 
        net15099, net15100, net15101, net15102, net15103, net15104, net15105, 
        net15106, net15107, net15108, net15109, net15110, net15111, net15112, 
        net15113, net15114, net15115, net15116, net15117, net15118, net15119, 
        net15120, net15121, net15122, net15123, net15124, net15125, net15126, 
        net15127, net15128, net15129, net15130, net15131, net15132, net15133, 
        net15134, net15135, net15136, net15137, net15138, net15139, net15140, 
        net15141, net15142, net15143, net15144, net15145, net15146, net15147})
         );
  dff_SIZE64 i_a4stg_rnd_frac_pre1 ( .din({a4stg_rnd_frac_pre1_in, 1'b0, 1'b0}), .clk(clk), .q(a4stg_rnd_frac_pre1), .se(se), .si({net15020, net15021, 
        net15022, net15023, net15024, net15025, net15026, net15027, net15028, 
        net15029, net15030, net15031, net15032, net15033, net15034, net15035, 
        net15036, net15037, net15038, net15039, net15040, net15041, net15042, 
        net15043, net15044, net15045, net15046, net15047, net15048, net15049, 
        net15050, net15051, net15052, net15053, net15054, net15055, net15056, 
        net15057, net15058, net15059, net15060, net15061, net15062, net15063, 
        net15064, net15065, net15066, net15067, net15068, net15069, net15070, 
        net15071, net15072, net15073, net15074, net15075, net15076, net15077, 
        net15078, net15079, net15080, net15081, net15082, net15083}) );
  dff_SIZE64 i_a4stg_rnd_frac_pre3 ( .din({a4stg_rnd_frac_pre3_in, 1'b0}), 
        .clk(clk), .q(a4stg_rnd_frac_pre3), .se(se), .si({net14956, net14957, 
        net14958, net14959, net14960, net14961, net14962, net14963, net14964, 
        net14965, net14966, net14967, net14968, net14969, net14970, net14971, 
        net14972, net14973, net14974, net14975, net14976, net14977, net14978, 
        net14979, net14980, net14981, net14982, net14983, net14984, net14985, 
        net14986, net14987, net14988, net14989, net14990, net14991, net14992, 
        net14993, net14994, net14995, net14996, net14997, net14998, net14999, 
        net15000, net15001, net15002, net15003, net15004, net15005, net15006, 
        net15007, net15008, net15009, net15010, net15011, net15012, net15013, 
        net15014, net15015, net15016, net15017, net15018, net15019}) );
  dff_SIZE64 i_a4stg_rnd_frac_pre2 ( .din(a4stg_rnd_frac_pre2_in), .clk(clk), 
        .q(a4stg_rnd_frac_pre2), .se(se), .si({net14892, net14893, net14894, 
        net14895, net14896, net14897, net14898, net14899, net14900, net14901, 
        net14902, net14903, net14904, net14905, net14906, net14907, net14908, 
        net14909, net14910, net14911, net14912, net14913, net14914, net14915, 
        net14916, net14917, net14918, net14919, net14920, net14921, net14922, 
        net14923, net14924, net14925, net14926, net14927, net14928, net14929, 
        net14930, net14931, net14932, net14933, net14934, net14935, net14936, 
        net14937, net14938, net14939, net14940, net14941, net14942, net14943, 
        net14944, net14945, net14946, net14947, net14948, net14949, net14950, 
        net14951, net14952, net14953, net14954, net14955}) );
  dffe_SIZE64 i_a4stg_shl_data ( .din(a4stg_shl_data_in), .en(a6stg_step), 
        .clk(clk), .q(a4stg_shl_data), .se(se), .si({net14828, net14829, 
        net14830, net14831, net14832, net14833, net14834, net14835, net14836, 
        net14837, net14838, net14839, net14840, net14841, net14842, net14843, 
        net14844, net14845, net14846, net14847, net14848, net14849, net14850, 
        net14851, net14852, net14853, net14854, net14855, net14856, net14857, 
        net14858, net14859, net14860, net14861, net14862, net14863, net14864, 
        net14865, net14866, net14867, net14868, net14869, net14870, net14871, 
        net14872, net14873, net14874, net14875, net14876, net14877, net14878, 
        net14879, net14880, net14881, net14882, net14883, net14884, net14885, 
        net14886, net14887, net14888, net14889, net14890, net14891}) );
  ASH_UNS_UNS_OP sll_979 ( .A(a4stg_shl_tmp4), .SH(a4stg_shl_cnt[3:0]), .Z(
        a4stg_shl) );
  dffe_SIZE58 i_a5stg_rndadd ( .din({a4stg_rndadd_cout, add_frac_out_rndadd, 
        add_frac_out_rnd_frac, a4stg_in_of, add_frac_out_shl, a4stg_to_0, 
        a4stg_rndadd_tmp}), .en(a6stg_step), .clk(clk), .q({add_of_out_cout, 
        a5stg_frac_out_rndadd, a5stg_frac_out_rnd_frac, a5stg_in_of, 
        a5stg_frac_out_shl, a5stg_to_0, a5stg_rndadd}), .se(se), .si({net14770, 
        net14771, net14772, net14773, net14774, net14775, net14776, net14777, 
        net14778, net14779, net14780, net14781, net14782, net14783, net14784, 
        net14785, net14786, net14787, net14788, net14789, net14790, net14791, 
        net14792, net14793, net14794, net14795, net14796, net14797, net14798, 
        net14799, net14800, net14801, net14802, net14803, net14804, net14805, 
        net14806, net14807, net14808, net14809, net14810, net14811, net14812, 
        net14813, net14814, net14815, net14816, net14817, net14818, net14819, 
        net14820, net14821, net14822, net14823, net14824, net14825, net14826, 
        net14827}) );
  dffe_SIZE64 i_a5stg_rnd_frac ( .din({a4stg_rnd_frac_63, a4stg_rnd_frac_62, 
        a4stg_rnd_frac_61, a4stg_rnd_frac_60, a4stg_rnd_frac_59, 
        a4stg_rnd_frac_58, a4stg_rnd_frac_57, a4stg_rnd_frac_56, 
        a4stg_rnd_frac_55, a4stg_rnd_frac_54, a4stg_rnd_frac_53, 
        a4stg_rnd_frac_52, a4stg_rnd_frac_51, a4stg_rnd_frac_50, 
        a4stg_rnd_frac_49, a4stg_rnd_frac_48, a4stg_rnd_frac_47, 
        a4stg_rnd_frac_46, a4stg_rnd_frac_45, a4stg_rnd_frac_44, 
        a4stg_rnd_frac_43, a4stg_rnd_frac_42, a4stg_rnd_frac_41, 
        a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac, 
        a4stg_rnd_frac_11, a4stg_rnd_frac_10, a4stg_rnd_frac_9, 
        a4stg_rnd_frac_8, a4stg_rnd_frac_7, a4stg_rnd_frac_6, a4stg_rnd_frac_5, 
        a4stg_rnd_frac_4, a4stg_rnd_frac_3, a4stg_rnd_frac_2, a4stg_rnd_frac_1, 
        a4stg_rnd_frac_0}), .en(a6stg_step), .clk(clk), .q(a5stg_rnd_frac), 
        .se(se), .si({net14706, net14707, net14708, net14709, net14710, 
        net14711, net14712, net14713, net14714, net14715, net14716, net14717, 
        net14718, net14719, net14720, net14721, net14722, net14723, net14724, 
        net14725, net14726, net14727, net14728, net14729, net14730, net14731, 
        net14732, net14733, net14734, net14735, net14736, net14737, net14738, 
        net14739, net14740, net14741, net14742, net14743, net14744, net14745, 
        net14746, net14747, net14748, net14749, net14750, net14751, net14752, 
        net14753, net14754, net14755, net14756, net14757, net14758, net14759, 
        net14760, net14761, net14762, net14763, net14764, net14765, net14766, 
        net14767, net14768, net14769}) );
  dffe_SIZE64 i_a5stg_shl ( .din(a4stg_shl), .en(a6stg_step), .clk(clk), .q(
        a5stg_shl), .se(se), .si({net14642, net14643, net14644, net14645, 
        net14646, net14647, net14648, net14649, net14650, net14651, net14652, 
        net14653, net14654, net14655, net14656, net14657, net14658, net14659, 
        net14660, net14661, net14662, net14663, net14664, net14665, net14666, 
        net14667, net14668, net14669, net14670, net14671, net14672, net14673, 
        net14674, net14675, net14676, net14677, net14678, net14679, net14680, 
        net14681, net14682, net14683, net14684, net14685, net14686, net14687, 
        net14688, net14689, net14690, net14691, net14692, net14693, net14694, 
        net14695, net14696, net14697, net14698, net14699, net14700, net14701, 
        net14702, net14703, net14704, net14705}) );
  ADD_UNS_OP add_767 ( .A(a3stg_frac1), .B(a3stg_frac2), .Z({N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66}) );
  ADD_UNS_OP add_679 ( .A(a2stg_frac1), .B(a2stg_fracadd_in2), .Z({N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, N4, N3, N2}) );
  ADD_UNS_OP add_956 ( .A({a4stg_rnd_frac_62, a4stg_rnd_frac_61, 
        a4stg_rnd_frac_60, a4stg_rnd_frac_59, a4stg_rnd_frac_58, 
        a4stg_rnd_frac_57, a4stg_rnd_frac_56, a4stg_rnd_frac_55, 
        a4stg_rnd_frac_54, a4stg_rnd_frac_53, a4stg_rnd_frac_52, 
        a4stg_rnd_frac_51, a4stg_rnd_frac_50, a4stg_rnd_frac_49, 
        a4stg_rnd_frac_48, a4stg_rnd_frac_47, a4stg_rnd_frac_46, 
        a4stg_rnd_frac_45, a4stg_rnd_frac_44, a4stg_rnd_frac_43, 
        a4stg_rnd_frac_42, a4stg_rnd_frac_41, a4stg_rnd_frac_40, 
        a4stg_rnd_frac_39, a4stg_rnd_frac, a4stg_rnd_frac_11}), .B({
        a4stg_rnd_sng, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, a4stg_rnd_dbl}), .Z({
        a4stg_rndadd_cout, a4stg_rndadd_tmp}) );
  ADD_UNS_OP add_767_2 ( .A({N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66}), .B(a3stg_suba), .Z(a3stg_fracadd) );
  ADD_UNS_OP add_679_2 ( .A({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2}), .B(
        a2stg_fracadd_cin), .Z(a2stg_fracadd) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_AND2 C1540 ( .A(N161), .B(N164), .Z(a1stg_in2_eq_in1_exp) );
  GTECH_AND2 C1541 ( .A(N157), .B(N160), .Z(N161) );
  GTECH_AND2 C1542 ( .A(N153), .B(N156), .Z(N157) );
  GTECH_AND2 C1543 ( .A(N150), .B(N152), .Z(N153) );
  GTECH_AND2 C1544 ( .A(N147), .B(N149), .Z(N150) );
  GTECH_AND2 C1545 ( .A(N144), .B(N146), .Z(N147) );
  GTECH_AND2 C1546 ( .A(N141), .B(N143), .Z(N144) );
  GTECH_AND2 C1547 ( .A(N138), .B(N140), .Z(N141) );
  GTECH_AND2 C1548 ( .A(N135), .B(N137), .Z(N138) );
  GTECH_AND2 C1549 ( .A(N132), .B(N134), .Z(N135) );
  GTECH_NOT I_1 ( .A(N131), .Z(N132) );
  GTECH_XOR2 C1551 ( .A(a1stg_in1[62]), .B(a1stg_in2[62]), .Z(N131) );
  GTECH_NOT I_2 ( .A(N133), .Z(N134) );
  GTECH_XOR2 C1553 ( .A(a1stg_in1[61]), .B(a1stg_in2[61]), .Z(N133) );
  GTECH_NOT I_3 ( .A(N136), .Z(N137) );
  GTECH_XOR2 C1555 ( .A(a1stg_in1[60]), .B(a1stg_in2[60]), .Z(N136) );
  GTECH_NOT I_4 ( .A(N139), .Z(N140) );
  GTECH_XOR2 C1557 ( .A(a1stg_in1[59]), .B(a1stg_in2[59]), .Z(N139) );
  GTECH_NOT I_5 ( .A(N142), .Z(N143) );
  GTECH_XOR2 C1559 ( .A(a1stg_in1[58]), .B(a1stg_in2[58]), .Z(N142) );
  GTECH_NOT I_6 ( .A(N145), .Z(N146) );
  GTECH_XOR2 C1561 ( .A(a1stg_in1[57]), .B(a1stg_in2[57]), .Z(N145) );
  GTECH_NOT I_7 ( .A(N148), .Z(N149) );
  GTECH_XOR2 C1563 ( .A(a1stg_in1[56]), .B(a1stg_in2[56]), .Z(N148) );
  GTECH_NOT I_8 ( .A(N151), .Z(N152) );
  GTECH_XOR2 C1565 ( .A(a1stg_in1[55]), .B(a1stg_in2[55]), .Z(N151) );
  GTECH_OR2 C1566 ( .A(N155), .B(a1stg_sngop), .Z(N156) );
  GTECH_NOT I_9 ( .A(N154), .Z(N155) );
  GTECH_XOR2 C1568 ( .A(a1stg_in1[54]), .B(a1stg_in2[54]), .Z(N154) );
  GTECH_OR2 C1569 ( .A(N159), .B(a1stg_sngop), .Z(N160) );
  GTECH_NOT I_10 ( .A(N158), .Z(N159) );
  GTECH_XOR2 C1571 ( .A(a1stg_in1[53]), .B(a1stg_in2[53]), .Z(N158) );
  GTECH_OR2 C1572 ( .A(N163), .B(a1stg_sngop), .Z(N164) );
  GTECH_NOT I_11 ( .A(N162), .Z(N163) );
  GTECH_XOR2 C1574 ( .A(a1stg_in1[52]), .B(a1stg_in2[52]), .Z(N162) );
  GTECH_OR2 C1575 ( .A(N167), .B(N168), .Z(a1stg_norm_frac1[63]) );
  GTECH_OR2 C1576 ( .A(N166), .B(a1stg_norm_sng_in1), .Z(N167) );
  GTECH_OR2 C1577 ( .A(a1stg_norm_dbl_in1), .B(N165), .Z(N166) );
  GTECH_AND2 C1578 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[51]), .Z(N165) );
  GTECH_AND2 C1579 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[54]), .Z(N168) );
  GTECH_OR2 C1580 ( .A(N173), .B(N174), .Z(a1stg_norm_frac1[62]) );
  GTECH_OR2 C1581 ( .A(N171), .B(N172), .Z(N173) );
  GTECH_OR2 C1582 ( .A(N169), .B(N170), .Z(N171) );
  GTECH_AND2 C1583 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[51]), .Z(N169) );
  GTECH_AND2 C1584 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[50]), .Z(N170) );
  GTECH_AND2 C1585 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[54]), .Z(N172) );
  GTECH_AND2 C1586 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[53]), .Z(N174) );
  GTECH_OR2 C1587 ( .A(N179), .B(N180), .Z(a1stg_norm_frac1[61]) );
  GTECH_OR2 C1588 ( .A(N177), .B(N178), .Z(N179) );
  GTECH_OR2 C1589 ( .A(N175), .B(N176), .Z(N177) );
  GTECH_AND2 C1590 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[50]), .Z(N175) );
  GTECH_AND2 C1591 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[49]), .Z(N176) );
  GTECH_AND2 C1592 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[53]), .Z(N178) );
  GTECH_AND2 C1593 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[52]), .Z(N180) );
  GTECH_OR2 C1594 ( .A(N185), .B(N186), .Z(a1stg_norm_frac1[60]) );
  GTECH_OR2 C1595 ( .A(N183), .B(N184), .Z(N185) );
  GTECH_OR2 C1596 ( .A(N181), .B(N182), .Z(N183) );
  GTECH_AND2 C1597 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[49]), .Z(N181) );
  GTECH_AND2 C1598 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[48]), .Z(N182) );
  GTECH_AND2 C1599 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[52]), .Z(N184) );
  GTECH_AND2 C1600 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[51]), .Z(N186) );
  GTECH_OR2 C1601 ( .A(N191), .B(N192), .Z(a1stg_norm_frac1[59]) );
  GTECH_OR2 C1602 ( .A(N189), .B(N190), .Z(N191) );
  GTECH_OR2 C1603 ( .A(N187), .B(N188), .Z(N189) );
  GTECH_AND2 C1604 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[48]), .Z(N187) );
  GTECH_AND2 C1605 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[47]), .Z(N188) );
  GTECH_AND2 C1606 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[51]), .Z(N190) );
  GTECH_AND2 C1607 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[50]), .Z(N192) );
  GTECH_OR2 C1608 ( .A(N197), .B(N198), .Z(a1stg_norm_frac1[58]) );
  GTECH_OR2 C1609 ( .A(N195), .B(N196), .Z(N197) );
  GTECH_OR2 C1610 ( .A(N193), .B(N194), .Z(N195) );
  GTECH_AND2 C1611 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[47]), .Z(N193) );
  GTECH_AND2 C1612 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[46]), .Z(N194) );
  GTECH_AND2 C1613 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[50]), .Z(N196) );
  GTECH_AND2 C1614 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[49]), .Z(N198) );
  GTECH_OR2 C1615 ( .A(N203), .B(N204), .Z(a1stg_norm_frac1[57]) );
  GTECH_OR2 C1616 ( .A(N201), .B(N202), .Z(N203) );
  GTECH_OR2 C1617 ( .A(N199), .B(N200), .Z(N201) );
  GTECH_AND2 C1618 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[46]), .Z(N199) );
  GTECH_AND2 C1619 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[45]), .Z(N200) );
  GTECH_AND2 C1620 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[49]), .Z(N202) );
  GTECH_AND2 C1621 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[48]), .Z(N204) );
  GTECH_OR2 C1622 ( .A(N209), .B(N210), .Z(a1stg_norm_frac1[56]) );
  GTECH_OR2 C1623 ( .A(N207), .B(N208), .Z(N209) );
  GTECH_OR2 C1624 ( .A(N205), .B(N206), .Z(N207) );
  GTECH_AND2 C1625 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[45]), .Z(N205) );
  GTECH_AND2 C1626 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[44]), .Z(N206) );
  GTECH_AND2 C1627 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[48]), .Z(N208) );
  GTECH_AND2 C1628 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[47]), .Z(N210) );
  GTECH_OR2 C1629 ( .A(N215), .B(N216), .Z(a1stg_norm_frac1[55]) );
  GTECH_OR2 C1630 ( .A(N213), .B(N214), .Z(N215) );
  GTECH_OR2 C1631 ( .A(N211), .B(N212), .Z(N213) );
  GTECH_AND2 C1632 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[44]), .Z(N211) );
  GTECH_AND2 C1633 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[43]), .Z(N212) );
  GTECH_AND2 C1634 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[47]), .Z(N214) );
  GTECH_AND2 C1635 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[46]), .Z(N216) );
  GTECH_OR2 C1636 ( .A(N221), .B(N222), .Z(a1stg_norm_frac1[54]) );
  GTECH_OR2 C1637 ( .A(N219), .B(N220), .Z(N221) );
  GTECH_OR2 C1638 ( .A(N217), .B(N218), .Z(N219) );
  GTECH_AND2 C1639 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[43]), .Z(N217) );
  GTECH_AND2 C1640 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[42]), .Z(N218) );
  GTECH_AND2 C1641 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[46]), .Z(N220) );
  GTECH_AND2 C1642 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[45]), .Z(N222) );
  GTECH_OR2 C1643 ( .A(N227), .B(N228), .Z(a1stg_norm_frac1[53]) );
  GTECH_OR2 C1644 ( .A(N225), .B(N226), .Z(N227) );
  GTECH_OR2 C1645 ( .A(N223), .B(N224), .Z(N225) );
  GTECH_AND2 C1646 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[42]), .Z(N223) );
  GTECH_AND2 C1647 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[41]), .Z(N224) );
  GTECH_AND2 C1648 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[45]), .Z(N226) );
  GTECH_AND2 C1649 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[44]), .Z(N228) );
  GTECH_OR2 C1650 ( .A(N233), .B(N234), .Z(a1stg_norm_frac1[52]) );
  GTECH_OR2 C1651 ( .A(N231), .B(N232), .Z(N233) );
  GTECH_OR2 C1652 ( .A(N229), .B(N230), .Z(N231) );
  GTECH_AND2 C1653 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[41]), .Z(N229) );
  GTECH_AND2 C1654 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[40]), .Z(N230) );
  GTECH_AND2 C1655 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[44]), .Z(N232) );
  GTECH_AND2 C1656 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[43]), .Z(N234) );
  GTECH_OR2 C1657 ( .A(N239), .B(N240), .Z(a1stg_norm_frac1[51]) );
  GTECH_OR2 C1658 ( .A(N237), .B(N238), .Z(N239) );
  GTECH_OR2 C1659 ( .A(N235), .B(N236), .Z(N237) );
  GTECH_AND2 C1660 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[40]), .Z(N235) );
  GTECH_AND2 C1661 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[39]), .Z(N236) );
  GTECH_AND2 C1662 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[43]), .Z(N238) );
  GTECH_AND2 C1663 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[42]), .Z(N240) );
  GTECH_OR2 C1664 ( .A(N245), .B(N246), .Z(a1stg_norm_frac1[50]) );
  GTECH_OR2 C1665 ( .A(N243), .B(N244), .Z(N245) );
  GTECH_OR2 C1666 ( .A(N241), .B(N242), .Z(N243) );
  GTECH_AND2 C1667 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[39]), .Z(N241) );
  GTECH_AND2 C1668 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[38]), .Z(N242) );
  GTECH_AND2 C1669 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[42]), .Z(N244) );
  GTECH_AND2 C1670 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[41]), .Z(N246) );
  GTECH_OR2 C1671 ( .A(N251), .B(N252), .Z(a1stg_norm_frac1[49]) );
  GTECH_OR2 C1672 ( .A(N249), .B(N250), .Z(N251) );
  GTECH_OR2 C1673 ( .A(N247), .B(N248), .Z(N249) );
  GTECH_AND2 C1674 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[38]), .Z(N247) );
  GTECH_AND2 C1675 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[37]), .Z(N248) );
  GTECH_AND2 C1676 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[41]), .Z(N250) );
  GTECH_AND2 C1677 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[40]), .Z(N252) );
  GTECH_OR2 C1678 ( .A(N257), .B(N258), .Z(a1stg_norm_frac1[48]) );
  GTECH_OR2 C1679 ( .A(N255), .B(N256), .Z(N257) );
  GTECH_OR2 C1680 ( .A(N253), .B(N254), .Z(N255) );
  GTECH_AND2 C1681 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[37]), .Z(N253) );
  GTECH_AND2 C1682 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[36]), .Z(N254) );
  GTECH_AND2 C1683 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[40]), .Z(N256) );
  GTECH_AND2 C1684 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[39]), .Z(N258) );
  GTECH_OR2 C1685 ( .A(N263), .B(N264), .Z(a1stg_norm_frac1[47]) );
  GTECH_OR2 C1686 ( .A(N261), .B(N262), .Z(N263) );
  GTECH_OR2 C1687 ( .A(N259), .B(N260), .Z(N261) );
  GTECH_AND2 C1688 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[36]), .Z(N259) );
  GTECH_AND2 C1689 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[35]), .Z(N260) );
  GTECH_AND2 C1690 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[39]), .Z(N262) );
  GTECH_AND2 C1691 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[38]), .Z(N264) );
  GTECH_OR2 C1692 ( .A(N269), .B(N270), .Z(a1stg_norm_frac1[46]) );
  GTECH_OR2 C1693 ( .A(N267), .B(N268), .Z(N269) );
  GTECH_OR2 C1694 ( .A(N265), .B(N266), .Z(N267) );
  GTECH_AND2 C1695 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[35]), .Z(N265) );
  GTECH_AND2 C1696 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[34]), .Z(N266) );
  GTECH_AND2 C1697 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[38]), .Z(N268) );
  GTECH_AND2 C1698 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[37]), .Z(N270) );
  GTECH_OR2 C1699 ( .A(N275), .B(N276), .Z(a1stg_norm_frac1[45]) );
  GTECH_OR2 C1700 ( .A(N273), .B(N274), .Z(N275) );
  GTECH_OR2 C1701 ( .A(N271), .B(N272), .Z(N273) );
  GTECH_AND2 C1702 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[34]), .Z(N271) );
  GTECH_AND2 C1703 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[33]), .Z(N272) );
  GTECH_AND2 C1704 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[37]), .Z(N274) );
  GTECH_AND2 C1705 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[36]), .Z(N276) );
  GTECH_OR2 C1706 ( .A(N281), .B(N282), .Z(a1stg_norm_frac1[44]) );
  GTECH_OR2 C1707 ( .A(N279), .B(N280), .Z(N281) );
  GTECH_OR2 C1708 ( .A(N277), .B(N278), .Z(N279) );
  GTECH_AND2 C1709 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[33]), .Z(N277) );
  GTECH_AND2 C1710 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[32]), .Z(N278) );
  GTECH_AND2 C1711 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[36]), .Z(N280) );
  GTECH_AND2 C1712 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[35]), .Z(N282) );
  GTECH_OR2 C1713 ( .A(N287), .B(N288), .Z(a1stg_norm_frac1[43]) );
  GTECH_OR2 C1714 ( .A(N285), .B(N286), .Z(N287) );
  GTECH_OR2 C1715 ( .A(N283), .B(N284), .Z(N285) );
  GTECH_AND2 C1716 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[32]), .Z(N283) );
  GTECH_AND2 C1717 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[31]), .Z(N284) );
  GTECH_AND2 C1718 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[35]), .Z(N286) );
  GTECH_AND2 C1719 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[34]), .Z(N288) );
  GTECH_OR2 C1720 ( .A(N293), .B(N294), .Z(a1stg_norm_frac1[42]) );
  GTECH_OR2 C1721 ( .A(N291), .B(N292), .Z(N293) );
  GTECH_OR2 C1722 ( .A(N289), .B(N290), .Z(N291) );
  GTECH_AND2 C1723 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[31]), .Z(N289) );
  GTECH_AND2 C1724 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[30]), .Z(N290) );
  GTECH_AND2 C1725 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[34]), .Z(N292) );
  GTECH_AND2 C1726 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[33]), .Z(N294) );
  GTECH_OR2 C1727 ( .A(N299), .B(N300), .Z(a1stg_norm_frac1[41]) );
  GTECH_OR2 C1728 ( .A(N297), .B(N298), .Z(N299) );
  GTECH_OR2 C1729 ( .A(N295), .B(N296), .Z(N297) );
  GTECH_AND2 C1730 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[30]), .Z(N295) );
  GTECH_AND2 C1731 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[29]), .Z(N296) );
  GTECH_AND2 C1732 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[33]), .Z(N298) );
  GTECH_AND2 C1733 ( .A(a1stg_denorm_sng_in1), .B(a1stg_in1[32]), .Z(N300) );
  GTECH_OR2 C1734 ( .A(N303), .B(N304), .Z(a1stg_norm_frac1[40]) );
  GTECH_OR2 C1735 ( .A(N301), .B(N302), .Z(N303) );
  GTECH_AND2 C1736 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[29]), .Z(N301) );
  GTECH_AND2 C1737 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[28]), .Z(N302) );
  GTECH_AND2 C1738 ( .A(a1stg_norm_sng_in1), .B(a1stg_in1[32]), .Z(N304) );
  GTECH_OR2 C1739 ( .A(N305), .B(N306), .Z(a1stg_norm_frac1[39]) );
  GTECH_AND2 C1740 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[28]), .Z(N305) );
  GTECH_AND2 C1741 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[27]), .Z(N306) );
  GTECH_OR2 C1742 ( .A(N307), .B(N308), .Z(a1stg_norm_frac1[38]) );
  GTECH_AND2 C1743 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[27]), .Z(N307) );
  GTECH_AND2 C1744 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[26]), .Z(N308) );
  GTECH_OR2 C1745 ( .A(N309), .B(N310), .Z(a1stg_norm_frac1[37]) );
  GTECH_AND2 C1746 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[26]), .Z(N309) );
  GTECH_AND2 C1747 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[25]), .Z(N310) );
  GTECH_OR2 C1748 ( .A(N311), .B(N312), .Z(a1stg_norm_frac1[36]) );
  GTECH_AND2 C1749 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[25]), .Z(N311) );
  GTECH_AND2 C1750 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[24]), .Z(N312) );
  GTECH_OR2 C1751 ( .A(N313), .B(N314), .Z(a1stg_norm_frac1[35]) );
  GTECH_AND2 C1752 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[24]), .Z(N313) );
  GTECH_AND2 C1753 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[23]), .Z(N314) );
  GTECH_OR2 C1754 ( .A(N315), .B(N316), .Z(a1stg_norm_frac1[34]) );
  GTECH_AND2 C1755 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[23]), .Z(N315) );
  GTECH_AND2 C1756 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[22]), .Z(N316) );
  GTECH_OR2 C1757 ( .A(N317), .B(N318), .Z(a1stg_norm_frac1[33]) );
  GTECH_AND2 C1758 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[22]), .Z(N317) );
  GTECH_AND2 C1759 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[21]), .Z(N318) );
  GTECH_OR2 C1760 ( .A(N319), .B(N320), .Z(a1stg_norm_frac1[32]) );
  GTECH_AND2 C1761 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[21]), .Z(N319) );
  GTECH_AND2 C1762 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[20]), .Z(N320) );
  GTECH_OR2 C1763 ( .A(N321), .B(N322), .Z(a1stg_norm_frac1[31]) );
  GTECH_AND2 C1764 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[20]), .Z(N321) );
  GTECH_AND2 C1765 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[19]), .Z(N322) );
  GTECH_OR2 C1766 ( .A(N323), .B(N324), .Z(a1stg_norm_frac1[30]) );
  GTECH_AND2 C1767 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[19]), .Z(N323) );
  GTECH_AND2 C1768 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[18]), .Z(N324) );
  GTECH_OR2 C1769 ( .A(N325), .B(N326), .Z(a1stg_norm_frac1[29]) );
  GTECH_AND2 C1770 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[18]), .Z(N325) );
  GTECH_AND2 C1771 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[17]), .Z(N326) );
  GTECH_OR2 C1772 ( .A(N327), .B(N328), .Z(a1stg_norm_frac1[28]) );
  GTECH_AND2 C1773 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[17]), .Z(N327) );
  GTECH_AND2 C1774 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[16]), .Z(N328) );
  GTECH_OR2 C1775 ( .A(N329), .B(N330), .Z(a1stg_norm_frac1[27]) );
  GTECH_AND2 C1776 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[16]), .Z(N329) );
  GTECH_AND2 C1777 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[15]), .Z(N330) );
  GTECH_OR2 C1778 ( .A(N331), .B(N332), .Z(a1stg_norm_frac1[26]) );
  GTECH_AND2 C1779 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[15]), .Z(N331) );
  GTECH_AND2 C1780 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[14]), .Z(N332) );
  GTECH_OR2 C1781 ( .A(N333), .B(N334), .Z(a1stg_norm_frac1[25]) );
  GTECH_AND2 C1782 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[14]), .Z(N333) );
  GTECH_AND2 C1783 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[13]), .Z(N334) );
  GTECH_OR2 C1784 ( .A(N335), .B(N336), .Z(a1stg_norm_frac1[24]) );
  GTECH_AND2 C1785 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[13]), .Z(N335) );
  GTECH_AND2 C1786 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[12]), .Z(N336) );
  GTECH_OR2 C1787 ( .A(N337), .B(N338), .Z(a1stg_norm_frac1[23]) );
  GTECH_AND2 C1788 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[12]), .Z(N337) );
  GTECH_AND2 C1789 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[11]), .Z(N338) );
  GTECH_OR2 C1790 ( .A(N339), .B(N340), .Z(a1stg_norm_frac1[22]) );
  GTECH_AND2 C1791 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[11]), .Z(N339) );
  GTECH_AND2 C1792 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[10]), .Z(N340) );
  GTECH_OR2 C1793 ( .A(N341), .B(N342), .Z(a1stg_norm_frac1[21]) );
  GTECH_AND2 C1794 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[10]), .Z(N341) );
  GTECH_AND2 C1795 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[9]), .Z(N342) );
  GTECH_OR2 C1796 ( .A(N343), .B(N344), .Z(a1stg_norm_frac1[20]) );
  GTECH_AND2 C1797 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[9]), .Z(N343) );
  GTECH_AND2 C1798 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[8]), .Z(N344) );
  GTECH_OR2 C1799 ( .A(N345), .B(N346), .Z(a1stg_norm_frac1[19]) );
  GTECH_AND2 C1800 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[8]), .Z(N345) );
  GTECH_AND2 C1801 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[7]), .Z(N346) );
  GTECH_OR2 C1802 ( .A(N347), .B(N348), .Z(a1stg_norm_frac1[18]) );
  GTECH_AND2 C1803 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[7]), .Z(N347) );
  GTECH_AND2 C1804 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[6]), .Z(N348) );
  GTECH_OR2 C1805 ( .A(N349), .B(N350), .Z(a1stg_norm_frac1[17]) );
  GTECH_AND2 C1806 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[6]), .Z(N349) );
  GTECH_AND2 C1807 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[5]), .Z(N350) );
  GTECH_OR2 C1808 ( .A(N351), .B(N352), .Z(a1stg_norm_frac1[16]) );
  GTECH_AND2 C1809 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[5]), .Z(N351) );
  GTECH_AND2 C1810 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[4]), .Z(N352) );
  GTECH_OR2 C1811 ( .A(N353), .B(N354), .Z(a1stg_norm_frac1[15]) );
  GTECH_AND2 C1812 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[4]), .Z(N353) );
  GTECH_AND2 C1813 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[3]), .Z(N354) );
  GTECH_OR2 C1814 ( .A(N355), .B(N356), .Z(a1stg_norm_frac1[14]) );
  GTECH_AND2 C1815 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[3]), .Z(N355) );
  GTECH_AND2 C1816 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[2]), .Z(N356) );
  GTECH_OR2 C1817 ( .A(N357), .B(N358), .Z(a1stg_norm_frac1[13]) );
  GTECH_AND2 C1818 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[2]), .Z(N357) );
  GTECH_AND2 C1819 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[1]), .Z(N358) );
  GTECH_OR2 C1820 ( .A(N359), .B(N360), .Z(a1stg_norm_frac1[12]) );
  GTECH_AND2 C1821 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[1]), .Z(N359) );
  GTECH_AND2 C1822 ( .A(a1stg_denorm_dbl_in1), .B(a1stg_in1[0]), .Z(N360) );
  GTECH_AND2 C1823 ( .A(a1stg_norm_dbl_in1), .B(a1stg_in1[0]), .Z(
        a1stg_norm_frac1[11]) );
  GTECH_OR2 C1824 ( .A(N365), .B(N366), .Z(a1stg_norm_frac2[63]) );
  GTECH_OR2 C1825 ( .A(N363), .B(N364), .Z(N365) );
  GTECH_OR2 C1826 ( .A(N362), .B(a1stg_norm_sng_in2), .Z(N363) );
  GTECH_OR2 C1827 ( .A(a1stg_norm_dbl_in2), .B(N361), .Z(N362) );
  GTECH_AND2 C1828 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[51]), .Z(N361) );
  GTECH_AND2 C1829 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[54]), .Z(N364) );
  GTECH_AND2 C1830 ( .A(a1stg_intlngop), .B(a1stg_in2[63]), .Z(N366) );
  GTECH_OR2 C1831 ( .A(N373), .B(N374), .Z(a1stg_norm_frac2[62]) );
  GTECH_OR2 C1832 ( .A(N371), .B(N372), .Z(N373) );
  GTECH_OR2 C1833 ( .A(N369), .B(N370), .Z(N371) );
  GTECH_OR2 C1834 ( .A(N367), .B(N368), .Z(N369) );
  GTECH_AND2 C1835 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[51]), .Z(N367) );
  GTECH_AND2 C1836 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[50]), .Z(N368) );
  GTECH_AND2 C1837 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[54]), .Z(N370) );
  GTECH_AND2 C1838 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[53]), .Z(N372) );
  GTECH_AND2 C1839 ( .A(a1stg_intlngop), .B(a1stg_in2[62]), .Z(N374) );
  GTECH_OR2 C1840 ( .A(N381), .B(N382), .Z(a1stg_norm_frac2[61]) );
  GTECH_OR2 C1841 ( .A(N379), .B(N380), .Z(N381) );
  GTECH_OR2 C1842 ( .A(N377), .B(N378), .Z(N379) );
  GTECH_OR2 C1843 ( .A(N375), .B(N376), .Z(N377) );
  GTECH_AND2 C1844 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[50]), .Z(N375) );
  GTECH_AND2 C1845 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[49]), .Z(N376) );
  GTECH_AND2 C1846 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[53]), .Z(N378) );
  GTECH_AND2 C1847 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[52]), .Z(N380) );
  GTECH_AND2 C1848 ( .A(a1stg_intlngop), .B(a1stg_in2[61]), .Z(N382) );
  GTECH_OR2 C1849 ( .A(N389), .B(N390), .Z(a1stg_norm_frac2[60]) );
  GTECH_OR2 C1850 ( .A(N387), .B(N388), .Z(N389) );
  GTECH_OR2 C1851 ( .A(N385), .B(N386), .Z(N387) );
  GTECH_OR2 C1852 ( .A(N383), .B(N384), .Z(N385) );
  GTECH_AND2 C1853 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[49]), .Z(N383) );
  GTECH_AND2 C1854 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[48]), .Z(N384) );
  GTECH_AND2 C1855 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[52]), .Z(N386) );
  GTECH_AND2 C1856 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[51]), .Z(N388) );
  GTECH_AND2 C1857 ( .A(a1stg_intlngop), .B(a1stg_in2[60]), .Z(N390) );
  GTECH_OR2 C1858 ( .A(N397), .B(N398), .Z(a1stg_norm_frac2[59]) );
  GTECH_OR2 C1859 ( .A(N395), .B(N396), .Z(N397) );
  GTECH_OR2 C1860 ( .A(N393), .B(N394), .Z(N395) );
  GTECH_OR2 C1861 ( .A(N391), .B(N392), .Z(N393) );
  GTECH_AND2 C1862 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[48]), .Z(N391) );
  GTECH_AND2 C1863 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[47]), .Z(N392) );
  GTECH_AND2 C1864 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[51]), .Z(N394) );
  GTECH_AND2 C1865 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[50]), .Z(N396) );
  GTECH_AND2 C1866 ( .A(a1stg_intlngop), .B(a1stg_in2[59]), .Z(N398) );
  GTECH_OR2 C1867 ( .A(N405), .B(N406), .Z(a1stg_norm_frac2[58]) );
  GTECH_OR2 C1868 ( .A(N403), .B(N404), .Z(N405) );
  GTECH_OR2 C1869 ( .A(N401), .B(N402), .Z(N403) );
  GTECH_OR2 C1870 ( .A(N399), .B(N400), .Z(N401) );
  GTECH_AND2 C1871 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[47]), .Z(N399) );
  GTECH_AND2 C1872 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[46]), .Z(N400) );
  GTECH_AND2 C1873 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[50]), .Z(N402) );
  GTECH_AND2 C1874 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[49]), .Z(N404) );
  GTECH_AND2 C1875 ( .A(a1stg_intlngop), .B(a1stg_in2[58]), .Z(N406) );
  GTECH_OR2 C1876 ( .A(N413), .B(N414), .Z(a1stg_norm_frac2[57]) );
  GTECH_OR2 C1877 ( .A(N411), .B(N412), .Z(N413) );
  GTECH_OR2 C1878 ( .A(N409), .B(N410), .Z(N411) );
  GTECH_OR2 C1879 ( .A(N407), .B(N408), .Z(N409) );
  GTECH_AND2 C1880 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[46]), .Z(N407) );
  GTECH_AND2 C1881 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[45]), .Z(N408) );
  GTECH_AND2 C1882 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[49]), .Z(N410) );
  GTECH_AND2 C1883 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[48]), .Z(N412) );
  GTECH_AND2 C1884 ( .A(a1stg_intlngop), .B(a1stg_in2[57]), .Z(N414) );
  GTECH_OR2 C1885 ( .A(N421), .B(N422), .Z(a1stg_norm_frac2[56]) );
  GTECH_OR2 C1886 ( .A(N419), .B(N420), .Z(N421) );
  GTECH_OR2 C1887 ( .A(N417), .B(N418), .Z(N419) );
  GTECH_OR2 C1888 ( .A(N415), .B(N416), .Z(N417) );
  GTECH_AND2 C1889 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[45]), .Z(N415) );
  GTECH_AND2 C1890 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[44]), .Z(N416) );
  GTECH_AND2 C1891 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[48]), .Z(N418) );
  GTECH_AND2 C1892 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[47]), .Z(N420) );
  GTECH_AND2 C1893 ( .A(a1stg_intlngop), .B(a1stg_in2[56]), .Z(N422) );
  GTECH_OR2 C1894 ( .A(N429), .B(N430), .Z(a1stg_norm_frac2[55]) );
  GTECH_OR2 C1895 ( .A(N427), .B(N428), .Z(N429) );
  GTECH_OR2 C1896 ( .A(N425), .B(N426), .Z(N427) );
  GTECH_OR2 C1897 ( .A(N423), .B(N424), .Z(N425) );
  GTECH_AND2 C1898 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[44]), .Z(N423) );
  GTECH_AND2 C1899 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[43]), .Z(N424) );
  GTECH_AND2 C1900 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[47]), .Z(N426) );
  GTECH_AND2 C1901 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[46]), .Z(N428) );
  GTECH_AND2 C1902 ( .A(a1stg_intlngop), .B(a1stg_in2[55]), .Z(N430) );
  GTECH_OR2 C1903 ( .A(N437), .B(N438), .Z(a1stg_norm_frac2[54]) );
  GTECH_OR2 C1904 ( .A(N435), .B(N436), .Z(N437) );
  GTECH_OR2 C1905 ( .A(N433), .B(N434), .Z(N435) );
  GTECH_OR2 C1906 ( .A(N431), .B(N432), .Z(N433) );
  GTECH_AND2 C1907 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[43]), .Z(N431) );
  GTECH_AND2 C1908 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[42]), .Z(N432) );
  GTECH_AND2 C1909 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[46]), .Z(N434) );
  GTECH_AND2 C1910 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[45]), .Z(N436) );
  GTECH_AND2 C1911 ( .A(a1stg_intlngop), .B(a1stg_in2[54]), .Z(N438) );
  GTECH_OR2 C1912 ( .A(N445), .B(N446), .Z(a1stg_norm_frac2[53]) );
  GTECH_OR2 C1913 ( .A(N443), .B(N444), .Z(N445) );
  GTECH_OR2 C1914 ( .A(N441), .B(N442), .Z(N443) );
  GTECH_OR2 C1915 ( .A(N439), .B(N440), .Z(N441) );
  GTECH_AND2 C1916 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[42]), .Z(N439) );
  GTECH_AND2 C1917 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[41]), .Z(N440) );
  GTECH_AND2 C1918 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[45]), .Z(N442) );
  GTECH_AND2 C1919 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[44]), .Z(N444) );
  GTECH_AND2 C1920 ( .A(a1stg_intlngop), .B(a1stg_in2[53]), .Z(N446) );
  GTECH_OR2 C1921 ( .A(N453), .B(N454), .Z(a1stg_norm_frac2[52]) );
  GTECH_OR2 C1922 ( .A(N451), .B(N452), .Z(N453) );
  GTECH_OR2 C1923 ( .A(N449), .B(N450), .Z(N451) );
  GTECH_OR2 C1924 ( .A(N447), .B(N448), .Z(N449) );
  GTECH_AND2 C1925 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[41]), .Z(N447) );
  GTECH_AND2 C1926 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[40]), .Z(N448) );
  GTECH_AND2 C1927 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[44]), .Z(N450) );
  GTECH_AND2 C1928 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[43]), .Z(N452) );
  GTECH_AND2 C1929 ( .A(a1stg_intlngop), .B(a1stg_in2[52]), .Z(N454) );
  GTECH_OR2 C1930 ( .A(N461), .B(N462), .Z(a1stg_norm_frac2[51]) );
  GTECH_OR2 C1931 ( .A(N459), .B(N460), .Z(N461) );
  GTECH_OR2 C1932 ( .A(N457), .B(N458), .Z(N459) );
  GTECH_OR2 C1933 ( .A(N455), .B(N456), .Z(N457) );
  GTECH_AND2 C1934 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[40]), .Z(N455) );
  GTECH_AND2 C1935 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[39]), .Z(N456) );
  GTECH_AND2 C1936 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[43]), .Z(N458) );
  GTECH_AND2 C1937 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[42]), .Z(N460) );
  GTECH_AND2 C1938 ( .A(a1stg_intlngop), .B(a1stg_in2[51]), .Z(N462) );
  GTECH_OR2 C1939 ( .A(N469), .B(N470), .Z(a1stg_norm_frac2[50]) );
  GTECH_OR2 C1940 ( .A(N467), .B(N468), .Z(N469) );
  GTECH_OR2 C1941 ( .A(N465), .B(N466), .Z(N467) );
  GTECH_OR2 C1942 ( .A(N463), .B(N464), .Z(N465) );
  GTECH_AND2 C1943 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[39]), .Z(N463) );
  GTECH_AND2 C1944 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[38]), .Z(N464) );
  GTECH_AND2 C1945 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[42]), .Z(N466) );
  GTECH_AND2 C1946 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[41]), .Z(N468) );
  GTECH_AND2 C1947 ( .A(a1stg_intlngop), .B(a1stg_in2[50]), .Z(N470) );
  GTECH_OR2 C1948 ( .A(N477), .B(N478), .Z(a1stg_norm_frac2[49]) );
  GTECH_OR2 C1949 ( .A(N475), .B(N476), .Z(N477) );
  GTECH_OR2 C1950 ( .A(N473), .B(N474), .Z(N475) );
  GTECH_OR2 C1951 ( .A(N471), .B(N472), .Z(N473) );
  GTECH_AND2 C1952 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[38]), .Z(N471) );
  GTECH_AND2 C1953 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[37]), .Z(N472) );
  GTECH_AND2 C1954 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[41]), .Z(N474) );
  GTECH_AND2 C1955 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[40]), .Z(N476) );
  GTECH_AND2 C1956 ( .A(a1stg_intlngop), .B(a1stg_in2[49]), .Z(N478) );
  GTECH_OR2 C1957 ( .A(N485), .B(N486), .Z(a1stg_norm_frac2[48]) );
  GTECH_OR2 C1958 ( .A(N483), .B(N484), .Z(N485) );
  GTECH_OR2 C1959 ( .A(N481), .B(N482), .Z(N483) );
  GTECH_OR2 C1960 ( .A(N479), .B(N480), .Z(N481) );
  GTECH_AND2 C1961 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[37]), .Z(N479) );
  GTECH_AND2 C1962 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[36]), .Z(N480) );
  GTECH_AND2 C1963 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[40]), .Z(N482) );
  GTECH_AND2 C1964 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[39]), .Z(N484) );
  GTECH_AND2 C1965 ( .A(a1stg_intlngop), .B(a1stg_in2[48]), .Z(N486) );
  GTECH_OR2 C1966 ( .A(N493), .B(N494), .Z(a1stg_norm_frac2[47]) );
  GTECH_OR2 C1967 ( .A(N491), .B(N492), .Z(N493) );
  GTECH_OR2 C1968 ( .A(N489), .B(N490), .Z(N491) );
  GTECH_OR2 C1969 ( .A(N487), .B(N488), .Z(N489) );
  GTECH_AND2 C1970 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[36]), .Z(N487) );
  GTECH_AND2 C1971 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[35]), .Z(N488) );
  GTECH_AND2 C1972 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[39]), .Z(N490) );
  GTECH_AND2 C1973 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[38]), .Z(N492) );
  GTECH_AND2 C1974 ( .A(a1stg_intlngop), .B(a1stg_in2[47]), .Z(N494) );
  GTECH_OR2 C1975 ( .A(N501), .B(N502), .Z(a1stg_norm_frac2[46]) );
  GTECH_OR2 C1976 ( .A(N499), .B(N500), .Z(N501) );
  GTECH_OR2 C1977 ( .A(N497), .B(N498), .Z(N499) );
  GTECH_OR2 C1978 ( .A(N495), .B(N496), .Z(N497) );
  GTECH_AND2 C1979 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[35]), .Z(N495) );
  GTECH_AND2 C1980 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[34]), .Z(N496) );
  GTECH_AND2 C1981 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[38]), .Z(N498) );
  GTECH_AND2 C1982 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[37]), .Z(N500) );
  GTECH_AND2 C1983 ( .A(a1stg_intlngop), .B(a1stg_in2[46]), .Z(N502) );
  GTECH_OR2 C1984 ( .A(N509), .B(N510), .Z(a1stg_norm_frac2[45]) );
  GTECH_OR2 C1985 ( .A(N507), .B(N508), .Z(N509) );
  GTECH_OR2 C1986 ( .A(N505), .B(N506), .Z(N507) );
  GTECH_OR2 C1987 ( .A(N503), .B(N504), .Z(N505) );
  GTECH_AND2 C1988 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[34]), .Z(N503) );
  GTECH_AND2 C1989 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[33]), .Z(N504) );
  GTECH_AND2 C1990 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[37]), .Z(N506) );
  GTECH_AND2 C1991 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[36]), .Z(N508) );
  GTECH_AND2 C1992 ( .A(a1stg_intlngop), .B(a1stg_in2[45]), .Z(N510) );
  GTECH_OR2 C1993 ( .A(N517), .B(N518), .Z(a1stg_norm_frac2[44]) );
  GTECH_OR2 C1994 ( .A(N515), .B(N516), .Z(N517) );
  GTECH_OR2 C1995 ( .A(N513), .B(N514), .Z(N515) );
  GTECH_OR2 C1996 ( .A(N511), .B(N512), .Z(N513) );
  GTECH_AND2 C1997 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[33]), .Z(N511) );
  GTECH_AND2 C1998 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[32]), .Z(N512) );
  GTECH_AND2 C1999 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[36]), .Z(N514) );
  GTECH_AND2 C2000 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[35]), .Z(N516) );
  GTECH_AND2 C2001 ( .A(a1stg_intlngop), .B(a1stg_in2[44]), .Z(N518) );
  GTECH_OR2 C2002 ( .A(N525), .B(N526), .Z(a1stg_norm_frac2[43]) );
  GTECH_OR2 C2003 ( .A(N523), .B(N524), .Z(N525) );
  GTECH_OR2 C2004 ( .A(N521), .B(N522), .Z(N523) );
  GTECH_OR2 C2005 ( .A(N519), .B(N520), .Z(N521) );
  GTECH_AND2 C2006 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[32]), .Z(N519) );
  GTECH_AND2 C2007 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[31]), .Z(N520) );
  GTECH_AND2 C2008 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[35]), .Z(N522) );
  GTECH_AND2 C2009 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[34]), .Z(N524) );
  GTECH_AND2 C2010 ( .A(a1stg_intlngop), .B(a1stg_in2[43]), .Z(N526) );
  GTECH_OR2 C2011 ( .A(N533), .B(N534), .Z(a1stg_norm_frac2[42]) );
  GTECH_OR2 C2012 ( .A(N531), .B(N532), .Z(N533) );
  GTECH_OR2 C2013 ( .A(N529), .B(N530), .Z(N531) );
  GTECH_OR2 C2014 ( .A(N527), .B(N528), .Z(N529) );
  GTECH_AND2 C2015 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[31]), .Z(N527) );
  GTECH_AND2 C2016 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[30]), .Z(N528) );
  GTECH_AND2 C2017 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[34]), .Z(N530) );
  GTECH_AND2 C2018 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[33]), .Z(N532) );
  GTECH_AND2 C2019 ( .A(a1stg_intlngop), .B(a1stg_in2[42]), .Z(N534) );
  GTECH_OR2 C2020 ( .A(N541), .B(N542), .Z(a1stg_norm_frac2[41]) );
  GTECH_OR2 C2021 ( .A(N539), .B(N540), .Z(N541) );
  GTECH_OR2 C2022 ( .A(N537), .B(N538), .Z(N539) );
  GTECH_OR2 C2023 ( .A(N535), .B(N536), .Z(N537) );
  GTECH_AND2 C2024 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[30]), .Z(N535) );
  GTECH_AND2 C2025 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[29]), .Z(N536) );
  GTECH_AND2 C2026 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[33]), .Z(N538) );
  GTECH_AND2 C2027 ( .A(a1stg_denorm_sng_in2), .B(a1stg_in2[32]), .Z(N540) );
  GTECH_AND2 C2028 ( .A(a1stg_intlngop), .B(a1stg_in2[41]), .Z(N542) );
  GTECH_OR2 C2029 ( .A(N547), .B(N548), .Z(a1stg_norm_frac2[40]) );
  GTECH_OR2 C2030 ( .A(N545), .B(N546), .Z(N547) );
  GTECH_OR2 C2031 ( .A(N543), .B(N544), .Z(N545) );
  GTECH_AND2 C2032 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[29]), .Z(N543) );
  GTECH_AND2 C2033 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[28]), .Z(N544) );
  GTECH_AND2 C2034 ( .A(a1stg_norm_sng_in2), .B(a1stg_in2[32]), .Z(N546) );
  GTECH_AND2 C2035 ( .A(a1stg_intlngop), .B(a1stg_in2[40]), .Z(N548) );
  GTECH_OR2 C2036 ( .A(N551), .B(N552), .Z(a1stg_norm_frac2[39]) );
  GTECH_OR2 C2037 ( .A(N549), .B(N550), .Z(N551) );
  GTECH_AND2 C2038 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[28]), .Z(N549) );
  GTECH_AND2 C2039 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[27]), .Z(N550) );
  GTECH_AND2 C2040 ( .A(a1stg_intlngop), .B(a1stg_in2[39]), .Z(N552) );
  GTECH_OR2 C2041 ( .A(N555), .B(N556), .Z(a1stg_norm_frac2[38]) );
  GTECH_OR2 C2042 ( .A(N553), .B(N554), .Z(N555) );
  GTECH_AND2 C2043 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[27]), .Z(N553) );
  GTECH_AND2 C2044 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[26]), .Z(N554) );
  GTECH_AND2 C2045 ( .A(a1stg_intlngop), .B(a1stg_in2[38]), .Z(N556) );
  GTECH_OR2 C2046 ( .A(N559), .B(N560), .Z(a1stg_norm_frac2[37]) );
  GTECH_OR2 C2047 ( .A(N557), .B(N558), .Z(N559) );
  GTECH_AND2 C2048 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[26]), .Z(N557) );
  GTECH_AND2 C2049 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[25]), .Z(N558) );
  GTECH_AND2 C2050 ( .A(a1stg_intlngop), .B(a1stg_in2[37]), .Z(N560) );
  GTECH_OR2 C2051 ( .A(N563), .B(N564), .Z(a1stg_norm_frac2[36]) );
  GTECH_OR2 C2052 ( .A(N561), .B(N562), .Z(N563) );
  GTECH_AND2 C2053 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[25]), .Z(N561) );
  GTECH_AND2 C2054 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[24]), .Z(N562) );
  GTECH_AND2 C2055 ( .A(a1stg_intlngop), .B(a1stg_in2[36]), .Z(N564) );
  GTECH_OR2 C2056 ( .A(N567), .B(N568), .Z(a1stg_norm_frac2[35]) );
  GTECH_OR2 C2057 ( .A(N565), .B(N566), .Z(N567) );
  GTECH_AND2 C2058 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[24]), .Z(N565) );
  GTECH_AND2 C2059 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[23]), .Z(N566) );
  GTECH_AND2 C2060 ( .A(a1stg_intlngop), .B(a1stg_in2[35]), .Z(N568) );
  GTECH_OR2 C2061 ( .A(N571), .B(N572), .Z(a1stg_norm_frac2[34]) );
  GTECH_OR2 C2062 ( .A(N569), .B(N570), .Z(N571) );
  GTECH_AND2 C2063 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[23]), .Z(N569) );
  GTECH_AND2 C2064 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[22]), .Z(N570) );
  GTECH_AND2 C2065 ( .A(a1stg_intlngop), .B(a1stg_in2[34]), .Z(N572) );
  GTECH_OR2 C2066 ( .A(N575), .B(N576), .Z(a1stg_norm_frac2[33]) );
  GTECH_OR2 C2067 ( .A(N573), .B(N574), .Z(N575) );
  GTECH_AND2 C2068 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[22]), .Z(N573) );
  GTECH_AND2 C2069 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[21]), .Z(N574) );
  GTECH_AND2 C2070 ( .A(a1stg_intlngop), .B(a1stg_in2[33]), .Z(N576) );
  GTECH_OR2 C2071 ( .A(N579), .B(N580), .Z(a1stg_norm_frac2[32]) );
  GTECH_OR2 C2072 ( .A(N577), .B(N578), .Z(N579) );
  GTECH_AND2 C2073 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[21]), .Z(N577) );
  GTECH_AND2 C2074 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[20]), .Z(N578) );
  GTECH_AND2 C2075 ( .A(a1stg_intlngop), .B(a1stg_in2[32]), .Z(N580) );
  GTECH_OR2 C2076 ( .A(N583), .B(N584), .Z(a1stg_norm_frac2[31]) );
  GTECH_OR2 C2077 ( .A(N581), .B(N582), .Z(N583) );
  GTECH_AND2 C2078 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[20]), .Z(N581) );
  GTECH_AND2 C2079 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[19]), .Z(N582) );
  GTECH_AND2 C2080 ( .A(a1stg_intlngop), .B(a1stg_in2[31]), .Z(N584) );
  GTECH_OR2 C2081 ( .A(N587), .B(N588), .Z(a1stg_norm_frac2[30]) );
  GTECH_OR2 C2082 ( .A(N585), .B(N586), .Z(N587) );
  GTECH_AND2 C2083 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[19]), .Z(N585) );
  GTECH_AND2 C2084 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[18]), .Z(N586) );
  GTECH_AND2 C2085 ( .A(a1stg_intlngop), .B(a1stg_in2[30]), .Z(N588) );
  GTECH_OR2 C2086 ( .A(N591), .B(N592), .Z(a1stg_norm_frac2[29]) );
  GTECH_OR2 C2087 ( .A(N589), .B(N590), .Z(N591) );
  GTECH_AND2 C2088 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[18]), .Z(N589) );
  GTECH_AND2 C2089 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[17]), .Z(N590) );
  GTECH_AND2 C2090 ( .A(a1stg_intlngop), .B(a1stg_in2[29]), .Z(N592) );
  GTECH_OR2 C2091 ( .A(N595), .B(N596), .Z(a1stg_norm_frac2[28]) );
  GTECH_OR2 C2092 ( .A(N593), .B(N594), .Z(N595) );
  GTECH_AND2 C2093 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[17]), .Z(N593) );
  GTECH_AND2 C2094 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[16]), .Z(N594) );
  GTECH_AND2 C2095 ( .A(a1stg_intlngop), .B(a1stg_in2[28]), .Z(N596) );
  GTECH_OR2 C2096 ( .A(N599), .B(N600), .Z(a1stg_norm_frac2[27]) );
  GTECH_OR2 C2097 ( .A(N597), .B(N598), .Z(N599) );
  GTECH_AND2 C2098 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[16]), .Z(N597) );
  GTECH_AND2 C2099 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[15]), .Z(N598) );
  GTECH_AND2 C2100 ( .A(a1stg_intlngop), .B(a1stg_in2[27]), .Z(N600) );
  GTECH_OR2 C2101 ( .A(N603), .B(N604), .Z(a1stg_norm_frac2[26]) );
  GTECH_OR2 C2102 ( .A(N601), .B(N602), .Z(N603) );
  GTECH_AND2 C2103 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[15]), .Z(N601) );
  GTECH_AND2 C2104 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[14]), .Z(N602) );
  GTECH_AND2 C2105 ( .A(a1stg_intlngop), .B(a1stg_in2[26]), .Z(N604) );
  GTECH_OR2 C2106 ( .A(N607), .B(N608), .Z(a1stg_norm_frac2[25]) );
  GTECH_OR2 C2107 ( .A(N605), .B(N606), .Z(N607) );
  GTECH_AND2 C2108 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[14]), .Z(N605) );
  GTECH_AND2 C2109 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[13]), .Z(N606) );
  GTECH_AND2 C2110 ( .A(a1stg_intlngop), .B(a1stg_in2[25]), .Z(N608) );
  GTECH_OR2 C2111 ( .A(N611), .B(N612), .Z(a1stg_norm_frac2[24]) );
  GTECH_OR2 C2112 ( .A(N609), .B(N610), .Z(N611) );
  GTECH_AND2 C2113 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[13]), .Z(N609) );
  GTECH_AND2 C2114 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[12]), .Z(N610) );
  GTECH_AND2 C2115 ( .A(a1stg_intlngop), .B(a1stg_in2[24]), .Z(N612) );
  GTECH_OR2 C2116 ( .A(N615), .B(N616), .Z(a1stg_norm_frac2[23]) );
  GTECH_OR2 C2117 ( .A(N613), .B(N614), .Z(N615) );
  GTECH_AND2 C2118 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[12]), .Z(N613) );
  GTECH_AND2 C2119 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[11]), .Z(N614) );
  GTECH_AND2 C2120 ( .A(a1stg_intlngop), .B(a1stg_in2[23]), .Z(N616) );
  GTECH_OR2 C2121 ( .A(N619), .B(N620), .Z(a1stg_norm_frac2[22]) );
  GTECH_OR2 C2122 ( .A(N617), .B(N618), .Z(N619) );
  GTECH_AND2 C2123 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[11]), .Z(N617) );
  GTECH_AND2 C2124 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[10]), .Z(N618) );
  GTECH_AND2 C2125 ( .A(a1stg_intlngop), .B(a1stg_in2[22]), .Z(N620) );
  GTECH_OR2 C2126 ( .A(N623), .B(N624), .Z(a1stg_norm_frac2[21]) );
  GTECH_OR2 C2127 ( .A(N621), .B(N622), .Z(N623) );
  GTECH_AND2 C2128 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[10]), .Z(N621) );
  GTECH_AND2 C2129 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[9]), .Z(N622) );
  GTECH_AND2 C2130 ( .A(a1stg_intlngop), .B(a1stg_in2[21]), .Z(N624) );
  GTECH_OR2 C2131 ( .A(N627), .B(N628), .Z(a1stg_norm_frac2[20]) );
  GTECH_OR2 C2132 ( .A(N625), .B(N626), .Z(N627) );
  GTECH_AND2 C2133 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[9]), .Z(N625) );
  GTECH_AND2 C2134 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[8]), .Z(N626) );
  GTECH_AND2 C2135 ( .A(a1stg_intlngop), .B(a1stg_in2[20]), .Z(N628) );
  GTECH_OR2 C2136 ( .A(N631), .B(N632), .Z(a1stg_norm_frac2[19]) );
  GTECH_OR2 C2137 ( .A(N629), .B(N630), .Z(N631) );
  GTECH_AND2 C2138 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[8]), .Z(N629) );
  GTECH_AND2 C2139 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[7]), .Z(N630) );
  GTECH_AND2 C2140 ( .A(a1stg_intlngop), .B(a1stg_in2[19]), .Z(N632) );
  GTECH_OR2 C2141 ( .A(N635), .B(N636), .Z(a1stg_norm_frac2[18]) );
  GTECH_OR2 C2142 ( .A(N633), .B(N634), .Z(N635) );
  GTECH_AND2 C2143 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[7]), .Z(N633) );
  GTECH_AND2 C2144 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[6]), .Z(N634) );
  GTECH_AND2 C2145 ( .A(a1stg_intlngop), .B(a1stg_in2[18]), .Z(N636) );
  GTECH_OR2 C2146 ( .A(N639), .B(N640), .Z(a1stg_norm_frac2[17]) );
  GTECH_OR2 C2147 ( .A(N637), .B(N638), .Z(N639) );
  GTECH_AND2 C2148 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[6]), .Z(N637) );
  GTECH_AND2 C2149 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[5]), .Z(N638) );
  GTECH_AND2 C2150 ( .A(a1stg_intlngop), .B(a1stg_in2[17]), .Z(N640) );
  GTECH_OR2 C2151 ( .A(N643), .B(N644), .Z(a1stg_norm_frac2[16]) );
  GTECH_OR2 C2152 ( .A(N641), .B(N642), .Z(N643) );
  GTECH_AND2 C2153 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[5]), .Z(N641) );
  GTECH_AND2 C2154 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[4]), .Z(N642) );
  GTECH_AND2 C2155 ( .A(a1stg_intlngop), .B(a1stg_in2[16]), .Z(N644) );
  GTECH_OR2 C2156 ( .A(N647), .B(N648), .Z(a1stg_norm_frac2[15]) );
  GTECH_OR2 C2157 ( .A(N645), .B(N646), .Z(N647) );
  GTECH_AND2 C2158 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[4]), .Z(N645) );
  GTECH_AND2 C2159 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[3]), .Z(N646) );
  GTECH_AND2 C2160 ( .A(a1stg_intlngop), .B(a1stg_in2[15]), .Z(N648) );
  GTECH_OR2 C2161 ( .A(N651), .B(N652), .Z(a1stg_norm_frac2[14]) );
  GTECH_OR2 C2162 ( .A(N649), .B(N650), .Z(N651) );
  GTECH_AND2 C2163 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[3]), .Z(N649) );
  GTECH_AND2 C2164 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[2]), .Z(N650) );
  GTECH_AND2 C2165 ( .A(a1stg_intlngop), .B(a1stg_in2[14]), .Z(N652) );
  GTECH_OR2 C2166 ( .A(N655), .B(N656), .Z(a1stg_norm_frac2[13]) );
  GTECH_OR2 C2167 ( .A(N653), .B(N654), .Z(N655) );
  GTECH_AND2 C2168 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[2]), .Z(N653) );
  GTECH_AND2 C2169 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[1]), .Z(N654) );
  GTECH_AND2 C2170 ( .A(a1stg_intlngop), .B(a1stg_in2[13]), .Z(N656) );
  GTECH_OR2 C2171 ( .A(N659), .B(N660), .Z(a1stg_norm_frac2[12]) );
  GTECH_OR2 C2172 ( .A(N657), .B(N658), .Z(N659) );
  GTECH_AND2 C2173 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[1]), .Z(N657) );
  GTECH_AND2 C2174 ( .A(a1stg_denorm_dbl_in2), .B(a1stg_in2[0]), .Z(N658) );
  GTECH_AND2 C2175 ( .A(a1stg_intlngop), .B(a1stg_in2[12]), .Z(N660) );
  GTECH_OR2 C2176 ( .A(N661), .B(N662), .Z(a1stg_norm_frac2[11]) );
  GTECH_AND2 C2177 ( .A(a1stg_norm_dbl_in2), .B(a1stg_in2[0]), .Z(N661) );
  GTECH_AND2 C2178 ( .A(a1stg_intlngop), .B(a1stg_in2[11]), .Z(N662) );
  GTECH_AND2 C2179 ( .A(a1stg_intlngop), .B(a1stg_in2[10]), .Z(
        a1stg_norm_frac2[10]) );
  GTECH_AND2 C2180 ( .A(a1stg_intlngop), .B(a1stg_in2[9]), .Z(
        a1stg_norm_frac2[9]) );
  GTECH_AND2 C2181 ( .A(a1stg_intlngop), .B(a1stg_in2[8]), .Z(
        a1stg_norm_frac2[8]) );
  GTECH_AND2 C2182 ( .A(a1stg_intlngop), .B(a1stg_in2[7]), .Z(
        a1stg_norm_frac2[7]) );
  GTECH_AND2 C2183 ( .A(a1stg_intlngop), .B(a1stg_in2[6]), .Z(
        a1stg_norm_frac2[6]) );
  GTECH_AND2 C2184 ( .A(a1stg_intlngop), .B(a1stg_in2[5]), .Z(
        a1stg_norm_frac2[5]) );
  GTECH_AND2 C2185 ( .A(a1stg_intlngop), .B(a1stg_in2[4]), .Z(
        a1stg_norm_frac2[4]) );
  GTECH_AND2 C2186 ( .A(a1stg_intlngop), .B(a1stg_in2[3]), .Z(
        a1stg_norm_frac2[3]) );
  GTECH_AND2 C2187 ( .A(a1stg_intlngop), .B(a1stg_in2[2]), .Z(
        a1stg_norm_frac2[2]) );
  GTECH_AND2 C2188 ( .A(a1stg_intlngop), .B(a1stg_in2[1]), .Z(
        a1stg_norm_frac2[1]) );
  GTECH_AND2 C2189 ( .A(a1stg_intlngop), .B(a1stg_in2[0]), .Z(
        a1stg_norm_frac2[0]) );
  GTECH_OR2 C2190 ( .A(N667), .B(N670), .Z(a2stg_frac1_in[63]) );
  GTECH_AND2 C2191 ( .A(N666), .B(a1stg_norm_frac1[63]), .Z(N667) );
  GTECH_OR2 C2192 ( .A(a1stg_faddsubop_inv), .B(N665), .Z(N666) );
  GTECH_NOT I_12 ( .A(N664), .Z(N665) );
  GTECH_OR2 C2194 ( .A(N663), .B(a2stg_frac1_in_frac1), .Z(N664) );
  GTECH_AND2 C2195 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N663) );
  GTECH_AND2 C2196 ( .A(N669), .B(a1stg_norm_frac2[63]), .Z(N670) );
  GTECH_AND2 C2197 ( .A(a2stg_frac1_in_frac2), .B(N668), .Z(N669) );
  GTECH_OR2 C2198 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N668)
         );
  GTECH_OR2 C2199 ( .A(N676), .B(N680), .Z(a2stg_frac1_in[62]) );
  GTECH_AND2 C2200 ( .A(N674), .B(N675), .Z(N676) );
  GTECH_OR2 C2201 ( .A(a1stg_faddsubop_inv), .B(N673), .Z(N674) );
  GTECH_NOT I_13 ( .A(N672), .Z(N673) );
  GTECH_OR2 C2203 ( .A(N671), .B(a2stg_frac1_in_frac1), .Z(N672) );
  GTECH_AND2 C2204 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N671) );
  GTECH_OR2 C2205 ( .A(a1stg_norm_frac1[62]), .B(a2stg_frac1_in_qnan), .Z(N675) );
  GTECH_AND2 C2206 ( .A(N678), .B(N679), .Z(N680) );
  GTECH_AND2 C2207 ( .A(a2stg_frac1_in_frac2), .B(N677), .Z(N678) );
  GTECH_OR2 C2208 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N677)
         );
  GTECH_OR2 C2209 ( .A(a1stg_norm_frac2[62]), .B(a2stg_frac1_in_qnan), .Z(N679) );
  GTECH_OR2 C2210 ( .A(N686), .B(N690), .Z(a2stg_frac1_in[61]) );
  GTECH_AND2 C2211 ( .A(N684), .B(N685), .Z(N686) );
  GTECH_OR2 C2212 ( .A(a1stg_faddsubop_inv), .B(N683), .Z(N684) );
  GTECH_NOT I_14 ( .A(N682), .Z(N683) );
  GTECH_OR2 C2214 ( .A(N681), .B(a2stg_frac1_in_frac1), .Z(N682) );
  GTECH_AND2 C2215 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N681) );
  GTECH_OR2 C2216 ( .A(a1stg_norm_frac1[61]), .B(a2stg_frac1_in_nv), .Z(N685)
         );
  GTECH_AND2 C2217 ( .A(N688), .B(N689), .Z(N690) );
  GTECH_AND2 C2218 ( .A(a2stg_frac1_in_frac2), .B(N687), .Z(N688) );
  GTECH_OR2 C2219 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N687)
         );
  GTECH_OR2 C2220 ( .A(a1stg_norm_frac2[61]), .B(a2stg_frac1_in_nv), .Z(N689)
         );
  GTECH_OR2 C2221 ( .A(N696), .B(N700), .Z(a2stg_frac1_in[60]) );
  GTECH_AND2 C2222 ( .A(N694), .B(N695), .Z(N696) );
  GTECH_OR2 C2223 ( .A(a1stg_faddsubop_inv), .B(N693), .Z(N694) );
  GTECH_NOT I_15 ( .A(N692), .Z(N693) );
  GTECH_OR2 C2225 ( .A(N691), .B(a2stg_frac1_in_frac1), .Z(N692) );
  GTECH_AND2 C2226 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N691) );
  GTECH_OR2 C2227 ( .A(a1stg_norm_frac1[60]), .B(a2stg_frac1_in_nv), .Z(N695)
         );
  GTECH_AND2 C2228 ( .A(N698), .B(N699), .Z(N700) );
  GTECH_AND2 C2229 ( .A(a2stg_frac1_in_frac2), .B(N697), .Z(N698) );
  GTECH_OR2 C2230 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N697)
         );
  GTECH_OR2 C2231 ( .A(a1stg_norm_frac2[60]), .B(a2stg_frac1_in_nv), .Z(N699)
         );
  GTECH_OR2 C2232 ( .A(N706), .B(N710), .Z(a2stg_frac1_in[59]) );
  GTECH_AND2 C2233 ( .A(N704), .B(N705), .Z(N706) );
  GTECH_OR2 C2234 ( .A(a1stg_faddsubop_inv), .B(N703), .Z(N704) );
  GTECH_NOT I_16 ( .A(N702), .Z(N703) );
  GTECH_OR2 C2236 ( .A(N701), .B(a2stg_frac1_in_frac1), .Z(N702) );
  GTECH_AND2 C2237 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N701) );
  GTECH_OR2 C2238 ( .A(a1stg_norm_frac1[59]), .B(a2stg_frac1_in_nv), .Z(N705)
         );
  GTECH_AND2 C2239 ( .A(N708), .B(N709), .Z(N710) );
  GTECH_AND2 C2240 ( .A(a2stg_frac1_in_frac2), .B(N707), .Z(N708) );
  GTECH_OR2 C2241 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N707)
         );
  GTECH_OR2 C2242 ( .A(a1stg_norm_frac2[59]), .B(a2stg_frac1_in_nv), .Z(N709)
         );
  GTECH_OR2 C2243 ( .A(N716), .B(N720), .Z(a2stg_frac1_in[58]) );
  GTECH_AND2 C2244 ( .A(N714), .B(N715), .Z(N716) );
  GTECH_OR2 C2245 ( .A(a1stg_faddsubop_inv), .B(N713), .Z(N714) );
  GTECH_NOT I_17 ( .A(N712), .Z(N713) );
  GTECH_OR2 C2247 ( .A(N711), .B(a2stg_frac1_in_frac1), .Z(N712) );
  GTECH_AND2 C2248 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N711) );
  GTECH_OR2 C2249 ( .A(a1stg_norm_frac1[58]), .B(a2stg_frac1_in_nv), .Z(N715)
         );
  GTECH_AND2 C2250 ( .A(N718), .B(N719), .Z(N720) );
  GTECH_AND2 C2251 ( .A(a2stg_frac1_in_frac2), .B(N717), .Z(N718) );
  GTECH_OR2 C2252 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N717)
         );
  GTECH_OR2 C2253 ( .A(a1stg_norm_frac2[58]), .B(a2stg_frac1_in_nv), .Z(N719)
         );
  GTECH_OR2 C2254 ( .A(N726), .B(N730), .Z(a2stg_frac1_in[57]) );
  GTECH_AND2 C2255 ( .A(N724), .B(N725), .Z(N726) );
  GTECH_OR2 C2256 ( .A(a1stg_faddsubop_inv), .B(N723), .Z(N724) );
  GTECH_NOT I_18 ( .A(N722), .Z(N723) );
  GTECH_OR2 C2258 ( .A(N721), .B(a2stg_frac1_in_frac1), .Z(N722) );
  GTECH_AND2 C2259 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N721) );
  GTECH_OR2 C2260 ( .A(a1stg_norm_frac1[57]), .B(a2stg_frac1_in_nv), .Z(N725)
         );
  GTECH_AND2 C2261 ( .A(N728), .B(N729), .Z(N730) );
  GTECH_AND2 C2262 ( .A(a2stg_frac1_in_frac2), .B(N727), .Z(N728) );
  GTECH_OR2 C2263 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N727)
         );
  GTECH_OR2 C2264 ( .A(a1stg_norm_frac2[57]), .B(a2stg_frac1_in_nv), .Z(N729)
         );
  GTECH_OR2 C2265 ( .A(N736), .B(N740), .Z(a2stg_frac1_in[56]) );
  GTECH_AND2 C2266 ( .A(N734), .B(N735), .Z(N736) );
  GTECH_OR2 C2267 ( .A(a1stg_faddsubop_inv), .B(N733), .Z(N734) );
  GTECH_NOT I_19 ( .A(N732), .Z(N733) );
  GTECH_OR2 C2269 ( .A(N731), .B(a2stg_frac1_in_frac1), .Z(N732) );
  GTECH_AND2 C2270 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N731) );
  GTECH_OR2 C2271 ( .A(a1stg_norm_frac1[56]), .B(a2stg_frac1_in_nv), .Z(N735)
         );
  GTECH_AND2 C2272 ( .A(N738), .B(N739), .Z(N740) );
  GTECH_AND2 C2273 ( .A(a2stg_frac1_in_frac2), .B(N737), .Z(N738) );
  GTECH_OR2 C2274 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N737)
         );
  GTECH_OR2 C2275 ( .A(a1stg_norm_frac2[56]), .B(a2stg_frac1_in_nv), .Z(N739)
         );
  GTECH_OR2 C2276 ( .A(N746), .B(N750), .Z(a2stg_frac1_in[55]) );
  GTECH_AND2 C2277 ( .A(N744), .B(N745), .Z(N746) );
  GTECH_OR2 C2278 ( .A(a1stg_faddsubop_inv), .B(N743), .Z(N744) );
  GTECH_NOT I_20 ( .A(N742), .Z(N743) );
  GTECH_OR2 C2280 ( .A(N741), .B(a2stg_frac1_in_frac1), .Z(N742) );
  GTECH_AND2 C2281 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N741) );
  GTECH_OR2 C2282 ( .A(a1stg_norm_frac1[55]), .B(a2stg_frac1_in_nv), .Z(N745)
         );
  GTECH_AND2 C2283 ( .A(N748), .B(N749), .Z(N750) );
  GTECH_AND2 C2284 ( .A(a2stg_frac1_in_frac2), .B(N747), .Z(N748) );
  GTECH_OR2 C2285 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N747)
         );
  GTECH_OR2 C2286 ( .A(a1stg_norm_frac2[55]), .B(a2stg_frac1_in_nv), .Z(N749)
         );
  GTECH_OR2 C2287 ( .A(N756), .B(N760), .Z(a2stg_frac1_in[54]) );
  GTECH_AND2 C2288 ( .A(N754), .B(N755), .Z(N756) );
  GTECH_OR2 C2289 ( .A(a1stg_faddsubop_inv), .B(N753), .Z(N754) );
  GTECH_NOT I_21 ( .A(N752), .Z(N753) );
  GTECH_OR2 C2291 ( .A(N751), .B(a2stg_frac1_in_frac1), .Z(N752) );
  GTECH_AND2 C2292 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N751) );
  GTECH_OR2 C2293 ( .A(a1stg_norm_frac1[54]), .B(a2stg_frac1_in_nv), .Z(N755)
         );
  GTECH_AND2 C2294 ( .A(N758), .B(N759), .Z(N760) );
  GTECH_AND2 C2295 ( .A(a2stg_frac1_in_frac2), .B(N757), .Z(N758) );
  GTECH_OR2 C2296 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N757)
         );
  GTECH_OR2 C2297 ( .A(a1stg_norm_frac2[54]), .B(a2stg_frac1_in_nv), .Z(N759)
         );
  GTECH_OR2 C2298 ( .A(N766), .B(N770), .Z(a2stg_frac1_in[53]) );
  GTECH_AND2 C2299 ( .A(N764), .B(N765), .Z(N766) );
  GTECH_OR2 C2300 ( .A(a1stg_faddsubop_inv), .B(N763), .Z(N764) );
  GTECH_NOT I_22 ( .A(N762), .Z(N763) );
  GTECH_OR2 C2302 ( .A(N761), .B(a2stg_frac1_in_frac1), .Z(N762) );
  GTECH_AND2 C2303 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N761) );
  GTECH_OR2 C2304 ( .A(a1stg_norm_frac1[53]), .B(a2stg_frac1_in_nv), .Z(N765)
         );
  GTECH_AND2 C2305 ( .A(N768), .B(N769), .Z(N770) );
  GTECH_AND2 C2306 ( .A(a2stg_frac1_in_frac2), .B(N767), .Z(N768) );
  GTECH_OR2 C2307 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N767)
         );
  GTECH_OR2 C2308 ( .A(a1stg_norm_frac2[53]), .B(a2stg_frac1_in_nv), .Z(N769)
         );
  GTECH_OR2 C2309 ( .A(N776), .B(N780), .Z(a2stg_frac1_in[52]) );
  GTECH_AND2 C2310 ( .A(N774), .B(N775), .Z(N776) );
  GTECH_OR2 C2311 ( .A(a1stg_faddsubop_inv), .B(N773), .Z(N774) );
  GTECH_NOT I_23 ( .A(N772), .Z(N773) );
  GTECH_OR2 C2313 ( .A(N771), .B(a2stg_frac1_in_frac1), .Z(N772) );
  GTECH_AND2 C2314 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N771) );
  GTECH_OR2 C2315 ( .A(a1stg_norm_frac1[52]), .B(a2stg_frac1_in_nv), .Z(N775)
         );
  GTECH_AND2 C2316 ( .A(N778), .B(N779), .Z(N780) );
  GTECH_AND2 C2317 ( .A(a2stg_frac1_in_frac2), .B(N777), .Z(N778) );
  GTECH_OR2 C2318 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N777)
         );
  GTECH_OR2 C2319 ( .A(a1stg_norm_frac2[52]), .B(a2stg_frac1_in_nv), .Z(N779)
         );
  GTECH_OR2 C2320 ( .A(N786), .B(N790), .Z(a2stg_frac1_in[51]) );
  GTECH_AND2 C2321 ( .A(N784), .B(N785), .Z(N786) );
  GTECH_OR2 C2322 ( .A(a1stg_faddsubop_inv), .B(N783), .Z(N784) );
  GTECH_NOT I_24 ( .A(N782), .Z(N783) );
  GTECH_OR2 C2324 ( .A(N781), .B(a2stg_frac1_in_frac1), .Z(N782) );
  GTECH_AND2 C2325 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N781) );
  GTECH_OR2 C2326 ( .A(a1stg_norm_frac1[51]), .B(a2stg_frac1_in_nv), .Z(N785)
         );
  GTECH_AND2 C2327 ( .A(N788), .B(N789), .Z(N790) );
  GTECH_AND2 C2328 ( .A(a2stg_frac1_in_frac2), .B(N787), .Z(N788) );
  GTECH_OR2 C2329 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N787)
         );
  GTECH_OR2 C2330 ( .A(a1stg_norm_frac2[51]), .B(a2stg_frac1_in_nv), .Z(N789)
         );
  GTECH_OR2 C2331 ( .A(N796), .B(N800), .Z(a2stg_frac1_in[50]) );
  GTECH_AND2 C2332 ( .A(N794), .B(N795), .Z(N796) );
  GTECH_OR2 C2333 ( .A(a1stg_faddsubop_inv), .B(N793), .Z(N794) );
  GTECH_NOT I_25 ( .A(N792), .Z(N793) );
  GTECH_OR2 C2335 ( .A(N791), .B(a2stg_frac1_in_frac1), .Z(N792) );
  GTECH_AND2 C2336 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N791) );
  GTECH_OR2 C2337 ( .A(a1stg_norm_frac1[50]), .B(a2stg_frac1_in_nv), .Z(N795)
         );
  GTECH_AND2 C2338 ( .A(N798), .B(N799), .Z(N800) );
  GTECH_AND2 C2339 ( .A(a2stg_frac1_in_frac2), .B(N797), .Z(N798) );
  GTECH_OR2 C2340 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N797)
         );
  GTECH_OR2 C2341 ( .A(a1stg_norm_frac2[50]), .B(a2stg_frac1_in_nv), .Z(N799)
         );
  GTECH_OR2 C2342 ( .A(N806), .B(N810), .Z(a2stg_frac1_in[49]) );
  GTECH_AND2 C2343 ( .A(N804), .B(N805), .Z(N806) );
  GTECH_OR2 C2344 ( .A(a1stg_faddsubop_inv), .B(N803), .Z(N804) );
  GTECH_NOT I_26 ( .A(N802), .Z(N803) );
  GTECH_OR2 C2346 ( .A(N801), .B(a2stg_frac1_in_frac1), .Z(N802) );
  GTECH_AND2 C2347 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N801) );
  GTECH_OR2 C2348 ( .A(a1stg_norm_frac1[49]), .B(a2stg_frac1_in_nv), .Z(N805)
         );
  GTECH_AND2 C2349 ( .A(N808), .B(N809), .Z(N810) );
  GTECH_AND2 C2350 ( .A(a2stg_frac1_in_frac2), .B(N807), .Z(N808) );
  GTECH_OR2 C2351 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N807)
         );
  GTECH_OR2 C2352 ( .A(a1stg_norm_frac2[49]), .B(a2stg_frac1_in_nv), .Z(N809)
         );
  GTECH_OR2 C2353 ( .A(N816), .B(N820), .Z(a2stg_frac1_in[48]) );
  GTECH_AND2 C2354 ( .A(N814), .B(N815), .Z(N816) );
  GTECH_OR2 C2355 ( .A(a1stg_faddsubop_inv), .B(N813), .Z(N814) );
  GTECH_NOT I_27 ( .A(N812), .Z(N813) );
  GTECH_OR2 C2357 ( .A(N811), .B(a2stg_frac1_in_frac1), .Z(N812) );
  GTECH_AND2 C2358 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N811) );
  GTECH_OR2 C2359 ( .A(a1stg_norm_frac1[48]), .B(a2stg_frac1_in_nv), .Z(N815)
         );
  GTECH_AND2 C2360 ( .A(N818), .B(N819), .Z(N820) );
  GTECH_AND2 C2361 ( .A(a2stg_frac1_in_frac2), .B(N817), .Z(N818) );
  GTECH_OR2 C2362 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N817)
         );
  GTECH_OR2 C2363 ( .A(a1stg_norm_frac2[48]), .B(a2stg_frac1_in_nv), .Z(N819)
         );
  GTECH_OR2 C2364 ( .A(N826), .B(N830), .Z(a2stg_frac1_in[47]) );
  GTECH_AND2 C2365 ( .A(N824), .B(N825), .Z(N826) );
  GTECH_OR2 C2366 ( .A(a1stg_faddsubop_inv), .B(N823), .Z(N824) );
  GTECH_NOT I_28 ( .A(N822), .Z(N823) );
  GTECH_OR2 C2368 ( .A(N821), .B(a2stg_frac1_in_frac1), .Z(N822) );
  GTECH_AND2 C2369 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N821) );
  GTECH_OR2 C2370 ( .A(a1stg_norm_frac1[47]), .B(a2stg_frac1_in_nv), .Z(N825)
         );
  GTECH_AND2 C2371 ( .A(N828), .B(N829), .Z(N830) );
  GTECH_AND2 C2372 ( .A(a2stg_frac1_in_frac2), .B(N827), .Z(N828) );
  GTECH_OR2 C2373 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N827)
         );
  GTECH_OR2 C2374 ( .A(a1stg_norm_frac2[47]), .B(a2stg_frac1_in_nv), .Z(N829)
         );
  GTECH_OR2 C2375 ( .A(N836), .B(N840), .Z(a2stg_frac1_in[46]) );
  GTECH_AND2 C2376 ( .A(N834), .B(N835), .Z(N836) );
  GTECH_OR2 C2377 ( .A(a1stg_faddsubop_inv), .B(N833), .Z(N834) );
  GTECH_NOT I_29 ( .A(N832), .Z(N833) );
  GTECH_OR2 C2379 ( .A(N831), .B(a2stg_frac1_in_frac1), .Z(N832) );
  GTECH_AND2 C2380 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N831) );
  GTECH_OR2 C2381 ( .A(a1stg_norm_frac1[46]), .B(a2stg_frac1_in_nv), .Z(N835)
         );
  GTECH_AND2 C2382 ( .A(N838), .B(N839), .Z(N840) );
  GTECH_AND2 C2383 ( .A(a2stg_frac1_in_frac2), .B(N837), .Z(N838) );
  GTECH_OR2 C2384 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N837)
         );
  GTECH_OR2 C2385 ( .A(a1stg_norm_frac2[46]), .B(a2stg_frac1_in_nv), .Z(N839)
         );
  GTECH_OR2 C2386 ( .A(N846), .B(N850), .Z(a2stg_frac1_in[45]) );
  GTECH_AND2 C2387 ( .A(N844), .B(N845), .Z(N846) );
  GTECH_OR2 C2388 ( .A(a1stg_faddsubop_inv), .B(N843), .Z(N844) );
  GTECH_NOT I_30 ( .A(N842), .Z(N843) );
  GTECH_OR2 C2390 ( .A(N841), .B(a2stg_frac1_in_frac1), .Z(N842) );
  GTECH_AND2 C2391 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N841) );
  GTECH_OR2 C2392 ( .A(a1stg_norm_frac1[45]), .B(a2stg_frac1_in_nv), .Z(N845)
         );
  GTECH_AND2 C2393 ( .A(N848), .B(N849), .Z(N850) );
  GTECH_AND2 C2394 ( .A(a2stg_frac1_in_frac2), .B(N847), .Z(N848) );
  GTECH_OR2 C2395 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N847)
         );
  GTECH_OR2 C2396 ( .A(a1stg_norm_frac2[45]), .B(a2stg_frac1_in_nv), .Z(N849)
         );
  GTECH_OR2 C2397 ( .A(N856), .B(N860), .Z(a2stg_frac1_in[44]) );
  GTECH_AND2 C2398 ( .A(N854), .B(N855), .Z(N856) );
  GTECH_OR2 C2399 ( .A(a1stg_faddsubop_inv), .B(N853), .Z(N854) );
  GTECH_NOT I_31 ( .A(N852), .Z(N853) );
  GTECH_OR2 C2401 ( .A(N851), .B(a2stg_frac1_in_frac1), .Z(N852) );
  GTECH_AND2 C2402 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N851) );
  GTECH_OR2 C2403 ( .A(a1stg_norm_frac1[44]), .B(a2stg_frac1_in_nv), .Z(N855)
         );
  GTECH_AND2 C2404 ( .A(N858), .B(N859), .Z(N860) );
  GTECH_AND2 C2405 ( .A(a2stg_frac1_in_frac2), .B(N857), .Z(N858) );
  GTECH_OR2 C2406 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N857)
         );
  GTECH_OR2 C2407 ( .A(a1stg_norm_frac2[44]), .B(a2stg_frac1_in_nv), .Z(N859)
         );
  GTECH_OR2 C2408 ( .A(N866), .B(N870), .Z(a2stg_frac1_in[43]) );
  GTECH_AND2 C2409 ( .A(N864), .B(N865), .Z(N866) );
  GTECH_OR2 C2410 ( .A(a1stg_faddsubop_inv), .B(N863), .Z(N864) );
  GTECH_NOT I_32 ( .A(N862), .Z(N863) );
  GTECH_OR2 C2412 ( .A(N861), .B(a2stg_frac1_in_frac1), .Z(N862) );
  GTECH_AND2 C2413 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N861) );
  GTECH_OR2 C2414 ( .A(a1stg_norm_frac1[43]), .B(a2stg_frac1_in_nv), .Z(N865)
         );
  GTECH_AND2 C2415 ( .A(N868), .B(N869), .Z(N870) );
  GTECH_AND2 C2416 ( .A(a2stg_frac1_in_frac2), .B(N867), .Z(N868) );
  GTECH_OR2 C2417 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N867)
         );
  GTECH_OR2 C2418 ( .A(a1stg_norm_frac2[43]), .B(a2stg_frac1_in_nv), .Z(N869)
         );
  GTECH_OR2 C2419 ( .A(N876), .B(N880), .Z(a2stg_frac1_in[42]) );
  GTECH_AND2 C2420 ( .A(N874), .B(N875), .Z(N876) );
  GTECH_OR2 C2421 ( .A(a1stg_faddsubop_inv), .B(N873), .Z(N874) );
  GTECH_NOT I_33 ( .A(N872), .Z(N873) );
  GTECH_OR2 C2423 ( .A(N871), .B(a2stg_frac1_in_frac1), .Z(N872) );
  GTECH_AND2 C2424 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N871) );
  GTECH_OR2 C2425 ( .A(a1stg_norm_frac1[42]), .B(a2stg_frac1_in_nv), .Z(N875)
         );
  GTECH_AND2 C2426 ( .A(N878), .B(N879), .Z(N880) );
  GTECH_AND2 C2427 ( .A(a2stg_frac1_in_frac2), .B(N877), .Z(N878) );
  GTECH_OR2 C2428 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N877)
         );
  GTECH_OR2 C2429 ( .A(a1stg_norm_frac2[42]), .B(a2stg_frac1_in_nv), .Z(N879)
         );
  GTECH_OR2 C2430 ( .A(N886), .B(N890), .Z(a2stg_frac1_in[41]) );
  GTECH_AND2 C2431 ( .A(N884), .B(N885), .Z(N886) );
  GTECH_OR2 C2432 ( .A(a1stg_faddsubop_inv), .B(N883), .Z(N884) );
  GTECH_NOT I_34 ( .A(N882), .Z(N883) );
  GTECH_OR2 C2434 ( .A(N881), .B(a2stg_frac1_in_frac1), .Z(N882) );
  GTECH_AND2 C2435 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N881) );
  GTECH_OR2 C2436 ( .A(a1stg_norm_frac1[41]), .B(a2stg_frac1_in_nv), .Z(N885)
         );
  GTECH_AND2 C2437 ( .A(N888), .B(N889), .Z(N890) );
  GTECH_AND2 C2438 ( .A(a2stg_frac1_in_frac2), .B(N887), .Z(N888) );
  GTECH_OR2 C2439 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N887)
         );
  GTECH_OR2 C2440 ( .A(a1stg_norm_frac2[41]), .B(a2stg_frac1_in_nv), .Z(N889)
         );
  GTECH_OR2 C2441 ( .A(N896), .B(N900), .Z(a2stg_frac1_in[40]) );
  GTECH_AND2 C2442 ( .A(N894), .B(N895), .Z(N896) );
  GTECH_OR2 C2443 ( .A(a1stg_faddsubop_inv), .B(N893), .Z(N894) );
  GTECH_NOT I_35 ( .A(N892), .Z(N893) );
  GTECH_OR2 C2445 ( .A(N891), .B(a2stg_frac1_in_frac1), .Z(N892) );
  GTECH_AND2 C2446 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N891) );
  GTECH_OR2 C2447 ( .A(a1stg_norm_frac1[40]), .B(a2stg_frac1_in_nv), .Z(N895)
         );
  GTECH_AND2 C2448 ( .A(N898), .B(N899), .Z(N900) );
  GTECH_AND2 C2449 ( .A(a2stg_frac1_in_frac2), .B(N897), .Z(N898) );
  GTECH_OR2 C2450 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N897)
         );
  GTECH_OR2 C2451 ( .A(a1stg_norm_frac2[40]), .B(a2stg_frac1_in_nv), .Z(N899)
         );
  GTECH_OR2 C2452 ( .A(N906), .B(N910), .Z(a2stg_frac1_in[39]) );
  GTECH_AND2 C2453 ( .A(N904), .B(N905), .Z(N906) );
  GTECH_OR2 C2454 ( .A(a1stg_faddsubop_inv), .B(N903), .Z(N904) );
  GTECH_NOT I_36 ( .A(N902), .Z(N903) );
  GTECH_OR2 C2456 ( .A(N901), .B(a2stg_frac1_in_frac1), .Z(N902) );
  GTECH_AND2 C2457 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N901) );
  GTECH_OR2 C2458 ( .A(a1stg_norm_frac1[39]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N905) );
  GTECH_AND2 C2459 ( .A(N908), .B(N909), .Z(N910) );
  GTECH_AND2 C2460 ( .A(a2stg_frac1_in_frac2), .B(N907), .Z(N908) );
  GTECH_OR2 C2461 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N907)
         );
  GTECH_OR2 C2462 ( .A(a1stg_norm_frac2[39]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N909) );
  GTECH_OR2 C2463 ( .A(N916), .B(N920), .Z(a2stg_frac1_in[38]) );
  GTECH_AND2 C2464 ( .A(N914), .B(N915), .Z(N916) );
  GTECH_OR2 C2465 ( .A(a1stg_faddsubop_inv), .B(N913), .Z(N914) );
  GTECH_NOT I_37 ( .A(N912), .Z(N913) );
  GTECH_OR2 C2467 ( .A(N911), .B(a2stg_frac1_in_frac1), .Z(N912) );
  GTECH_AND2 C2468 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N911) );
  GTECH_OR2 C2469 ( .A(a1stg_norm_frac1[38]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N915) );
  GTECH_AND2 C2470 ( .A(N918), .B(N919), .Z(N920) );
  GTECH_AND2 C2471 ( .A(a2stg_frac1_in_frac2), .B(N917), .Z(N918) );
  GTECH_OR2 C2472 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N917)
         );
  GTECH_OR2 C2473 ( .A(a1stg_norm_frac2[38]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N919) );
  GTECH_OR2 C2474 ( .A(N926), .B(N930), .Z(a2stg_frac1_in[37]) );
  GTECH_AND2 C2475 ( .A(N924), .B(N925), .Z(N926) );
  GTECH_OR2 C2476 ( .A(a1stg_faddsubop_inv), .B(N923), .Z(N924) );
  GTECH_NOT I_38 ( .A(N922), .Z(N923) );
  GTECH_OR2 C2478 ( .A(N921), .B(a2stg_frac1_in_frac1), .Z(N922) );
  GTECH_AND2 C2479 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N921) );
  GTECH_OR2 C2480 ( .A(a1stg_norm_frac1[37]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N925) );
  GTECH_AND2 C2481 ( .A(N928), .B(N929), .Z(N930) );
  GTECH_AND2 C2482 ( .A(a2stg_frac1_in_frac2), .B(N927), .Z(N928) );
  GTECH_OR2 C2483 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N927)
         );
  GTECH_OR2 C2484 ( .A(a1stg_norm_frac2[37]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N929) );
  GTECH_OR2 C2485 ( .A(N936), .B(N940), .Z(a2stg_frac1_in[36]) );
  GTECH_AND2 C2486 ( .A(N934), .B(N935), .Z(N936) );
  GTECH_OR2 C2487 ( .A(a1stg_faddsubop_inv), .B(N933), .Z(N934) );
  GTECH_NOT I_39 ( .A(N932), .Z(N933) );
  GTECH_OR2 C2489 ( .A(N931), .B(a2stg_frac1_in_frac1), .Z(N932) );
  GTECH_AND2 C2490 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N931) );
  GTECH_OR2 C2491 ( .A(a1stg_norm_frac1[36]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N935) );
  GTECH_AND2 C2492 ( .A(N938), .B(N939), .Z(N940) );
  GTECH_AND2 C2493 ( .A(a2stg_frac1_in_frac2), .B(N937), .Z(N938) );
  GTECH_OR2 C2494 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N937)
         );
  GTECH_OR2 C2495 ( .A(a1stg_norm_frac2[36]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N939) );
  GTECH_OR2 C2496 ( .A(N946), .B(N950), .Z(a2stg_frac1_in[35]) );
  GTECH_AND2 C2497 ( .A(N944), .B(N945), .Z(N946) );
  GTECH_OR2 C2498 ( .A(a1stg_faddsubop_inv), .B(N943), .Z(N944) );
  GTECH_NOT I_40 ( .A(N942), .Z(N943) );
  GTECH_OR2 C2500 ( .A(N941), .B(a2stg_frac1_in_frac1), .Z(N942) );
  GTECH_AND2 C2501 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N941) );
  GTECH_OR2 C2502 ( .A(a1stg_norm_frac1[35]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N945) );
  GTECH_AND2 C2503 ( .A(N948), .B(N949), .Z(N950) );
  GTECH_AND2 C2504 ( .A(a2stg_frac1_in_frac2), .B(N947), .Z(N948) );
  GTECH_OR2 C2505 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N947)
         );
  GTECH_OR2 C2506 ( .A(a1stg_norm_frac2[35]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N949) );
  GTECH_OR2 C2507 ( .A(N956), .B(N960), .Z(a2stg_frac1_in[34]) );
  GTECH_AND2 C2508 ( .A(N954), .B(N955), .Z(N956) );
  GTECH_OR2 C2509 ( .A(a1stg_faddsubop_inv), .B(N953), .Z(N954) );
  GTECH_NOT I_41 ( .A(N952), .Z(N953) );
  GTECH_OR2 C2511 ( .A(N951), .B(a2stg_frac1_in_frac1), .Z(N952) );
  GTECH_AND2 C2512 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N951) );
  GTECH_OR2 C2513 ( .A(a1stg_norm_frac1[34]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N955) );
  GTECH_AND2 C2514 ( .A(N958), .B(N959), .Z(N960) );
  GTECH_AND2 C2515 ( .A(a2stg_frac1_in_frac2), .B(N957), .Z(N958) );
  GTECH_OR2 C2516 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N957)
         );
  GTECH_OR2 C2517 ( .A(a1stg_norm_frac2[34]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N959) );
  GTECH_OR2 C2518 ( .A(N966), .B(N970), .Z(a2stg_frac1_in[33]) );
  GTECH_AND2 C2519 ( .A(N964), .B(N965), .Z(N966) );
  GTECH_OR2 C2520 ( .A(a1stg_faddsubop_inv), .B(N963), .Z(N964) );
  GTECH_NOT I_42 ( .A(N962), .Z(N963) );
  GTECH_OR2 C2522 ( .A(N961), .B(a2stg_frac1_in_frac1), .Z(N962) );
  GTECH_AND2 C2523 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N961) );
  GTECH_OR2 C2524 ( .A(a1stg_norm_frac1[33]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N965) );
  GTECH_AND2 C2525 ( .A(N968), .B(N969), .Z(N970) );
  GTECH_AND2 C2526 ( .A(a2stg_frac1_in_frac2), .B(N967), .Z(N968) );
  GTECH_OR2 C2527 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N967)
         );
  GTECH_OR2 C2528 ( .A(a1stg_norm_frac2[33]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N969) );
  GTECH_OR2 C2529 ( .A(N976), .B(N980), .Z(a2stg_frac1_in[32]) );
  GTECH_AND2 C2530 ( .A(N974), .B(N975), .Z(N976) );
  GTECH_OR2 C2531 ( .A(a1stg_faddsubop_inv), .B(N973), .Z(N974) );
  GTECH_NOT I_43 ( .A(N972), .Z(N973) );
  GTECH_OR2 C2533 ( .A(N971), .B(a2stg_frac1_in_frac1), .Z(N972) );
  GTECH_AND2 C2534 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N971) );
  GTECH_OR2 C2535 ( .A(a1stg_norm_frac1[32]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N975) );
  GTECH_AND2 C2536 ( .A(N978), .B(N979), .Z(N980) );
  GTECH_AND2 C2537 ( .A(a2stg_frac1_in_frac2), .B(N977), .Z(N978) );
  GTECH_OR2 C2538 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N977)
         );
  GTECH_OR2 C2539 ( .A(a1stg_norm_frac2[32]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N979) );
  GTECH_OR2 C2540 ( .A(N986), .B(N990), .Z(a2stg_frac1_in[31]) );
  GTECH_AND2 C2541 ( .A(N984), .B(N985), .Z(N986) );
  GTECH_OR2 C2542 ( .A(a1stg_faddsubop_inv), .B(N983), .Z(N984) );
  GTECH_NOT I_44 ( .A(N982), .Z(N983) );
  GTECH_OR2 C2544 ( .A(N981), .B(a2stg_frac1_in_frac1), .Z(N982) );
  GTECH_AND2 C2545 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N981) );
  GTECH_OR2 C2546 ( .A(a1stg_norm_frac1[31]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N985) );
  GTECH_AND2 C2547 ( .A(N988), .B(N989), .Z(N990) );
  GTECH_AND2 C2548 ( .A(a2stg_frac1_in_frac2), .B(N987), .Z(N988) );
  GTECH_OR2 C2549 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N987)
         );
  GTECH_OR2 C2550 ( .A(a1stg_norm_frac2[31]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N989) );
  GTECH_OR2 C2551 ( .A(N996), .B(N1000), .Z(a2stg_frac1_in[30]) );
  GTECH_AND2 C2552 ( .A(N994), .B(N995), .Z(N996) );
  GTECH_OR2 C2553 ( .A(a1stg_faddsubop_inv), .B(N993), .Z(N994) );
  GTECH_NOT I_45 ( .A(N992), .Z(N993) );
  GTECH_OR2 C2555 ( .A(N991), .B(a2stg_frac1_in_frac1), .Z(N992) );
  GTECH_AND2 C2556 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N991) );
  GTECH_OR2 C2557 ( .A(a1stg_norm_frac1[30]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N995) );
  GTECH_AND2 C2558 ( .A(N998), .B(N999), .Z(N1000) );
  GTECH_AND2 C2559 ( .A(a2stg_frac1_in_frac2), .B(N997), .Z(N998) );
  GTECH_OR2 C2560 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N997)
         );
  GTECH_OR2 C2561 ( .A(a1stg_norm_frac2[30]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N999) );
  GTECH_OR2 C2562 ( .A(N1006), .B(N1010), .Z(a2stg_frac1_in[29]) );
  GTECH_AND2 C2563 ( .A(N1004), .B(N1005), .Z(N1006) );
  GTECH_OR2 C2564 ( .A(a1stg_faddsubop_inv), .B(N1003), .Z(N1004) );
  GTECH_NOT I_46 ( .A(N1002), .Z(N1003) );
  GTECH_OR2 C2566 ( .A(N1001), .B(a2stg_frac1_in_frac1), .Z(N1002) );
  GTECH_AND2 C2567 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1001) );
  GTECH_OR2 C2568 ( .A(a1stg_norm_frac1[29]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1005) );
  GTECH_AND2 C2569 ( .A(N1008), .B(N1009), .Z(N1010) );
  GTECH_AND2 C2570 ( .A(a2stg_frac1_in_frac2), .B(N1007), .Z(N1008) );
  GTECH_OR2 C2571 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1007)
         );
  GTECH_OR2 C2572 ( .A(a1stg_norm_frac2[29]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1009) );
  GTECH_OR2 C2573 ( .A(N1016), .B(N1020), .Z(a2stg_frac1_in[28]) );
  GTECH_AND2 C2574 ( .A(N1014), .B(N1015), .Z(N1016) );
  GTECH_OR2 C2575 ( .A(a1stg_faddsubop_inv), .B(N1013), .Z(N1014) );
  GTECH_NOT I_47 ( .A(N1012), .Z(N1013) );
  GTECH_OR2 C2577 ( .A(N1011), .B(a2stg_frac1_in_frac1), .Z(N1012) );
  GTECH_AND2 C2578 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1011) );
  GTECH_OR2 C2579 ( .A(a1stg_norm_frac1[28]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1015) );
  GTECH_AND2 C2580 ( .A(N1018), .B(N1019), .Z(N1020) );
  GTECH_AND2 C2581 ( .A(a2stg_frac1_in_frac2), .B(N1017), .Z(N1018) );
  GTECH_OR2 C2582 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1017)
         );
  GTECH_OR2 C2583 ( .A(a1stg_norm_frac2[28]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1019) );
  GTECH_OR2 C2584 ( .A(N1026), .B(N1030), .Z(a2stg_frac1_in[27]) );
  GTECH_AND2 C2585 ( .A(N1024), .B(N1025), .Z(N1026) );
  GTECH_OR2 C2586 ( .A(a1stg_faddsubop_inv), .B(N1023), .Z(N1024) );
  GTECH_NOT I_48 ( .A(N1022), .Z(N1023) );
  GTECH_OR2 C2588 ( .A(N1021), .B(a2stg_frac1_in_frac1), .Z(N1022) );
  GTECH_AND2 C2589 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1021) );
  GTECH_OR2 C2590 ( .A(a1stg_norm_frac1[27]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1025) );
  GTECH_AND2 C2591 ( .A(N1028), .B(N1029), .Z(N1030) );
  GTECH_AND2 C2592 ( .A(a2stg_frac1_in_frac2), .B(N1027), .Z(N1028) );
  GTECH_OR2 C2593 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1027)
         );
  GTECH_OR2 C2594 ( .A(a1stg_norm_frac2[27]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1029) );
  GTECH_OR2 C2595 ( .A(N1036), .B(N1040), .Z(a2stg_frac1_in[26]) );
  GTECH_AND2 C2596 ( .A(N1034), .B(N1035), .Z(N1036) );
  GTECH_OR2 C2597 ( .A(a1stg_faddsubop_inv), .B(N1033), .Z(N1034) );
  GTECH_NOT I_49 ( .A(N1032), .Z(N1033) );
  GTECH_OR2 C2599 ( .A(N1031), .B(a2stg_frac1_in_frac1), .Z(N1032) );
  GTECH_AND2 C2600 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1031) );
  GTECH_OR2 C2601 ( .A(a1stg_norm_frac1[26]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1035) );
  GTECH_AND2 C2602 ( .A(N1038), .B(N1039), .Z(N1040) );
  GTECH_AND2 C2603 ( .A(a2stg_frac1_in_frac2), .B(N1037), .Z(N1038) );
  GTECH_OR2 C2604 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1037)
         );
  GTECH_OR2 C2605 ( .A(a1stg_norm_frac2[26]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1039) );
  GTECH_OR2 C2606 ( .A(N1046), .B(N1050), .Z(a2stg_frac1_in[25]) );
  GTECH_AND2 C2607 ( .A(N1044), .B(N1045), .Z(N1046) );
  GTECH_OR2 C2608 ( .A(a1stg_faddsubop_inv), .B(N1043), .Z(N1044) );
  GTECH_NOT I_50 ( .A(N1042), .Z(N1043) );
  GTECH_OR2 C2610 ( .A(N1041), .B(a2stg_frac1_in_frac1), .Z(N1042) );
  GTECH_AND2 C2611 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1041) );
  GTECH_OR2 C2612 ( .A(a1stg_norm_frac1[25]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1045) );
  GTECH_AND2 C2613 ( .A(N1048), .B(N1049), .Z(N1050) );
  GTECH_AND2 C2614 ( .A(a2stg_frac1_in_frac2), .B(N1047), .Z(N1048) );
  GTECH_OR2 C2615 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1047)
         );
  GTECH_OR2 C2616 ( .A(a1stg_norm_frac2[25]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1049) );
  GTECH_OR2 C2617 ( .A(N1056), .B(N1060), .Z(a2stg_frac1_in[24]) );
  GTECH_AND2 C2618 ( .A(N1054), .B(N1055), .Z(N1056) );
  GTECH_OR2 C2619 ( .A(a1stg_faddsubop_inv), .B(N1053), .Z(N1054) );
  GTECH_NOT I_51 ( .A(N1052), .Z(N1053) );
  GTECH_OR2 C2621 ( .A(N1051), .B(a2stg_frac1_in_frac1), .Z(N1052) );
  GTECH_AND2 C2622 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1051) );
  GTECH_OR2 C2623 ( .A(a1stg_norm_frac1[24]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1055) );
  GTECH_AND2 C2624 ( .A(N1058), .B(N1059), .Z(N1060) );
  GTECH_AND2 C2625 ( .A(a2stg_frac1_in_frac2), .B(N1057), .Z(N1058) );
  GTECH_OR2 C2626 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1057)
         );
  GTECH_OR2 C2627 ( .A(a1stg_norm_frac2[24]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1059) );
  GTECH_OR2 C2628 ( .A(N1066), .B(N1070), .Z(a2stg_frac1_in[23]) );
  GTECH_AND2 C2629 ( .A(N1064), .B(N1065), .Z(N1066) );
  GTECH_OR2 C2630 ( .A(a1stg_faddsubop_inv), .B(N1063), .Z(N1064) );
  GTECH_NOT I_52 ( .A(N1062), .Z(N1063) );
  GTECH_OR2 C2632 ( .A(N1061), .B(a2stg_frac1_in_frac1), .Z(N1062) );
  GTECH_AND2 C2633 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1061) );
  GTECH_OR2 C2634 ( .A(a1stg_norm_frac1[23]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1065) );
  GTECH_AND2 C2635 ( .A(N1068), .B(N1069), .Z(N1070) );
  GTECH_AND2 C2636 ( .A(a2stg_frac1_in_frac2), .B(N1067), .Z(N1068) );
  GTECH_OR2 C2637 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1067)
         );
  GTECH_OR2 C2638 ( .A(a1stg_norm_frac2[23]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1069) );
  GTECH_OR2 C2639 ( .A(N1076), .B(N1080), .Z(a2stg_frac1_in[22]) );
  GTECH_AND2 C2640 ( .A(N1074), .B(N1075), .Z(N1076) );
  GTECH_OR2 C2641 ( .A(a1stg_faddsubop_inv), .B(N1073), .Z(N1074) );
  GTECH_NOT I_53 ( .A(N1072), .Z(N1073) );
  GTECH_OR2 C2643 ( .A(N1071), .B(a2stg_frac1_in_frac1), .Z(N1072) );
  GTECH_AND2 C2644 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1071) );
  GTECH_OR2 C2645 ( .A(a1stg_norm_frac1[22]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1075) );
  GTECH_AND2 C2646 ( .A(N1078), .B(N1079), .Z(N1080) );
  GTECH_AND2 C2647 ( .A(a2stg_frac1_in_frac2), .B(N1077), .Z(N1078) );
  GTECH_OR2 C2648 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1077)
         );
  GTECH_OR2 C2649 ( .A(a1stg_norm_frac2[22]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1079) );
  GTECH_OR2 C2650 ( .A(N1086), .B(N1090), .Z(a2stg_frac1_in[21]) );
  GTECH_AND2 C2651 ( .A(N1084), .B(N1085), .Z(N1086) );
  GTECH_OR2 C2652 ( .A(a1stg_faddsubop_inv), .B(N1083), .Z(N1084) );
  GTECH_NOT I_54 ( .A(N1082), .Z(N1083) );
  GTECH_OR2 C2654 ( .A(N1081), .B(a2stg_frac1_in_frac1), .Z(N1082) );
  GTECH_AND2 C2655 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1081) );
  GTECH_OR2 C2656 ( .A(a1stg_norm_frac1[21]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1085) );
  GTECH_AND2 C2657 ( .A(N1088), .B(N1089), .Z(N1090) );
  GTECH_AND2 C2658 ( .A(a2stg_frac1_in_frac2), .B(N1087), .Z(N1088) );
  GTECH_OR2 C2659 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1087)
         );
  GTECH_OR2 C2660 ( .A(a1stg_norm_frac2[21]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1089) );
  GTECH_OR2 C2661 ( .A(N1096), .B(N1100), .Z(a2stg_frac1_in[20]) );
  GTECH_AND2 C2662 ( .A(N1094), .B(N1095), .Z(N1096) );
  GTECH_OR2 C2663 ( .A(a1stg_faddsubop_inv), .B(N1093), .Z(N1094) );
  GTECH_NOT I_55 ( .A(N1092), .Z(N1093) );
  GTECH_OR2 C2665 ( .A(N1091), .B(a2stg_frac1_in_frac1), .Z(N1092) );
  GTECH_AND2 C2666 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1091) );
  GTECH_OR2 C2667 ( .A(a1stg_norm_frac1[20]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1095) );
  GTECH_AND2 C2668 ( .A(N1098), .B(N1099), .Z(N1100) );
  GTECH_AND2 C2669 ( .A(a2stg_frac1_in_frac2), .B(N1097), .Z(N1098) );
  GTECH_OR2 C2670 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1097)
         );
  GTECH_OR2 C2671 ( .A(a1stg_norm_frac2[20]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1099) );
  GTECH_OR2 C2672 ( .A(N1106), .B(N1110), .Z(a2stg_frac1_in[19]) );
  GTECH_AND2 C2673 ( .A(N1104), .B(N1105), .Z(N1106) );
  GTECH_OR2 C2674 ( .A(a1stg_faddsubop_inv), .B(N1103), .Z(N1104) );
  GTECH_NOT I_56 ( .A(N1102), .Z(N1103) );
  GTECH_OR2 C2676 ( .A(N1101), .B(a2stg_frac1_in_frac1), .Z(N1102) );
  GTECH_AND2 C2677 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1101) );
  GTECH_OR2 C2678 ( .A(a1stg_norm_frac1[19]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1105) );
  GTECH_AND2 C2679 ( .A(N1108), .B(N1109), .Z(N1110) );
  GTECH_AND2 C2680 ( .A(a2stg_frac1_in_frac2), .B(N1107), .Z(N1108) );
  GTECH_OR2 C2681 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1107)
         );
  GTECH_OR2 C2682 ( .A(a1stg_norm_frac2[19]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1109) );
  GTECH_OR2 C2683 ( .A(N1116), .B(N1120), .Z(a2stg_frac1_in[18]) );
  GTECH_AND2 C2684 ( .A(N1114), .B(N1115), .Z(N1116) );
  GTECH_OR2 C2685 ( .A(a1stg_faddsubop_inv), .B(N1113), .Z(N1114) );
  GTECH_NOT I_57 ( .A(N1112), .Z(N1113) );
  GTECH_OR2 C2687 ( .A(N1111), .B(a2stg_frac1_in_frac1), .Z(N1112) );
  GTECH_AND2 C2688 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1111) );
  GTECH_OR2 C2689 ( .A(a1stg_norm_frac1[18]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1115) );
  GTECH_AND2 C2690 ( .A(N1118), .B(N1119), .Z(N1120) );
  GTECH_AND2 C2691 ( .A(a2stg_frac1_in_frac2), .B(N1117), .Z(N1118) );
  GTECH_OR2 C2692 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1117)
         );
  GTECH_OR2 C2693 ( .A(a1stg_norm_frac2[18]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1119) );
  GTECH_OR2 C2694 ( .A(N1126), .B(N1130), .Z(a2stg_frac1_in[17]) );
  GTECH_AND2 C2695 ( .A(N1124), .B(N1125), .Z(N1126) );
  GTECH_OR2 C2696 ( .A(a1stg_faddsubop_inv), .B(N1123), .Z(N1124) );
  GTECH_NOT I_58 ( .A(N1122), .Z(N1123) );
  GTECH_OR2 C2698 ( .A(N1121), .B(a2stg_frac1_in_frac1), .Z(N1122) );
  GTECH_AND2 C2699 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1121) );
  GTECH_OR2 C2700 ( .A(a1stg_norm_frac1[17]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1125) );
  GTECH_AND2 C2701 ( .A(N1128), .B(N1129), .Z(N1130) );
  GTECH_AND2 C2702 ( .A(a2stg_frac1_in_frac2), .B(N1127), .Z(N1128) );
  GTECH_OR2 C2703 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1127)
         );
  GTECH_OR2 C2704 ( .A(a1stg_norm_frac2[17]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1129) );
  GTECH_OR2 C2705 ( .A(N1136), .B(N1140), .Z(a2stg_frac1_in[16]) );
  GTECH_AND2 C2706 ( .A(N1134), .B(N1135), .Z(N1136) );
  GTECH_OR2 C2707 ( .A(a1stg_faddsubop_inv), .B(N1133), .Z(N1134) );
  GTECH_NOT I_59 ( .A(N1132), .Z(N1133) );
  GTECH_OR2 C2709 ( .A(N1131), .B(a2stg_frac1_in_frac1), .Z(N1132) );
  GTECH_AND2 C2710 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1131) );
  GTECH_OR2 C2711 ( .A(a1stg_norm_frac1[16]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1135) );
  GTECH_AND2 C2712 ( .A(N1138), .B(N1139), .Z(N1140) );
  GTECH_AND2 C2713 ( .A(a2stg_frac1_in_frac2), .B(N1137), .Z(N1138) );
  GTECH_OR2 C2714 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1137)
         );
  GTECH_OR2 C2715 ( .A(a1stg_norm_frac2[16]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1139) );
  GTECH_OR2 C2716 ( .A(N1146), .B(N1150), .Z(a2stg_frac1_in[15]) );
  GTECH_AND2 C2717 ( .A(N1144), .B(N1145), .Z(N1146) );
  GTECH_OR2 C2718 ( .A(a1stg_faddsubop_inv), .B(N1143), .Z(N1144) );
  GTECH_NOT I_60 ( .A(N1142), .Z(N1143) );
  GTECH_OR2 C2720 ( .A(N1141), .B(a2stg_frac1_in_frac1), .Z(N1142) );
  GTECH_AND2 C2721 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1141) );
  GTECH_OR2 C2722 ( .A(a1stg_norm_frac1[15]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1145) );
  GTECH_AND2 C2723 ( .A(N1148), .B(N1149), .Z(N1150) );
  GTECH_AND2 C2724 ( .A(a2stg_frac1_in_frac2), .B(N1147), .Z(N1148) );
  GTECH_OR2 C2725 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1147)
         );
  GTECH_OR2 C2726 ( .A(a1stg_norm_frac2[15]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1149) );
  GTECH_OR2 C2727 ( .A(N1156), .B(N1160), .Z(a2stg_frac1_in[14]) );
  GTECH_AND2 C2728 ( .A(N1154), .B(N1155), .Z(N1156) );
  GTECH_OR2 C2729 ( .A(a1stg_faddsubop_inv), .B(N1153), .Z(N1154) );
  GTECH_NOT I_61 ( .A(N1152), .Z(N1153) );
  GTECH_OR2 C2731 ( .A(N1151), .B(a2stg_frac1_in_frac1), .Z(N1152) );
  GTECH_AND2 C2732 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1151) );
  GTECH_OR2 C2733 ( .A(a1stg_norm_frac1[14]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1155) );
  GTECH_AND2 C2734 ( .A(N1158), .B(N1159), .Z(N1160) );
  GTECH_AND2 C2735 ( .A(a2stg_frac1_in_frac2), .B(N1157), .Z(N1158) );
  GTECH_OR2 C2736 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1157)
         );
  GTECH_OR2 C2737 ( .A(a1stg_norm_frac2[14]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1159) );
  GTECH_OR2 C2738 ( .A(N1166), .B(N1170), .Z(a2stg_frac1_in[13]) );
  GTECH_AND2 C2739 ( .A(N1164), .B(N1165), .Z(N1166) );
  GTECH_OR2 C2740 ( .A(a1stg_faddsubop_inv), .B(N1163), .Z(N1164) );
  GTECH_NOT I_62 ( .A(N1162), .Z(N1163) );
  GTECH_OR2 C2742 ( .A(N1161), .B(a2stg_frac1_in_frac1), .Z(N1162) );
  GTECH_AND2 C2743 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1161) );
  GTECH_OR2 C2744 ( .A(a1stg_norm_frac1[13]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1165) );
  GTECH_AND2 C2745 ( .A(N1168), .B(N1169), .Z(N1170) );
  GTECH_AND2 C2746 ( .A(a2stg_frac1_in_frac2), .B(N1167), .Z(N1168) );
  GTECH_OR2 C2747 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1167)
         );
  GTECH_OR2 C2748 ( .A(a1stg_norm_frac2[13]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1169) );
  GTECH_OR2 C2749 ( .A(N1176), .B(N1180), .Z(a2stg_frac1_in[12]) );
  GTECH_AND2 C2750 ( .A(N1174), .B(N1175), .Z(N1176) );
  GTECH_OR2 C2751 ( .A(a1stg_faddsubop_inv), .B(N1173), .Z(N1174) );
  GTECH_NOT I_63 ( .A(N1172), .Z(N1173) );
  GTECH_OR2 C2753 ( .A(N1171), .B(a2stg_frac1_in_frac1), .Z(N1172) );
  GTECH_AND2 C2754 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1171) );
  GTECH_OR2 C2755 ( .A(a1stg_norm_frac1[12]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1175) );
  GTECH_AND2 C2756 ( .A(N1178), .B(N1179), .Z(N1180) );
  GTECH_AND2 C2757 ( .A(a2stg_frac1_in_frac2), .B(N1177), .Z(N1178) );
  GTECH_OR2 C2758 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1177)
         );
  GTECH_OR2 C2759 ( .A(a1stg_norm_frac2[12]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1179) );
  GTECH_OR2 C2760 ( .A(N1186), .B(N1190), .Z(a2stg_frac1_in[11]) );
  GTECH_AND2 C2761 ( .A(N1184), .B(N1185), .Z(N1186) );
  GTECH_OR2 C2762 ( .A(a1stg_faddsubop_inv), .B(N1183), .Z(N1184) );
  GTECH_NOT I_64 ( .A(N1182), .Z(N1183) );
  GTECH_OR2 C2764 ( .A(N1181), .B(a2stg_frac1_in_frac1), .Z(N1182) );
  GTECH_AND2 C2765 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1181) );
  GTECH_OR2 C2766 ( .A(a1stg_norm_frac1[11]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1185) );
  GTECH_AND2 C2767 ( .A(N1188), .B(N1189), .Z(N1190) );
  GTECH_AND2 C2768 ( .A(a2stg_frac1_in_frac2), .B(N1187), .Z(N1188) );
  GTECH_OR2 C2769 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1187)
         );
  GTECH_OR2 C2770 ( .A(a1stg_norm_frac2[11]), .B(a2stg_frac1_in_nv_dbl), .Z(
        N1189) );
  GTECH_OR2 C2771 ( .A(N1195), .B(N1198), .Z(a2stg_frac1_in[10]) );
  GTECH_AND2 C2772 ( .A(N1194), .B(1'b0), .Z(N1195) );
  GTECH_OR2 C2773 ( .A(a1stg_faddsubop_inv), .B(N1193), .Z(N1194) );
  GTECH_NOT I_65 ( .A(N1192), .Z(N1193) );
  GTECH_OR2 C2775 ( .A(N1191), .B(a2stg_frac1_in_frac1), .Z(N1192) );
  GTECH_AND2 C2776 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1191) );
  GTECH_AND2 C2777 ( .A(N1197), .B(a1stg_norm_frac2[10]), .Z(N1198) );
  GTECH_AND2 C2778 ( .A(a2stg_frac1_in_frac2), .B(N1196), .Z(N1197) );
  GTECH_OR2 C2779 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1196)
         );
  GTECH_OR2 C2780 ( .A(N1203), .B(N1206), .Z(a2stg_frac1_in[9]) );
  GTECH_AND2 C2781 ( .A(N1202), .B(1'b0), .Z(N1203) );
  GTECH_OR2 C2782 ( .A(a1stg_faddsubop_inv), .B(N1201), .Z(N1202) );
  GTECH_NOT I_66 ( .A(N1200), .Z(N1201) );
  GTECH_OR2 C2784 ( .A(N1199), .B(a2stg_frac1_in_frac1), .Z(N1200) );
  GTECH_AND2 C2785 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1199) );
  GTECH_AND2 C2786 ( .A(N1205), .B(a1stg_norm_frac2[9]), .Z(N1206) );
  GTECH_AND2 C2787 ( .A(a2stg_frac1_in_frac2), .B(N1204), .Z(N1205) );
  GTECH_OR2 C2788 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1204)
         );
  GTECH_OR2 C2789 ( .A(N1211), .B(N1214), .Z(a2stg_frac1_in[8]) );
  GTECH_AND2 C2790 ( .A(N1210), .B(1'b0), .Z(N1211) );
  GTECH_OR2 C2791 ( .A(a1stg_faddsubop_inv), .B(N1209), .Z(N1210) );
  GTECH_NOT I_67 ( .A(N1208), .Z(N1209) );
  GTECH_OR2 C2793 ( .A(N1207), .B(a2stg_frac1_in_frac1), .Z(N1208) );
  GTECH_AND2 C2794 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1207) );
  GTECH_AND2 C2795 ( .A(N1213), .B(a1stg_norm_frac2[8]), .Z(N1214) );
  GTECH_AND2 C2796 ( .A(a2stg_frac1_in_frac2), .B(N1212), .Z(N1213) );
  GTECH_OR2 C2797 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1212)
         );
  GTECH_OR2 C2798 ( .A(N1219), .B(N1222), .Z(a2stg_frac1_in[7]) );
  GTECH_AND2 C2799 ( .A(N1218), .B(1'b0), .Z(N1219) );
  GTECH_OR2 C2800 ( .A(a1stg_faddsubop_inv), .B(N1217), .Z(N1218) );
  GTECH_NOT I_68 ( .A(N1216), .Z(N1217) );
  GTECH_OR2 C2802 ( .A(N1215), .B(a2stg_frac1_in_frac1), .Z(N1216) );
  GTECH_AND2 C2803 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1215) );
  GTECH_AND2 C2804 ( .A(N1221), .B(a1stg_norm_frac2[7]), .Z(N1222) );
  GTECH_AND2 C2805 ( .A(a2stg_frac1_in_frac2), .B(N1220), .Z(N1221) );
  GTECH_OR2 C2806 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1220)
         );
  GTECH_OR2 C2807 ( .A(N1227), .B(N1230), .Z(a2stg_frac1_in[6]) );
  GTECH_AND2 C2808 ( .A(N1226), .B(1'b0), .Z(N1227) );
  GTECH_OR2 C2809 ( .A(a1stg_faddsubop_inv), .B(N1225), .Z(N1226) );
  GTECH_NOT I_69 ( .A(N1224), .Z(N1225) );
  GTECH_OR2 C2811 ( .A(N1223), .B(a2stg_frac1_in_frac1), .Z(N1224) );
  GTECH_AND2 C2812 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1223) );
  GTECH_AND2 C2813 ( .A(N1229), .B(a1stg_norm_frac2[6]), .Z(N1230) );
  GTECH_AND2 C2814 ( .A(a2stg_frac1_in_frac2), .B(N1228), .Z(N1229) );
  GTECH_OR2 C2815 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1228)
         );
  GTECH_OR2 C2816 ( .A(N1235), .B(N1238), .Z(a2stg_frac1_in[5]) );
  GTECH_AND2 C2817 ( .A(N1234), .B(1'b0), .Z(N1235) );
  GTECH_OR2 C2818 ( .A(a1stg_faddsubop_inv), .B(N1233), .Z(N1234) );
  GTECH_NOT I_70 ( .A(N1232), .Z(N1233) );
  GTECH_OR2 C2820 ( .A(N1231), .B(a2stg_frac1_in_frac1), .Z(N1232) );
  GTECH_AND2 C2821 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1231) );
  GTECH_AND2 C2822 ( .A(N1237), .B(a1stg_norm_frac2[5]), .Z(N1238) );
  GTECH_AND2 C2823 ( .A(a2stg_frac1_in_frac2), .B(N1236), .Z(N1237) );
  GTECH_OR2 C2824 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1236)
         );
  GTECH_OR2 C2825 ( .A(N1243), .B(N1246), .Z(a2stg_frac1_in[4]) );
  GTECH_AND2 C2826 ( .A(N1242), .B(1'b0), .Z(N1243) );
  GTECH_OR2 C2827 ( .A(a1stg_faddsubop_inv), .B(N1241), .Z(N1242) );
  GTECH_NOT I_71 ( .A(N1240), .Z(N1241) );
  GTECH_OR2 C2829 ( .A(N1239), .B(a2stg_frac1_in_frac1), .Z(N1240) );
  GTECH_AND2 C2830 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1239) );
  GTECH_AND2 C2831 ( .A(N1245), .B(a1stg_norm_frac2[4]), .Z(N1246) );
  GTECH_AND2 C2832 ( .A(a2stg_frac1_in_frac2), .B(N1244), .Z(N1245) );
  GTECH_OR2 C2833 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1244)
         );
  GTECH_OR2 C2834 ( .A(N1251), .B(N1254), .Z(a2stg_frac1_in[3]) );
  GTECH_AND2 C2835 ( .A(N1250), .B(1'b0), .Z(N1251) );
  GTECH_OR2 C2836 ( .A(a1stg_faddsubop_inv), .B(N1249), .Z(N1250) );
  GTECH_NOT I_72 ( .A(N1248), .Z(N1249) );
  GTECH_OR2 C2838 ( .A(N1247), .B(a2stg_frac1_in_frac1), .Z(N1248) );
  GTECH_AND2 C2839 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1247) );
  GTECH_AND2 C2840 ( .A(N1253), .B(a1stg_norm_frac2[3]), .Z(N1254) );
  GTECH_AND2 C2841 ( .A(a2stg_frac1_in_frac2), .B(N1252), .Z(N1253) );
  GTECH_OR2 C2842 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1252)
         );
  GTECH_OR2 C2843 ( .A(N1259), .B(N1262), .Z(a2stg_frac1_in[2]) );
  GTECH_AND2 C2844 ( .A(N1258), .B(1'b0), .Z(N1259) );
  GTECH_OR2 C2845 ( .A(a1stg_faddsubop_inv), .B(N1257), .Z(N1258) );
  GTECH_NOT I_73 ( .A(N1256), .Z(N1257) );
  GTECH_OR2 C2847 ( .A(N1255), .B(a2stg_frac1_in_frac1), .Z(N1256) );
  GTECH_AND2 C2848 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1255) );
  GTECH_AND2 C2849 ( .A(N1261), .B(a1stg_norm_frac2[2]), .Z(N1262) );
  GTECH_AND2 C2850 ( .A(a2stg_frac1_in_frac2), .B(N1260), .Z(N1261) );
  GTECH_OR2 C2851 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1260)
         );
  GTECH_OR2 C2852 ( .A(N1267), .B(N1270), .Z(a2stg_frac1_in[1]) );
  GTECH_AND2 C2853 ( .A(N1266), .B(1'b0), .Z(N1267) );
  GTECH_OR2 C2854 ( .A(a1stg_faddsubop_inv), .B(N1265), .Z(N1266) );
  GTECH_NOT I_74 ( .A(N1264), .Z(N1265) );
  GTECH_OR2 C2856 ( .A(N1263), .B(a2stg_frac1_in_frac1), .Z(N1264) );
  GTECH_AND2 C2857 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1263) );
  GTECH_AND2 C2858 ( .A(N1269), .B(a1stg_norm_frac2[1]), .Z(N1270) );
  GTECH_AND2 C2859 ( .A(a2stg_frac1_in_frac2), .B(N1268), .Z(N1269) );
  GTECH_OR2 C2860 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1268)
         );
  GTECH_OR2 C2861 ( .A(N1275), .B(N1278), .Z(a2stg_frac1_in[0]) );
  GTECH_AND2 C2862 ( .A(N1274), .B(1'b0), .Z(N1275) );
  GTECH_OR2 C2863 ( .A(a1stg_faddsubop_inv), .B(N1273), .Z(N1274) );
  GTECH_NOT I_75 ( .A(N1272), .Z(N1273) );
  GTECH_OR2 C2865 ( .A(N1271), .B(a2stg_frac1_in_frac1), .Z(N1272) );
  GTECH_AND2 C2866 ( .A(a1stg_in2_gt_in1), .B(a1stg_2nan_in_inv), .Z(N1271) );
  GTECH_AND2 C2867 ( .A(N1277), .B(a1stg_norm_frac2[0]), .Z(N1278) );
  GTECH_AND2 C2868 ( .A(a2stg_frac1_in_frac2), .B(N1276), .Z(N1277) );
  GTECH_OR2 C2869 ( .A(a1stg_in2_gt_in1), .B(a2stg_frac1_in_frac1), .Z(N1276)
         );
  GTECH_OR2 C2870 ( .A(a1stg_norm_frac2[62]), .B(a2stg_frac2_in_qnan), .Z(N0)
         );
  GTECH_OR2 C2871 ( .A(N1283), .B(N1285), .Z(a2stg_frac2_in[63]) );
  GTECH_OR2 C2872 ( .A(N1279), .B(N1282), .Z(N1283) );
  GTECH_AND2 C2873 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[63]), .Z(
        N1279) );
  GTECH_AND2 C2874 ( .A(N1281), .B(a1stg_norm_frac2[63]), .Z(N1282) );
  GTECH_AND2 C2875 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1281) );
  GTECH_NOT I_76 ( .A(a1stg_in2_gt_in1), .Z(N1280) );
  GTECH_AND2 C2877 ( .A(N1284), .B(a1stg_norm_frac1[63]), .Z(N1285) );
  GTECH_AND2 C2878 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1284)
         );
  GTECH_OR2 C2879 ( .A(N1289), .B(N1291), .Z(a2stg_frac2_in[62]) );
  GTECH_OR2 C2880 ( .A(N1286), .B(N1288), .Z(N1289) );
  GTECH_AND2 C2881 ( .A(a1stg_faddsubop_inv), .B(N0), .Z(N1286) );
  GTECH_AND2 C2882 ( .A(N1287), .B(N0), .Z(N1288) );
  GTECH_AND2 C2883 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1287) );
  GTECH_AND2 C2885 ( .A(N1290), .B(a1stg_norm_frac1[62]), .Z(N1291) );
  GTECH_AND2 C2886 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1290)
         );
  GTECH_OR2 C2887 ( .A(N1295), .B(N1297), .Z(a2stg_frac2_in[61]) );
  GTECH_OR2 C2888 ( .A(N1292), .B(N1294), .Z(N1295) );
  GTECH_AND2 C2889 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[61]), .Z(
        N1292) );
  GTECH_AND2 C2890 ( .A(N1293), .B(a1stg_norm_frac2[61]), .Z(N1294) );
  GTECH_AND2 C2891 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1293) );
  GTECH_AND2 C2893 ( .A(N1296), .B(a1stg_norm_frac1[61]), .Z(N1297) );
  GTECH_AND2 C2894 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1296)
         );
  GTECH_OR2 C2895 ( .A(N1301), .B(N1303), .Z(a2stg_frac2_in[60]) );
  GTECH_OR2 C2896 ( .A(N1298), .B(N1300), .Z(N1301) );
  GTECH_AND2 C2897 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[60]), .Z(
        N1298) );
  GTECH_AND2 C2898 ( .A(N1299), .B(a1stg_norm_frac2[60]), .Z(N1300) );
  GTECH_AND2 C2899 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1299) );
  GTECH_AND2 C2901 ( .A(N1302), .B(a1stg_norm_frac1[60]), .Z(N1303) );
  GTECH_AND2 C2902 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1302)
         );
  GTECH_OR2 C2903 ( .A(N1307), .B(N1309), .Z(a2stg_frac2_in[59]) );
  GTECH_OR2 C2904 ( .A(N1304), .B(N1306), .Z(N1307) );
  GTECH_AND2 C2905 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[59]), .Z(
        N1304) );
  GTECH_AND2 C2906 ( .A(N1305), .B(a1stg_norm_frac2[59]), .Z(N1306) );
  GTECH_AND2 C2907 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1305) );
  GTECH_AND2 C2909 ( .A(N1308), .B(a1stg_norm_frac1[59]), .Z(N1309) );
  GTECH_AND2 C2910 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1308)
         );
  GTECH_OR2 C2911 ( .A(N1313), .B(N1315), .Z(a2stg_frac2_in[58]) );
  GTECH_OR2 C2912 ( .A(N1310), .B(N1312), .Z(N1313) );
  GTECH_AND2 C2913 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[58]), .Z(
        N1310) );
  GTECH_AND2 C2914 ( .A(N1311), .B(a1stg_norm_frac2[58]), .Z(N1312) );
  GTECH_AND2 C2915 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1311) );
  GTECH_AND2 C2917 ( .A(N1314), .B(a1stg_norm_frac1[58]), .Z(N1315) );
  GTECH_AND2 C2918 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1314)
         );
  GTECH_OR2 C2919 ( .A(N1319), .B(N1321), .Z(a2stg_frac2_in[57]) );
  GTECH_OR2 C2920 ( .A(N1316), .B(N1318), .Z(N1319) );
  GTECH_AND2 C2921 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[57]), .Z(
        N1316) );
  GTECH_AND2 C2922 ( .A(N1317), .B(a1stg_norm_frac2[57]), .Z(N1318) );
  GTECH_AND2 C2923 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1317) );
  GTECH_AND2 C2925 ( .A(N1320), .B(a1stg_norm_frac1[57]), .Z(N1321) );
  GTECH_AND2 C2926 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1320)
         );
  GTECH_OR2 C2927 ( .A(N1325), .B(N1327), .Z(a2stg_frac2_in[56]) );
  GTECH_OR2 C2928 ( .A(N1322), .B(N1324), .Z(N1325) );
  GTECH_AND2 C2929 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[56]), .Z(
        N1322) );
  GTECH_AND2 C2930 ( .A(N1323), .B(a1stg_norm_frac2[56]), .Z(N1324) );
  GTECH_AND2 C2931 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1323) );
  GTECH_AND2 C2933 ( .A(N1326), .B(a1stg_norm_frac1[56]), .Z(N1327) );
  GTECH_AND2 C2934 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1326)
         );
  GTECH_OR2 C2935 ( .A(N1331), .B(N1333), .Z(a2stg_frac2_in[55]) );
  GTECH_OR2 C2936 ( .A(N1328), .B(N1330), .Z(N1331) );
  GTECH_AND2 C2937 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[55]), .Z(
        N1328) );
  GTECH_AND2 C2938 ( .A(N1329), .B(a1stg_norm_frac2[55]), .Z(N1330) );
  GTECH_AND2 C2939 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1329) );
  GTECH_AND2 C2941 ( .A(N1332), .B(a1stg_norm_frac1[55]), .Z(N1333) );
  GTECH_AND2 C2942 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1332)
         );
  GTECH_OR2 C2943 ( .A(N1337), .B(N1339), .Z(a2stg_frac2_in[54]) );
  GTECH_OR2 C2944 ( .A(N1334), .B(N1336), .Z(N1337) );
  GTECH_AND2 C2945 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[54]), .Z(
        N1334) );
  GTECH_AND2 C2946 ( .A(N1335), .B(a1stg_norm_frac2[54]), .Z(N1336) );
  GTECH_AND2 C2947 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1335) );
  GTECH_AND2 C2949 ( .A(N1338), .B(a1stg_norm_frac1[54]), .Z(N1339) );
  GTECH_AND2 C2950 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1338)
         );
  GTECH_OR2 C2951 ( .A(N1343), .B(N1345), .Z(a2stg_frac2_in[53]) );
  GTECH_OR2 C2952 ( .A(N1340), .B(N1342), .Z(N1343) );
  GTECH_AND2 C2953 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[53]), .Z(
        N1340) );
  GTECH_AND2 C2954 ( .A(N1341), .B(a1stg_norm_frac2[53]), .Z(N1342) );
  GTECH_AND2 C2955 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1341) );
  GTECH_AND2 C2957 ( .A(N1344), .B(a1stg_norm_frac1[53]), .Z(N1345) );
  GTECH_AND2 C2958 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1344)
         );
  GTECH_OR2 C2959 ( .A(N1349), .B(N1351), .Z(a2stg_frac2_in[52]) );
  GTECH_OR2 C2960 ( .A(N1346), .B(N1348), .Z(N1349) );
  GTECH_AND2 C2961 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[52]), .Z(
        N1346) );
  GTECH_AND2 C2962 ( .A(N1347), .B(a1stg_norm_frac2[52]), .Z(N1348) );
  GTECH_AND2 C2963 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1347) );
  GTECH_AND2 C2965 ( .A(N1350), .B(a1stg_norm_frac1[52]), .Z(N1351) );
  GTECH_AND2 C2966 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1350)
         );
  GTECH_OR2 C2967 ( .A(N1355), .B(N1357), .Z(a2stg_frac2_in[51]) );
  GTECH_OR2 C2968 ( .A(N1352), .B(N1354), .Z(N1355) );
  GTECH_AND2 C2969 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[51]), .Z(
        N1352) );
  GTECH_AND2 C2970 ( .A(N1353), .B(a1stg_norm_frac2[51]), .Z(N1354) );
  GTECH_AND2 C2971 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1353) );
  GTECH_AND2 C2973 ( .A(N1356), .B(a1stg_norm_frac1[51]), .Z(N1357) );
  GTECH_AND2 C2974 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1356)
         );
  GTECH_OR2 C2975 ( .A(N1361), .B(N1363), .Z(a2stg_frac2_in[50]) );
  GTECH_OR2 C2976 ( .A(N1358), .B(N1360), .Z(N1361) );
  GTECH_AND2 C2977 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[50]), .Z(
        N1358) );
  GTECH_AND2 C2978 ( .A(N1359), .B(a1stg_norm_frac2[50]), .Z(N1360) );
  GTECH_AND2 C2979 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1359) );
  GTECH_AND2 C2981 ( .A(N1362), .B(a1stg_norm_frac1[50]), .Z(N1363) );
  GTECH_AND2 C2982 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1362)
         );
  GTECH_OR2 C2983 ( .A(N1367), .B(N1369), .Z(a2stg_frac2_in[49]) );
  GTECH_OR2 C2984 ( .A(N1364), .B(N1366), .Z(N1367) );
  GTECH_AND2 C2985 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[49]), .Z(
        N1364) );
  GTECH_AND2 C2986 ( .A(N1365), .B(a1stg_norm_frac2[49]), .Z(N1366) );
  GTECH_AND2 C2987 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1365) );
  GTECH_AND2 C2989 ( .A(N1368), .B(a1stg_norm_frac1[49]), .Z(N1369) );
  GTECH_AND2 C2990 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1368)
         );
  GTECH_OR2 C2991 ( .A(N1373), .B(N1375), .Z(a2stg_frac2_in[48]) );
  GTECH_OR2 C2992 ( .A(N1370), .B(N1372), .Z(N1373) );
  GTECH_AND2 C2993 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[48]), .Z(
        N1370) );
  GTECH_AND2 C2994 ( .A(N1371), .B(a1stg_norm_frac2[48]), .Z(N1372) );
  GTECH_AND2 C2995 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1371) );
  GTECH_AND2 C2997 ( .A(N1374), .B(a1stg_norm_frac1[48]), .Z(N1375) );
  GTECH_AND2 C2998 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1374)
         );
  GTECH_OR2 C2999 ( .A(N1379), .B(N1381), .Z(a2stg_frac2_in[47]) );
  GTECH_OR2 C3000 ( .A(N1376), .B(N1378), .Z(N1379) );
  GTECH_AND2 C3001 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[47]), .Z(
        N1376) );
  GTECH_AND2 C3002 ( .A(N1377), .B(a1stg_norm_frac2[47]), .Z(N1378) );
  GTECH_AND2 C3003 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1377) );
  GTECH_AND2 C3005 ( .A(N1380), .B(a1stg_norm_frac1[47]), .Z(N1381) );
  GTECH_AND2 C3006 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1380)
         );
  GTECH_OR2 C3007 ( .A(N1385), .B(N1387), .Z(a2stg_frac2_in[46]) );
  GTECH_OR2 C3008 ( .A(N1382), .B(N1384), .Z(N1385) );
  GTECH_AND2 C3009 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[46]), .Z(
        N1382) );
  GTECH_AND2 C3010 ( .A(N1383), .B(a1stg_norm_frac2[46]), .Z(N1384) );
  GTECH_AND2 C3011 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1383) );
  GTECH_AND2 C3013 ( .A(N1386), .B(a1stg_norm_frac1[46]), .Z(N1387) );
  GTECH_AND2 C3014 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1386)
         );
  GTECH_OR2 C3015 ( .A(N1391), .B(N1393), .Z(a2stg_frac2_in[45]) );
  GTECH_OR2 C3016 ( .A(N1388), .B(N1390), .Z(N1391) );
  GTECH_AND2 C3017 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[45]), .Z(
        N1388) );
  GTECH_AND2 C3018 ( .A(N1389), .B(a1stg_norm_frac2[45]), .Z(N1390) );
  GTECH_AND2 C3019 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1389) );
  GTECH_AND2 C3021 ( .A(N1392), .B(a1stg_norm_frac1[45]), .Z(N1393) );
  GTECH_AND2 C3022 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1392)
         );
  GTECH_OR2 C3023 ( .A(N1397), .B(N1399), .Z(a2stg_frac2_in[44]) );
  GTECH_OR2 C3024 ( .A(N1394), .B(N1396), .Z(N1397) );
  GTECH_AND2 C3025 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[44]), .Z(
        N1394) );
  GTECH_AND2 C3026 ( .A(N1395), .B(a1stg_norm_frac2[44]), .Z(N1396) );
  GTECH_AND2 C3027 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1395) );
  GTECH_AND2 C3029 ( .A(N1398), .B(a1stg_norm_frac1[44]), .Z(N1399) );
  GTECH_AND2 C3030 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1398)
         );
  GTECH_OR2 C3031 ( .A(N1403), .B(N1405), .Z(a2stg_frac2_in[43]) );
  GTECH_OR2 C3032 ( .A(N1400), .B(N1402), .Z(N1403) );
  GTECH_AND2 C3033 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[43]), .Z(
        N1400) );
  GTECH_AND2 C3034 ( .A(N1401), .B(a1stg_norm_frac2[43]), .Z(N1402) );
  GTECH_AND2 C3035 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1401) );
  GTECH_AND2 C3037 ( .A(N1404), .B(a1stg_norm_frac1[43]), .Z(N1405) );
  GTECH_AND2 C3038 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1404)
         );
  GTECH_OR2 C3039 ( .A(N1409), .B(N1411), .Z(a2stg_frac2_in[42]) );
  GTECH_OR2 C3040 ( .A(N1406), .B(N1408), .Z(N1409) );
  GTECH_AND2 C3041 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[42]), .Z(
        N1406) );
  GTECH_AND2 C3042 ( .A(N1407), .B(a1stg_norm_frac2[42]), .Z(N1408) );
  GTECH_AND2 C3043 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1407) );
  GTECH_AND2 C3045 ( .A(N1410), .B(a1stg_norm_frac1[42]), .Z(N1411) );
  GTECH_AND2 C3046 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1410)
         );
  GTECH_OR2 C3047 ( .A(N1415), .B(N1417), .Z(a2stg_frac2_in[41]) );
  GTECH_OR2 C3048 ( .A(N1412), .B(N1414), .Z(N1415) );
  GTECH_AND2 C3049 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[41]), .Z(
        N1412) );
  GTECH_AND2 C3050 ( .A(N1413), .B(a1stg_norm_frac2[41]), .Z(N1414) );
  GTECH_AND2 C3051 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1413) );
  GTECH_AND2 C3053 ( .A(N1416), .B(a1stg_norm_frac1[41]), .Z(N1417) );
  GTECH_AND2 C3054 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1416)
         );
  GTECH_OR2 C3055 ( .A(N1421), .B(N1423), .Z(a2stg_frac2_in[40]) );
  GTECH_OR2 C3056 ( .A(N1418), .B(N1420), .Z(N1421) );
  GTECH_AND2 C3057 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[40]), .Z(
        N1418) );
  GTECH_AND2 C3058 ( .A(N1419), .B(a1stg_norm_frac2[40]), .Z(N1420) );
  GTECH_AND2 C3059 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1419) );
  GTECH_AND2 C3061 ( .A(N1422), .B(a1stg_norm_frac1[40]), .Z(N1423) );
  GTECH_AND2 C3062 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1422)
         );
  GTECH_OR2 C3063 ( .A(N1427), .B(N1429), .Z(a2stg_frac2_in[39]) );
  GTECH_OR2 C3064 ( .A(N1424), .B(N1426), .Z(N1427) );
  GTECH_AND2 C3065 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[39]), .Z(
        N1424) );
  GTECH_AND2 C3066 ( .A(N1425), .B(a1stg_norm_frac2[39]), .Z(N1426) );
  GTECH_AND2 C3067 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1425) );
  GTECH_AND2 C3069 ( .A(N1428), .B(a1stg_norm_frac1[39]), .Z(N1429) );
  GTECH_AND2 C3070 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1428)
         );
  GTECH_OR2 C3071 ( .A(N1433), .B(N1435), .Z(a2stg_frac2_in[38]) );
  GTECH_OR2 C3072 ( .A(N1430), .B(N1432), .Z(N1433) );
  GTECH_AND2 C3073 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[38]), .Z(
        N1430) );
  GTECH_AND2 C3074 ( .A(N1431), .B(a1stg_norm_frac2[38]), .Z(N1432) );
  GTECH_AND2 C3075 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1431) );
  GTECH_AND2 C3077 ( .A(N1434), .B(a1stg_norm_frac1[38]), .Z(N1435) );
  GTECH_AND2 C3078 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1434)
         );
  GTECH_OR2 C3079 ( .A(N1439), .B(N1441), .Z(a2stg_frac2_in[37]) );
  GTECH_OR2 C3080 ( .A(N1436), .B(N1438), .Z(N1439) );
  GTECH_AND2 C3081 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[37]), .Z(
        N1436) );
  GTECH_AND2 C3082 ( .A(N1437), .B(a1stg_norm_frac2[37]), .Z(N1438) );
  GTECH_AND2 C3083 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1437) );
  GTECH_AND2 C3085 ( .A(N1440), .B(a1stg_norm_frac1[37]), .Z(N1441) );
  GTECH_AND2 C3086 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1440)
         );
  GTECH_OR2 C3087 ( .A(N1445), .B(N1447), .Z(a2stg_frac2_in[36]) );
  GTECH_OR2 C3088 ( .A(N1442), .B(N1444), .Z(N1445) );
  GTECH_AND2 C3089 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[36]), .Z(
        N1442) );
  GTECH_AND2 C3090 ( .A(N1443), .B(a1stg_norm_frac2[36]), .Z(N1444) );
  GTECH_AND2 C3091 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1443) );
  GTECH_AND2 C3093 ( .A(N1446), .B(a1stg_norm_frac1[36]), .Z(N1447) );
  GTECH_AND2 C3094 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1446)
         );
  GTECH_OR2 C3095 ( .A(N1451), .B(N1453), .Z(a2stg_frac2_in[35]) );
  GTECH_OR2 C3096 ( .A(N1448), .B(N1450), .Z(N1451) );
  GTECH_AND2 C3097 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[35]), .Z(
        N1448) );
  GTECH_AND2 C3098 ( .A(N1449), .B(a1stg_norm_frac2[35]), .Z(N1450) );
  GTECH_AND2 C3099 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1449) );
  GTECH_AND2 C3101 ( .A(N1452), .B(a1stg_norm_frac1[35]), .Z(N1453) );
  GTECH_AND2 C3102 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1452)
         );
  GTECH_OR2 C3103 ( .A(N1457), .B(N1459), .Z(a2stg_frac2_in[34]) );
  GTECH_OR2 C3104 ( .A(N1454), .B(N1456), .Z(N1457) );
  GTECH_AND2 C3105 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[34]), .Z(
        N1454) );
  GTECH_AND2 C3106 ( .A(N1455), .B(a1stg_norm_frac2[34]), .Z(N1456) );
  GTECH_AND2 C3107 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1455) );
  GTECH_AND2 C3109 ( .A(N1458), .B(a1stg_norm_frac1[34]), .Z(N1459) );
  GTECH_AND2 C3110 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1458)
         );
  GTECH_OR2 C3111 ( .A(N1463), .B(N1465), .Z(a2stg_frac2_in[33]) );
  GTECH_OR2 C3112 ( .A(N1460), .B(N1462), .Z(N1463) );
  GTECH_AND2 C3113 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[33]), .Z(
        N1460) );
  GTECH_AND2 C3114 ( .A(N1461), .B(a1stg_norm_frac2[33]), .Z(N1462) );
  GTECH_AND2 C3115 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1461) );
  GTECH_AND2 C3117 ( .A(N1464), .B(a1stg_norm_frac1[33]), .Z(N1465) );
  GTECH_AND2 C3118 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1464)
         );
  GTECH_OR2 C3119 ( .A(N1469), .B(N1471), .Z(a2stg_frac2_in[32]) );
  GTECH_OR2 C3120 ( .A(N1466), .B(N1468), .Z(N1469) );
  GTECH_AND2 C3121 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[32]), .Z(
        N1466) );
  GTECH_AND2 C3122 ( .A(N1467), .B(a1stg_norm_frac2[32]), .Z(N1468) );
  GTECH_AND2 C3123 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1467) );
  GTECH_AND2 C3125 ( .A(N1470), .B(a1stg_norm_frac1[32]), .Z(N1471) );
  GTECH_AND2 C3126 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1470)
         );
  GTECH_OR2 C3127 ( .A(N1475), .B(N1477), .Z(a2stg_frac2_in[31]) );
  GTECH_OR2 C3128 ( .A(N1472), .B(N1474), .Z(N1475) );
  GTECH_AND2 C3129 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[31]), .Z(
        N1472) );
  GTECH_AND2 C3130 ( .A(N1473), .B(a1stg_norm_frac2[31]), .Z(N1474) );
  GTECH_AND2 C3131 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1473) );
  GTECH_AND2 C3133 ( .A(N1476), .B(a1stg_norm_frac1[31]), .Z(N1477) );
  GTECH_AND2 C3134 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1476)
         );
  GTECH_OR2 C3135 ( .A(N1481), .B(N1483), .Z(a2stg_frac2_in[30]) );
  GTECH_OR2 C3136 ( .A(N1478), .B(N1480), .Z(N1481) );
  GTECH_AND2 C3137 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[30]), .Z(
        N1478) );
  GTECH_AND2 C3138 ( .A(N1479), .B(a1stg_norm_frac2[30]), .Z(N1480) );
  GTECH_AND2 C3139 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1479) );
  GTECH_AND2 C3141 ( .A(N1482), .B(a1stg_norm_frac1[30]), .Z(N1483) );
  GTECH_AND2 C3142 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1482)
         );
  GTECH_OR2 C3143 ( .A(N1487), .B(N1489), .Z(a2stg_frac2_in[29]) );
  GTECH_OR2 C3144 ( .A(N1484), .B(N1486), .Z(N1487) );
  GTECH_AND2 C3145 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[29]), .Z(
        N1484) );
  GTECH_AND2 C3146 ( .A(N1485), .B(a1stg_norm_frac2[29]), .Z(N1486) );
  GTECH_AND2 C3147 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1485) );
  GTECH_AND2 C3149 ( .A(N1488), .B(a1stg_norm_frac1[29]), .Z(N1489) );
  GTECH_AND2 C3150 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1488)
         );
  GTECH_OR2 C3151 ( .A(N1493), .B(N1495), .Z(a2stg_frac2_in[28]) );
  GTECH_OR2 C3152 ( .A(N1490), .B(N1492), .Z(N1493) );
  GTECH_AND2 C3153 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[28]), .Z(
        N1490) );
  GTECH_AND2 C3154 ( .A(N1491), .B(a1stg_norm_frac2[28]), .Z(N1492) );
  GTECH_AND2 C3155 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1491) );
  GTECH_AND2 C3157 ( .A(N1494), .B(a1stg_norm_frac1[28]), .Z(N1495) );
  GTECH_AND2 C3158 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1494)
         );
  GTECH_OR2 C3159 ( .A(N1499), .B(N1501), .Z(a2stg_frac2_in[27]) );
  GTECH_OR2 C3160 ( .A(N1496), .B(N1498), .Z(N1499) );
  GTECH_AND2 C3161 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[27]), .Z(
        N1496) );
  GTECH_AND2 C3162 ( .A(N1497), .B(a1stg_norm_frac2[27]), .Z(N1498) );
  GTECH_AND2 C3163 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1497) );
  GTECH_AND2 C3165 ( .A(N1500), .B(a1stg_norm_frac1[27]), .Z(N1501) );
  GTECH_AND2 C3166 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1500)
         );
  GTECH_OR2 C3167 ( .A(N1505), .B(N1507), .Z(a2stg_frac2_in[26]) );
  GTECH_OR2 C3168 ( .A(N1502), .B(N1504), .Z(N1505) );
  GTECH_AND2 C3169 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[26]), .Z(
        N1502) );
  GTECH_AND2 C3170 ( .A(N1503), .B(a1stg_norm_frac2[26]), .Z(N1504) );
  GTECH_AND2 C3171 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1503) );
  GTECH_AND2 C3173 ( .A(N1506), .B(a1stg_norm_frac1[26]), .Z(N1507) );
  GTECH_AND2 C3174 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1506)
         );
  GTECH_OR2 C3175 ( .A(N1511), .B(N1513), .Z(a2stg_frac2_in[25]) );
  GTECH_OR2 C3176 ( .A(N1508), .B(N1510), .Z(N1511) );
  GTECH_AND2 C3177 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[25]), .Z(
        N1508) );
  GTECH_AND2 C3178 ( .A(N1509), .B(a1stg_norm_frac2[25]), .Z(N1510) );
  GTECH_AND2 C3179 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1509) );
  GTECH_AND2 C3181 ( .A(N1512), .B(a1stg_norm_frac1[25]), .Z(N1513) );
  GTECH_AND2 C3182 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1512)
         );
  GTECH_OR2 C3183 ( .A(N1517), .B(N1519), .Z(a2stg_frac2_in[24]) );
  GTECH_OR2 C3184 ( .A(N1514), .B(N1516), .Z(N1517) );
  GTECH_AND2 C3185 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[24]), .Z(
        N1514) );
  GTECH_AND2 C3186 ( .A(N1515), .B(a1stg_norm_frac2[24]), .Z(N1516) );
  GTECH_AND2 C3187 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1515) );
  GTECH_AND2 C3189 ( .A(N1518), .B(a1stg_norm_frac1[24]), .Z(N1519) );
  GTECH_AND2 C3190 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1518)
         );
  GTECH_OR2 C3191 ( .A(N1523), .B(N1525), .Z(a2stg_frac2_in[23]) );
  GTECH_OR2 C3192 ( .A(N1520), .B(N1522), .Z(N1523) );
  GTECH_AND2 C3193 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[23]), .Z(
        N1520) );
  GTECH_AND2 C3194 ( .A(N1521), .B(a1stg_norm_frac2[23]), .Z(N1522) );
  GTECH_AND2 C3195 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1521) );
  GTECH_AND2 C3197 ( .A(N1524), .B(a1stg_norm_frac1[23]), .Z(N1525) );
  GTECH_AND2 C3198 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1524)
         );
  GTECH_OR2 C3199 ( .A(N1529), .B(N1531), .Z(a2stg_frac2_in[22]) );
  GTECH_OR2 C3200 ( .A(N1526), .B(N1528), .Z(N1529) );
  GTECH_AND2 C3201 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[22]), .Z(
        N1526) );
  GTECH_AND2 C3202 ( .A(N1527), .B(a1stg_norm_frac2[22]), .Z(N1528) );
  GTECH_AND2 C3203 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1527) );
  GTECH_AND2 C3205 ( .A(N1530), .B(a1stg_norm_frac1[22]), .Z(N1531) );
  GTECH_AND2 C3206 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1530)
         );
  GTECH_OR2 C3207 ( .A(N1535), .B(N1537), .Z(a2stg_frac2_in[21]) );
  GTECH_OR2 C3208 ( .A(N1532), .B(N1534), .Z(N1535) );
  GTECH_AND2 C3209 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[21]), .Z(
        N1532) );
  GTECH_AND2 C3210 ( .A(N1533), .B(a1stg_norm_frac2[21]), .Z(N1534) );
  GTECH_AND2 C3211 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1533) );
  GTECH_AND2 C3213 ( .A(N1536), .B(a1stg_norm_frac1[21]), .Z(N1537) );
  GTECH_AND2 C3214 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1536)
         );
  GTECH_OR2 C3215 ( .A(N1541), .B(N1543), .Z(a2stg_frac2_in[20]) );
  GTECH_OR2 C3216 ( .A(N1538), .B(N1540), .Z(N1541) );
  GTECH_AND2 C3217 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[20]), .Z(
        N1538) );
  GTECH_AND2 C3218 ( .A(N1539), .B(a1stg_norm_frac2[20]), .Z(N1540) );
  GTECH_AND2 C3219 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1539) );
  GTECH_AND2 C3221 ( .A(N1542), .B(a1stg_norm_frac1[20]), .Z(N1543) );
  GTECH_AND2 C3222 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1542)
         );
  GTECH_OR2 C3223 ( .A(N1547), .B(N1549), .Z(a2stg_frac2_in[19]) );
  GTECH_OR2 C3224 ( .A(N1544), .B(N1546), .Z(N1547) );
  GTECH_AND2 C3225 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[19]), .Z(
        N1544) );
  GTECH_AND2 C3226 ( .A(N1545), .B(a1stg_norm_frac2[19]), .Z(N1546) );
  GTECH_AND2 C3227 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1545) );
  GTECH_AND2 C3229 ( .A(N1548), .B(a1stg_norm_frac1[19]), .Z(N1549) );
  GTECH_AND2 C3230 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1548)
         );
  GTECH_OR2 C3231 ( .A(N1553), .B(N1555), .Z(a2stg_frac2_in[18]) );
  GTECH_OR2 C3232 ( .A(N1550), .B(N1552), .Z(N1553) );
  GTECH_AND2 C3233 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[18]), .Z(
        N1550) );
  GTECH_AND2 C3234 ( .A(N1551), .B(a1stg_norm_frac2[18]), .Z(N1552) );
  GTECH_AND2 C3235 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1551) );
  GTECH_AND2 C3237 ( .A(N1554), .B(a1stg_norm_frac1[18]), .Z(N1555) );
  GTECH_AND2 C3238 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1554)
         );
  GTECH_OR2 C3239 ( .A(N1559), .B(N1561), .Z(a2stg_frac2_in[17]) );
  GTECH_OR2 C3240 ( .A(N1556), .B(N1558), .Z(N1559) );
  GTECH_AND2 C3241 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[17]), .Z(
        N1556) );
  GTECH_AND2 C3242 ( .A(N1557), .B(a1stg_norm_frac2[17]), .Z(N1558) );
  GTECH_AND2 C3243 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1557) );
  GTECH_AND2 C3245 ( .A(N1560), .B(a1stg_norm_frac1[17]), .Z(N1561) );
  GTECH_AND2 C3246 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1560)
         );
  GTECH_OR2 C3247 ( .A(N1565), .B(N1567), .Z(a2stg_frac2_in[16]) );
  GTECH_OR2 C3248 ( .A(N1562), .B(N1564), .Z(N1565) );
  GTECH_AND2 C3249 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[16]), .Z(
        N1562) );
  GTECH_AND2 C3250 ( .A(N1563), .B(a1stg_norm_frac2[16]), .Z(N1564) );
  GTECH_AND2 C3251 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1563) );
  GTECH_AND2 C3253 ( .A(N1566), .B(a1stg_norm_frac1[16]), .Z(N1567) );
  GTECH_AND2 C3254 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1566)
         );
  GTECH_OR2 C3255 ( .A(N1571), .B(N1573), .Z(a2stg_frac2_in[15]) );
  GTECH_OR2 C3256 ( .A(N1568), .B(N1570), .Z(N1571) );
  GTECH_AND2 C3257 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[15]), .Z(
        N1568) );
  GTECH_AND2 C3258 ( .A(N1569), .B(a1stg_norm_frac2[15]), .Z(N1570) );
  GTECH_AND2 C3259 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1569) );
  GTECH_AND2 C3261 ( .A(N1572), .B(a1stg_norm_frac1[15]), .Z(N1573) );
  GTECH_AND2 C3262 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1572)
         );
  GTECH_OR2 C3263 ( .A(N1577), .B(N1579), .Z(a2stg_frac2_in[14]) );
  GTECH_OR2 C3264 ( .A(N1574), .B(N1576), .Z(N1577) );
  GTECH_AND2 C3265 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[14]), .Z(
        N1574) );
  GTECH_AND2 C3266 ( .A(N1575), .B(a1stg_norm_frac2[14]), .Z(N1576) );
  GTECH_AND2 C3267 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1575) );
  GTECH_AND2 C3269 ( .A(N1578), .B(a1stg_norm_frac1[14]), .Z(N1579) );
  GTECH_AND2 C3270 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1578)
         );
  GTECH_OR2 C3271 ( .A(N1583), .B(N1585), .Z(a2stg_frac2_in[13]) );
  GTECH_OR2 C3272 ( .A(N1580), .B(N1582), .Z(N1583) );
  GTECH_AND2 C3273 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[13]), .Z(
        N1580) );
  GTECH_AND2 C3274 ( .A(N1581), .B(a1stg_norm_frac2[13]), .Z(N1582) );
  GTECH_AND2 C3275 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1581) );
  GTECH_AND2 C3277 ( .A(N1584), .B(a1stg_norm_frac1[13]), .Z(N1585) );
  GTECH_AND2 C3278 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1584)
         );
  GTECH_OR2 C3279 ( .A(N1589), .B(N1591), .Z(a2stg_frac2_in[12]) );
  GTECH_OR2 C3280 ( .A(N1586), .B(N1588), .Z(N1589) );
  GTECH_AND2 C3281 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[12]), .Z(
        N1586) );
  GTECH_AND2 C3282 ( .A(N1587), .B(a1stg_norm_frac2[12]), .Z(N1588) );
  GTECH_AND2 C3283 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1587) );
  GTECH_AND2 C3285 ( .A(N1590), .B(a1stg_norm_frac1[12]), .Z(N1591) );
  GTECH_AND2 C3286 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1590)
         );
  GTECH_OR2 C3287 ( .A(N1595), .B(N1597), .Z(a2stg_frac2_in[11]) );
  GTECH_OR2 C3288 ( .A(N1592), .B(N1594), .Z(N1595) );
  GTECH_AND2 C3289 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[11]), .Z(
        N1592) );
  GTECH_AND2 C3290 ( .A(N1593), .B(a1stg_norm_frac2[11]), .Z(N1594) );
  GTECH_AND2 C3291 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1593) );
  GTECH_AND2 C3293 ( .A(N1596), .B(a1stg_norm_frac1[11]), .Z(N1597) );
  GTECH_AND2 C3294 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1596)
         );
  GTECH_OR2 C3295 ( .A(N1601), .B(N1603), .Z(a2stg_frac2_in[10]) );
  GTECH_OR2 C3296 ( .A(N1598), .B(N1600), .Z(N1601) );
  GTECH_AND2 C3297 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[10]), .Z(
        N1598) );
  GTECH_AND2 C3298 ( .A(N1599), .B(a1stg_norm_frac2[10]), .Z(N1600) );
  GTECH_AND2 C3299 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1599) );
  GTECH_AND2 C3301 ( .A(N1602), .B(1'b0), .Z(N1603) );
  GTECH_AND2 C3302 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1602)
         );
  GTECH_OR2 C3303 ( .A(N1607), .B(N1609), .Z(a2stg_frac2_in[9]) );
  GTECH_OR2 C3304 ( .A(N1604), .B(N1606), .Z(N1607) );
  GTECH_AND2 C3305 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[9]), .Z(
        N1604) );
  GTECH_AND2 C3306 ( .A(N1605), .B(a1stg_norm_frac2[9]), .Z(N1606) );
  GTECH_AND2 C3307 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1605) );
  GTECH_AND2 C3309 ( .A(N1608), .B(1'b0), .Z(N1609) );
  GTECH_AND2 C3310 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1608)
         );
  GTECH_OR2 C3311 ( .A(N1613), .B(N1615), .Z(a2stg_frac2_in[8]) );
  GTECH_OR2 C3312 ( .A(N1610), .B(N1612), .Z(N1613) );
  GTECH_AND2 C3313 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[8]), .Z(
        N1610) );
  GTECH_AND2 C3314 ( .A(N1611), .B(a1stg_norm_frac2[8]), .Z(N1612) );
  GTECH_AND2 C3315 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1611) );
  GTECH_AND2 C3317 ( .A(N1614), .B(1'b0), .Z(N1615) );
  GTECH_AND2 C3318 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1614)
         );
  GTECH_OR2 C3319 ( .A(N1619), .B(N1621), .Z(a2stg_frac2_in[7]) );
  GTECH_OR2 C3320 ( .A(N1616), .B(N1618), .Z(N1619) );
  GTECH_AND2 C3321 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[7]), .Z(
        N1616) );
  GTECH_AND2 C3322 ( .A(N1617), .B(a1stg_norm_frac2[7]), .Z(N1618) );
  GTECH_AND2 C3323 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1617) );
  GTECH_AND2 C3325 ( .A(N1620), .B(1'b0), .Z(N1621) );
  GTECH_AND2 C3326 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1620)
         );
  GTECH_OR2 C3327 ( .A(N1625), .B(N1627), .Z(a2stg_frac2_in[6]) );
  GTECH_OR2 C3328 ( .A(N1622), .B(N1624), .Z(N1625) );
  GTECH_AND2 C3329 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[6]), .Z(
        N1622) );
  GTECH_AND2 C3330 ( .A(N1623), .B(a1stg_norm_frac2[6]), .Z(N1624) );
  GTECH_AND2 C3331 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1623) );
  GTECH_AND2 C3333 ( .A(N1626), .B(1'b0), .Z(N1627) );
  GTECH_AND2 C3334 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1626)
         );
  GTECH_OR2 C3335 ( .A(N1631), .B(N1633), .Z(a2stg_frac2_in[5]) );
  GTECH_OR2 C3336 ( .A(N1628), .B(N1630), .Z(N1631) );
  GTECH_AND2 C3337 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[5]), .Z(
        N1628) );
  GTECH_AND2 C3338 ( .A(N1629), .B(a1stg_norm_frac2[5]), .Z(N1630) );
  GTECH_AND2 C3339 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1629) );
  GTECH_AND2 C3341 ( .A(N1632), .B(1'b0), .Z(N1633) );
  GTECH_AND2 C3342 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1632)
         );
  GTECH_OR2 C3343 ( .A(N1637), .B(N1639), .Z(a2stg_frac2_in[4]) );
  GTECH_OR2 C3344 ( .A(N1634), .B(N1636), .Z(N1637) );
  GTECH_AND2 C3345 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[4]), .Z(
        N1634) );
  GTECH_AND2 C3346 ( .A(N1635), .B(a1stg_norm_frac2[4]), .Z(N1636) );
  GTECH_AND2 C3347 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1635) );
  GTECH_AND2 C3349 ( .A(N1638), .B(1'b0), .Z(N1639) );
  GTECH_AND2 C3350 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1638)
         );
  GTECH_OR2 C3351 ( .A(N1643), .B(N1645), .Z(a2stg_frac2_in[3]) );
  GTECH_OR2 C3352 ( .A(N1640), .B(N1642), .Z(N1643) );
  GTECH_AND2 C3353 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[3]), .Z(
        N1640) );
  GTECH_AND2 C3354 ( .A(N1641), .B(a1stg_norm_frac2[3]), .Z(N1642) );
  GTECH_AND2 C3355 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1641) );
  GTECH_AND2 C3357 ( .A(N1644), .B(1'b0), .Z(N1645) );
  GTECH_AND2 C3358 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1644)
         );
  GTECH_OR2 C3359 ( .A(N1649), .B(N1651), .Z(a2stg_frac2_in[2]) );
  GTECH_OR2 C3360 ( .A(N1646), .B(N1648), .Z(N1649) );
  GTECH_AND2 C3361 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[2]), .Z(
        N1646) );
  GTECH_AND2 C3362 ( .A(N1647), .B(a1stg_norm_frac2[2]), .Z(N1648) );
  GTECH_AND2 C3363 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1647) );
  GTECH_AND2 C3365 ( .A(N1650), .B(1'b0), .Z(N1651) );
  GTECH_AND2 C3366 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1650)
         );
  GTECH_OR2 C3367 ( .A(N1655), .B(N1657), .Z(a2stg_frac2_in[1]) );
  GTECH_OR2 C3368 ( .A(N1652), .B(N1654), .Z(N1655) );
  GTECH_AND2 C3369 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[1]), .Z(
        N1652) );
  GTECH_AND2 C3370 ( .A(N1653), .B(a1stg_norm_frac2[1]), .Z(N1654) );
  GTECH_AND2 C3371 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1653) );
  GTECH_AND2 C3373 ( .A(N1656), .B(1'b0), .Z(N1657) );
  GTECH_AND2 C3374 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1656)
         );
  GTECH_OR2 C3375 ( .A(N1661), .B(N1663), .Z(a2stg_frac2_in[0]) );
  GTECH_OR2 C3376 ( .A(N1658), .B(N1660), .Z(N1661) );
  GTECH_AND2 C3377 ( .A(a1stg_faddsubop_inv), .B(a1stg_norm_frac2[0]), .Z(
        N1658) );
  GTECH_AND2 C3378 ( .A(N1659), .B(a1stg_norm_frac2[0]), .Z(N1660) );
  GTECH_AND2 C3379 ( .A(a2stg_frac2_in_frac1), .B(N1280), .Z(N1659) );
  GTECH_AND2 C3381 ( .A(N1662), .B(1'b0), .Z(N1663) );
  GTECH_AND2 C3382 ( .A(a2stg_frac2_in_frac1), .B(a1stg_in2_gt_in1), .Z(N1662)
         );
  GTECH_OR2 C3383 ( .A(N1692), .B(a2stg_frac2[32]), .Z(a2stg_frac2hi_neq_0) );
  GTECH_OR2 C3384 ( .A(N1691), .B(a2stg_frac2[33]), .Z(N1692) );
  GTECH_OR2 C3385 ( .A(N1690), .B(a2stg_frac2[34]), .Z(N1691) );
  GTECH_OR2 C3386 ( .A(N1689), .B(a2stg_frac2[35]), .Z(N1690) );
  GTECH_OR2 C3387 ( .A(N1688), .B(a2stg_frac2[36]), .Z(N1689) );
  GTECH_OR2 C3388 ( .A(N1687), .B(a2stg_frac2[37]), .Z(N1688) );
  GTECH_OR2 C3389 ( .A(N1686), .B(a2stg_frac2[38]), .Z(N1687) );
  GTECH_OR2 C3390 ( .A(N1685), .B(a2stg_frac2[39]), .Z(N1686) );
  GTECH_OR2 C3391 ( .A(N1684), .B(a2stg_frac2[40]), .Z(N1685) );
  GTECH_OR2 C3392 ( .A(N1683), .B(a2stg_frac2[41]), .Z(N1684) );
  GTECH_OR2 C3393 ( .A(N1682), .B(a2stg_frac2[42]), .Z(N1683) );
  GTECH_OR2 C3394 ( .A(N1681), .B(a2stg_frac2[43]), .Z(N1682) );
  GTECH_OR2 C3395 ( .A(N1680), .B(a2stg_frac2[44]), .Z(N1681) );
  GTECH_OR2 C3396 ( .A(N1679), .B(a2stg_frac2[45]), .Z(N1680) );
  GTECH_OR2 C3397 ( .A(N1678), .B(a2stg_frac2[46]), .Z(N1679) );
  GTECH_OR2 C3398 ( .A(N1677), .B(a2stg_frac2[47]), .Z(N1678) );
  GTECH_OR2 C3399 ( .A(N1676), .B(a2stg_frac2[48]), .Z(N1677) );
  GTECH_OR2 C3400 ( .A(N1675), .B(a2stg_frac2[49]), .Z(N1676) );
  GTECH_OR2 C3401 ( .A(N1674), .B(a2stg_frac2[50]), .Z(N1675) );
  GTECH_OR2 C3402 ( .A(N1673), .B(a2stg_frac2[51]), .Z(N1674) );
  GTECH_OR2 C3403 ( .A(N1672), .B(a2stg_frac2[52]), .Z(N1673) );
  GTECH_OR2 C3404 ( .A(N1671), .B(a2stg_frac2[53]), .Z(N1672) );
  GTECH_OR2 C3405 ( .A(N1670), .B(a2stg_frac2[54]), .Z(N1671) );
  GTECH_OR2 C3406 ( .A(N1669), .B(a2stg_frac2[55]), .Z(N1670) );
  GTECH_OR2 C3407 ( .A(N1668), .B(a2stg_frac2[56]), .Z(N1669) );
  GTECH_OR2 C3408 ( .A(N1667), .B(a2stg_frac2[57]), .Z(N1668) );
  GTECH_OR2 C3409 ( .A(N1666), .B(a2stg_frac2[58]), .Z(N1667) );
  GTECH_OR2 C3410 ( .A(N1665), .B(a2stg_frac2[59]), .Z(N1666) );
  GTECH_OR2 C3411 ( .A(N1664), .B(a2stg_frac2[60]), .Z(N1665) );
  GTECH_OR2 C3412 ( .A(a2stg_frac2[62]), .B(a2stg_frac2[61]), .Z(N1664) );
  GTECH_OR2 C3413 ( .A(N1711), .B(a2stg_frac2[11]), .Z(a2stg_frac2lo_neq_0) );
  GTECH_OR2 C3414 ( .A(N1710), .B(a2stg_frac2[12]), .Z(N1711) );
  GTECH_OR2 C3415 ( .A(N1709), .B(a2stg_frac2[13]), .Z(N1710) );
  GTECH_OR2 C3416 ( .A(N1708), .B(a2stg_frac2[14]), .Z(N1709) );
  GTECH_OR2 C3417 ( .A(N1707), .B(a2stg_frac2[15]), .Z(N1708) );
  GTECH_OR2 C3418 ( .A(N1706), .B(a2stg_frac2[16]), .Z(N1707) );
  GTECH_OR2 C3419 ( .A(N1705), .B(a2stg_frac2[17]), .Z(N1706) );
  GTECH_OR2 C3420 ( .A(N1704), .B(a2stg_frac2[18]), .Z(N1705) );
  GTECH_OR2 C3421 ( .A(N1703), .B(a2stg_frac2[19]), .Z(N1704) );
  GTECH_OR2 C3422 ( .A(N1702), .B(a2stg_frac2[20]), .Z(N1703) );
  GTECH_OR2 C3423 ( .A(N1701), .B(a2stg_frac2[21]), .Z(N1702) );
  GTECH_OR2 C3424 ( .A(N1700), .B(a2stg_frac2[22]), .Z(N1701) );
  GTECH_OR2 C3425 ( .A(N1699), .B(a2stg_frac2[23]), .Z(N1700) );
  GTECH_OR2 C3426 ( .A(N1698), .B(a2stg_frac2[24]), .Z(N1699) );
  GTECH_OR2 C3427 ( .A(N1697), .B(a2stg_frac2[25]), .Z(N1698) );
  GTECH_OR2 C3428 ( .A(N1696), .B(a2stg_frac2[26]), .Z(N1697) );
  GTECH_OR2 C3429 ( .A(N1695), .B(a2stg_frac2[27]), .Z(N1696) );
  GTECH_OR2 C3430 ( .A(N1694), .B(a2stg_frac2[28]), .Z(N1695) );
  GTECH_OR2 C3431 ( .A(N1693), .B(a2stg_frac2[29]), .Z(N1694) );
  GTECH_OR2 C3432 ( .A(a2stg_frac2[31]), .B(a2stg_frac2[30]), .Z(N1693) );
  GTECH_AND2 C3433 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[63]), .Z(
        a2stg_shr_tmp2[63]) );
  GTECH_AND2 C3434 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[62]), .Z(
        a2stg_shr_tmp2[62]) );
  GTECH_AND2 C3435 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[61]), .Z(
        a2stg_shr_tmp2[61]) );
  GTECH_AND2 C3436 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[60]), .Z(
        a2stg_shr_tmp2[60]) );
  GTECH_AND2 C3437 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[59]), .Z(
        a2stg_shr_tmp2[59]) );
  GTECH_AND2 C3438 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[58]), .Z(
        a2stg_shr_tmp2[58]) );
  GTECH_AND2 C3439 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[57]), .Z(
        a2stg_shr_tmp2[57]) );
  GTECH_AND2 C3440 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[56]), .Z(
        a2stg_shr_tmp2[56]) );
  GTECH_AND2 C3441 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[55]), .Z(
        a2stg_shr_tmp2[55]) );
  GTECH_AND2 C3442 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[54]), .Z(
        a2stg_shr_tmp2[54]) );
  GTECH_AND2 C3443 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[53]), .Z(
        a2stg_shr_tmp2[53]) );
  GTECH_AND2 C3444 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[52]), .Z(
        a2stg_shr_tmp2[52]) );
  GTECH_AND2 C3445 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[51]), .Z(
        a2stg_shr_tmp2[51]) );
  GTECH_AND2 C3446 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[50]), .Z(
        a2stg_shr_tmp2[50]) );
  GTECH_AND2 C3447 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[49]), .Z(
        a2stg_shr_tmp2[49]) );
  GTECH_AND2 C3448 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[48]), .Z(
        a2stg_shr_tmp2[48]) );
  GTECH_AND2 C3449 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[47]), .Z(
        a2stg_shr_tmp2[47]) );
  GTECH_AND2 C3450 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[46]), .Z(
        a2stg_shr_tmp2[46]) );
  GTECH_AND2 C3451 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[45]), .Z(
        a2stg_shr_tmp2[45]) );
  GTECH_AND2 C3452 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[44]), .Z(
        a2stg_shr_tmp2[44]) );
  GTECH_AND2 C3453 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[43]), .Z(
        a2stg_shr_tmp2[43]) );
  GTECH_AND2 C3454 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[42]), .Z(
        a2stg_shr_tmp2[42]) );
  GTECH_AND2 C3455 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[41]), .Z(
        a2stg_shr_tmp2[41]) );
  GTECH_AND2 C3456 ( .A(a2stg_shr_cnt_5_inv[0]), .B(a2stg_frac2a[40]), .Z(
        a2stg_shr_tmp2[40]) );
  GTECH_AND2 C3457 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[39]), .Z(
        a2stg_shr_tmp2[39]) );
  GTECH_AND2 C3458 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[38]), .Z(
        a2stg_shr_tmp2[38]) );
  GTECH_AND2 C3459 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[37]), .Z(
        a2stg_shr_tmp2[37]) );
  GTECH_AND2 C3460 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[36]), .Z(
        a2stg_shr_tmp2[36]) );
  GTECH_AND2 C3461 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[35]), .Z(
        a2stg_shr_tmp2[35]) );
  GTECH_AND2 C3462 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[34]), .Z(
        a2stg_shr_tmp2[34]) );
  GTECH_AND2 C3463 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[33]), .Z(
        a2stg_shr_tmp2[33]) );
  GTECH_AND2 C3464 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[32]), .Z(
        a2stg_shr_tmp2[32]) );
  GTECH_OR2 C3465 ( .A(N1712), .B(N1713), .Z(a2stg_shr_tmp2[31]) );
  GTECH_AND2 C3466 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[63]), .Z(N1712)
         );
  GTECH_AND2 C3467 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[31]), .Z(
        N1713) );
  GTECH_OR2 C3468 ( .A(N1714), .B(N1715), .Z(a2stg_shr_tmp2[30]) );
  GTECH_AND2 C3469 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[62]), .Z(N1714)
         );
  GTECH_AND2 C3470 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[30]), .Z(
        N1715) );
  GTECH_OR2 C3471 ( .A(N1716), .B(N1717), .Z(a2stg_shr_tmp2[29]) );
  GTECH_AND2 C3472 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[61]), .Z(N1716)
         );
  GTECH_AND2 C3473 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[29]), .Z(
        N1717) );
  GTECH_OR2 C3474 ( .A(N1718), .B(N1719), .Z(a2stg_shr_tmp2[28]) );
  GTECH_AND2 C3475 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[60]), .Z(N1718)
         );
  GTECH_AND2 C3476 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[28]), .Z(
        N1719) );
  GTECH_OR2 C3477 ( .A(N1720), .B(N1721), .Z(a2stg_shr_tmp2[27]) );
  GTECH_AND2 C3478 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[59]), .Z(N1720)
         );
  GTECH_AND2 C3479 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[27]), .Z(
        N1721) );
  GTECH_OR2 C3480 ( .A(N1722), .B(N1723), .Z(a2stg_shr_tmp2[26]) );
  GTECH_AND2 C3481 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[58]), .Z(N1722)
         );
  GTECH_AND2 C3482 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[26]), .Z(
        N1723) );
  GTECH_OR2 C3483 ( .A(N1724), .B(N1725), .Z(a2stg_shr_tmp2[25]) );
  GTECH_AND2 C3484 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[57]), .Z(N1724)
         );
  GTECH_AND2 C3485 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[25]), .Z(
        N1725) );
  GTECH_OR2 C3486 ( .A(N1726), .B(N1727), .Z(a2stg_shr_tmp2[24]) );
  GTECH_AND2 C3487 ( .A(a2stg_shr_cnt_5[1]), .B(a2stg_frac2a[56]), .Z(N1726)
         );
  GTECH_AND2 C3488 ( .A(a2stg_shr_cnt_5_inv[1]), .B(a2stg_frac2a[24]), .Z(
        N1727) );
  GTECH_OR2 C3489 ( .A(N1728), .B(N1729), .Z(a2stg_shr_tmp2[23]) );
  GTECH_AND2 C3490 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[55]), .Z(N1728)
         );
  GTECH_AND2 C3491 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[23]), .Z(
        N1729) );
  GTECH_OR2 C3492 ( .A(N1730), .B(N1731), .Z(a2stg_shr_tmp2[22]) );
  GTECH_AND2 C3493 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[54]), .Z(N1730)
         );
  GTECH_AND2 C3494 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[22]), .Z(
        N1731) );
  GTECH_OR2 C3495 ( .A(N1732), .B(N1733), .Z(a2stg_shr_tmp2[21]) );
  GTECH_AND2 C3496 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[53]), .Z(N1732)
         );
  GTECH_AND2 C3497 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[21]), .Z(
        N1733) );
  GTECH_OR2 C3498 ( .A(N1734), .B(N1735), .Z(a2stg_shr_tmp2[20]) );
  GTECH_AND2 C3499 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[52]), .Z(N1734)
         );
  GTECH_AND2 C3500 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[20]), .Z(
        N1735) );
  GTECH_OR2 C3501 ( .A(N1736), .B(N1737), .Z(a2stg_shr_tmp2[19]) );
  GTECH_AND2 C3502 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[51]), .Z(N1736)
         );
  GTECH_AND2 C3503 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[19]), .Z(
        N1737) );
  GTECH_OR2 C3504 ( .A(N1738), .B(N1739), .Z(a2stg_shr_tmp2[18]) );
  GTECH_AND2 C3505 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[50]), .Z(N1738)
         );
  GTECH_AND2 C3506 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[18]), .Z(
        N1739) );
  GTECH_OR2 C3507 ( .A(N1740), .B(N1741), .Z(a2stg_shr_tmp2[17]) );
  GTECH_AND2 C3508 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[49]), .Z(N1740)
         );
  GTECH_AND2 C3509 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[17]), .Z(
        N1741) );
  GTECH_OR2 C3510 ( .A(N1742), .B(N1743), .Z(a2stg_shr_tmp2[16]) );
  GTECH_AND2 C3511 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[48]), .Z(N1742)
         );
  GTECH_AND2 C3512 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[16]), .Z(
        N1743) );
  GTECH_OR2 C3513 ( .A(N1744), .B(N1745), .Z(a2stg_shr_tmp2[15]) );
  GTECH_AND2 C3514 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[47]), .Z(N1744)
         );
  GTECH_AND2 C3515 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[15]), .Z(
        N1745) );
  GTECH_OR2 C3516 ( .A(N1746), .B(N1747), .Z(a2stg_shr_tmp2[14]) );
  GTECH_AND2 C3517 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[46]), .Z(N1746)
         );
  GTECH_AND2 C3518 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[14]), .Z(
        N1747) );
  GTECH_OR2 C3519 ( .A(N1748), .B(N1749), .Z(a2stg_shr_tmp2[13]) );
  GTECH_AND2 C3520 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[45]), .Z(N1748)
         );
  GTECH_AND2 C3521 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[13]), .Z(
        N1749) );
  GTECH_OR2 C3522 ( .A(N1750), .B(N1751), .Z(a2stg_shr_tmp2[12]) );
  GTECH_AND2 C3523 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[44]), .Z(N1750)
         );
  GTECH_AND2 C3524 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[12]), .Z(
        N1751) );
  GTECH_OR2 C3525 ( .A(N1752), .B(N1753), .Z(a2stg_shr_tmp2[11]) );
  GTECH_AND2 C3526 ( .A(a2stg_shr_cnt_5[2]), .B(a2stg_frac2a[43]), .Z(N1752)
         );
  GTECH_AND2 C3527 ( .A(a2stg_shr_cnt_5_inv[2]), .B(a2stg_frac2a[11]), .Z(
        N1753) );
  GTECH_OR2 C3528 ( .A(N1754), .B(N1755), .Z(a2stg_shr_tmp2[10]) );
  GTECH_AND2 C3529 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[42]), .Z(N1754)
         );
  GTECH_AND2 C3530 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[10]), .Z(
        N1755) );
  GTECH_OR2 C3531 ( .A(N1756), .B(N1757), .Z(a2stg_shr_tmp2[9]) );
  GTECH_AND2 C3532 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[41]), .Z(N1756)
         );
  GTECH_AND2 C3533 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[9]), .Z(N1757) );
  GTECH_OR2 C3534 ( .A(N1758), .B(N1759), .Z(a2stg_shr_tmp2[8]) );
  GTECH_AND2 C3535 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[40]), .Z(N1758)
         );
  GTECH_AND2 C3536 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[8]), .Z(N1759) );
  GTECH_OR2 C3537 ( .A(N1760), .B(N1761), .Z(a2stg_shr_tmp2[7]) );
  GTECH_AND2 C3538 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[39]), .Z(N1760)
         );
  GTECH_AND2 C3539 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[7]), .Z(N1761) );
  GTECH_OR2 C3540 ( .A(N1762), .B(N1763), .Z(a2stg_shr_tmp2[6]) );
  GTECH_AND2 C3541 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[38]), .Z(N1762)
         );
  GTECH_AND2 C3542 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[6]), .Z(N1763) );
  GTECH_OR2 C3543 ( .A(N1764), .B(N1765), .Z(a2stg_shr_tmp2[5]) );
  GTECH_AND2 C3544 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[37]), .Z(N1764)
         );
  GTECH_AND2 C3545 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[5]), .Z(N1765) );
  GTECH_OR2 C3546 ( .A(N1766), .B(N1767), .Z(a2stg_shr_tmp2[4]) );
  GTECH_AND2 C3547 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[36]), .Z(N1766)
         );
  GTECH_AND2 C3548 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[4]), .Z(N1767) );
  GTECH_OR2 C3549 ( .A(N1768), .B(N1769), .Z(a2stg_shr_tmp2[3]) );
  GTECH_AND2 C3550 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[35]), .Z(N1768)
         );
  GTECH_AND2 C3551 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[3]), .Z(N1769) );
  GTECH_OR2 C3552 ( .A(N1770), .B(N1771), .Z(a2stg_shr_tmp2[2]) );
  GTECH_AND2 C3553 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[34]), .Z(N1770)
         );
  GTECH_AND2 C3554 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[2]), .Z(N1771) );
  GTECH_OR2 C3555 ( .A(N1772), .B(N1773), .Z(a2stg_shr_tmp2[1]) );
  GTECH_AND2 C3556 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[33]), .Z(N1772)
         );
  GTECH_AND2 C3557 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[1]), .Z(N1773) );
  GTECH_OR2 C3558 ( .A(N1774), .B(N1775), .Z(a2stg_shr_tmp2[0]) );
  GTECH_AND2 C3559 ( .A(a2stg_shr_cnt_5[3]), .B(a2stg_frac2a[32]), .Z(N1774)
         );
  GTECH_AND2 C3560 ( .A(a2stg_shr_cnt_5_inv[3]), .B(a2stg_frac2a[0]), .Z(N1775) );
  GTECH_NOT I_77 ( .A(a2stg_shr_cnt_4[4]), .Z(N1) );
  GTECH_AND2 C3562 ( .A(N1), .B(a2stg_shr_tmp2[63]), .Z(a2stg_shr_tmp4[63]) );
  GTECH_AND2 C3563 ( .A(N1), .B(a2stg_shr_tmp2[62]), .Z(a2stg_shr_tmp4[62]) );
  GTECH_AND2 C3564 ( .A(N1), .B(a2stg_shr_tmp2[61]), .Z(a2stg_shr_tmp4[61]) );
  GTECH_AND2 C3565 ( .A(N1), .B(a2stg_shr_tmp2[60]), .Z(a2stg_shr_tmp4[60]) );
  GTECH_AND2 C3566 ( .A(N1), .B(a2stg_shr_tmp2[59]), .Z(a2stg_shr_tmp4[59]) );
  GTECH_AND2 C3567 ( .A(N1), .B(a2stg_shr_tmp2[58]), .Z(a2stg_shr_tmp4[58]) );
  GTECH_AND2 C3568 ( .A(N1), .B(a2stg_shr_tmp2[57]), .Z(a2stg_shr_tmp4[57]) );
  GTECH_AND2 C3569 ( .A(N1), .B(a2stg_shr_tmp2[56]), .Z(a2stg_shr_tmp4[56]) );
  GTECH_AND2 C3570 ( .A(N1), .B(a2stg_shr_tmp2[55]), .Z(a2stg_shr_tmp4[55]) );
  GTECH_AND2 C3571 ( .A(N1), .B(a2stg_shr_tmp2[54]), .Z(a2stg_shr_tmp4[54]) );
  GTECH_AND2 C3572 ( .A(N1), .B(a2stg_shr_tmp2[53]), .Z(a2stg_shr_tmp4[53]) );
  GTECH_AND2 C3573 ( .A(N1), .B(a2stg_shr_tmp2[52]), .Z(a2stg_shr_tmp4[52]) );
  GTECH_AND2 C3574 ( .A(N1), .B(a2stg_shr_tmp2[51]), .Z(a2stg_shr_tmp4[51]) );
  GTECH_AND2 C3575 ( .A(N1), .B(a2stg_shr_tmp2[50]), .Z(a2stg_shr_tmp4[50]) );
  GTECH_AND2 C3576 ( .A(N1), .B(a2stg_shr_tmp2[49]), .Z(a2stg_shr_tmp4[49]) );
  GTECH_AND2 C3577 ( .A(N1), .B(a2stg_shr_tmp2[48]), .Z(a2stg_shr_tmp4[48]) );
  GTECH_OR2 C3578 ( .A(N1776), .B(N1777), .Z(a2stg_shr_tmp4[47]) );
  GTECH_AND2 C3579 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[63]), .Z(N1776)
         );
  GTECH_AND2 C3580 ( .A(N1), .B(a2stg_shr_tmp2[47]), .Z(N1777) );
  GTECH_OR2 C3581 ( .A(N1778), .B(N1779), .Z(a2stg_shr_tmp4[46]) );
  GTECH_AND2 C3582 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[62]), .Z(N1778)
         );
  GTECH_AND2 C3583 ( .A(N1), .B(a2stg_shr_tmp2[46]), .Z(N1779) );
  GTECH_OR2 C3584 ( .A(N1780), .B(N1781), .Z(a2stg_shr_tmp4[45]) );
  GTECH_AND2 C3585 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[61]), .Z(N1780)
         );
  GTECH_AND2 C3586 ( .A(N1), .B(a2stg_shr_tmp2[45]), .Z(N1781) );
  GTECH_OR2 C3587 ( .A(N1782), .B(N1783), .Z(a2stg_shr_tmp4[44]) );
  GTECH_AND2 C3588 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[60]), .Z(N1782)
         );
  GTECH_AND2 C3589 ( .A(N1), .B(a2stg_shr_tmp2[44]), .Z(N1783) );
  GTECH_OR2 C3590 ( .A(N1784), .B(N1785), .Z(a2stg_shr_tmp4[43]) );
  GTECH_AND2 C3591 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[59]), .Z(N1784)
         );
  GTECH_AND2 C3592 ( .A(N1), .B(a2stg_shr_tmp2[43]), .Z(N1785) );
  GTECH_OR2 C3593 ( .A(N1786), .B(N1787), .Z(a2stg_shr_tmp4[42]) );
  GTECH_AND2 C3594 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[58]), .Z(N1786)
         );
  GTECH_AND2 C3595 ( .A(N1), .B(a2stg_shr_tmp2[42]), .Z(N1787) );
  GTECH_OR2 C3596 ( .A(N1788), .B(N1789), .Z(a2stg_shr_tmp4[41]) );
  GTECH_AND2 C3597 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[57]), .Z(N1788)
         );
  GTECH_AND2 C3598 ( .A(N1), .B(a2stg_shr_tmp2[41]), .Z(N1789) );
  GTECH_OR2 C3599 ( .A(N1790), .B(N1791), .Z(a2stg_shr_tmp4[40]) );
  GTECH_AND2 C3600 ( .A(a2stg_shr_cnt_4[0]), .B(a2stg_shr_tmp2[56]), .Z(N1790)
         );
  GTECH_AND2 C3601 ( .A(N1), .B(a2stg_shr_tmp2[40]), .Z(N1791) );
  GTECH_OR2 C3602 ( .A(N1792), .B(N1793), .Z(a2stg_shr_tmp4[39]) );
  GTECH_AND2 C3603 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[55]), .Z(N1792)
         );
  GTECH_AND2 C3604 ( .A(N1), .B(a2stg_shr_tmp2[39]), .Z(N1793) );
  GTECH_OR2 C3605 ( .A(N1794), .B(N1795), .Z(a2stg_shr_tmp4[38]) );
  GTECH_AND2 C3606 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[54]), .Z(N1794)
         );
  GTECH_AND2 C3607 ( .A(N1), .B(a2stg_shr_tmp2[38]), .Z(N1795) );
  GTECH_OR2 C3608 ( .A(N1796), .B(N1797), .Z(a2stg_shr_tmp4[37]) );
  GTECH_AND2 C3609 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[53]), .Z(N1796)
         );
  GTECH_AND2 C3610 ( .A(N1), .B(a2stg_shr_tmp2[37]), .Z(N1797) );
  GTECH_OR2 C3611 ( .A(N1798), .B(N1799), .Z(a2stg_shr_tmp4[36]) );
  GTECH_AND2 C3612 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[52]), .Z(N1798)
         );
  GTECH_AND2 C3613 ( .A(N1), .B(a2stg_shr_tmp2[36]), .Z(N1799) );
  GTECH_OR2 C3614 ( .A(N1800), .B(N1801), .Z(a2stg_shr_tmp4[35]) );
  GTECH_AND2 C3615 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[51]), .Z(N1800)
         );
  GTECH_AND2 C3616 ( .A(N1), .B(a2stg_shr_tmp2[35]), .Z(N1801) );
  GTECH_OR2 C3617 ( .A(N1802), .B(N1803), .Z(a2stg_shr_tmp4[34]) );
  GTECH_AND2 C3618 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[50]), .Z(N1802)
         );
  GTECH_AND2 C3619 ( .A(N1), .B(a2stg_shr_tmp2[34]), .Z(N1803) );
  GTECH_OR2 C3620 ( .A(N1804), .B(N1805), .Z(a2stg_shr_tmp4[33]) );
  GTECH_AND2 C3621 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[49]), .Z(N1804)
         );
  GTECH_AND2 C3622 ( .A(N1), .B(a2stg_shr_tmp2[33]), .Z(N1805) );
  GTECH_OR2 C3623 ( .A(N1806), .B(N1807), .Z(a2stg_shr_tmp4[32]) );
  GTECH_AND2 C3624 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[48]), .Z(N1806)
         );
  GTECH_AND2 C3625 ( .A(N1), .B(a2stg_shr_tmp2[32]), .Z(N1807) );
  GTECH_OR2 C3626 ( .A(N1808), .B(N1809), .Z(a2stg_shr_tmp4[31]) );
  GTECH_AND2 C3627 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[47]), .Z(N1808)
         );
  GTECH_AND2 C3628 ( .A(N1), .B(a2stg_shr_tmp2[31]), .Z(N1809) );
  GTECH_OR2 C3629 ( .A(N1810), .B(N1811), .Z(a2stg_shr_tmp4[30]) );
  GTECH_AND2 C3630 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[46]), .Z(N1810)
         );
  GTECH_AND2 C3631 ( .A(N1), .B(a2stg_shr_tmp2[30]), .Z(N1811) );
  GTECH_OR2 C3632 ( .A(N1812), .B(N1813), .Z(a2stg_shr_tmp4[29]) );
  GTECH_AND2 C3633 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[45]), .Z(N1812)
         );
  GTECH_AND2 C3634 ( .A(N1), .B(a2stg_shr_tmp2[29]), .Z(N1813) );
  GTECH_OR2 C3635 ( .A(N1814), .B(N1815), .Z(a2stg_shr_tmp4[28]) );
  GTECH_AND2 C3636 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[44]), .Z(N1814)
         );
  GTECH_AND2 C3637 ( .A(N1), .B(a2stg_shr_tmp2[28]), .Z(N1815) );
  GTECH_OR2 C3638 ( .A(N1816), .B(N1817), .Z(a2stg_shr_tmp4[27]) );
  GTECH_AND2 C3639 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[43]), .Z(N1816)
         );
  GTECH_AND2 C3640 ( .A(N1), .B(a2stg_shr_tmp2[27]), .Z(N1817) );
  GTECH_OR2 C3641 ( .A(N1818), .B(N1819), .Z(a2stg_shr_tmp4[26]) );
  GTECH_AND2 C3642 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[42]), .Z(N1818)
         );
  GTECH_AND2 C3643 ( .A(N1), .B(a2stg_shr_tmp2[26]), .Z(N1819) );
  GTECH_OR2 C3644 ( .A(N1820), .B(N1821), .Z(a2stg_shr_tmp4[25]) );
  GTECH_AND2 C3645 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[41]), .Z(N1820)
         );
  GTECH_AND2 C3646 ( .A(N1), .B(a2stg_shr_tmp2[25]), .Z(N1821) );
  GTECH_OR2 C3647 ( .A(N1822), .B(N1823), .Z(a2stg_shr_tmp4[24]) );
  GTECH_AND2 C3648 ( .A(a2stg_shr_cnt_4[1]), .B(a2stg_shr_tmp2[40]), .Z(N1822)
         );
  GTECH_AND2 C3649 ( .A(N1), .B(a2stg_shr_tmp2[24]), .Z(N1823) );
  GTECH_OR2 C3650 ( .A(N1824), .B(N1825), .Z(a2stg_shr_tmp4[23]) );
  GTECH_AND2 C3651 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[39]), .Z(N1824)
         );
  GTECH_AND2 C3652 ( .A(N1), .B(a2stg_shr_tmp2[23]), .Z(N1825) );
  GTECH_OR2 C3653 ( .A(N1826), .B(N1827), .Z(a2stg_shr_tmp4[22]) );
  GTECH_AND2 C3654 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[38]), .Z(N1826)
         );
  GTECH_AND2 C3655 ( .A(N1), .B(a2stg_shr_tmp2[22]), .Z(N1827) );
  GTECH_OR2 C3656 ( .A(N1828), .B(N1829), .Z(a2stg_shr_tmp4[21]) );
  GTECH_AND2 C3657 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[37]), .Z(N1828)
         );
  GTECH_AND2 C3658 ( .A(N1), .B(a2stg_shr_tmp2[21]), .Z(N1829) );
  GTECH_OR2 C3659 ( .A(N1830), .B(N1831), .Z(a2stg_shr_tmp4[20]) );
  GTECH_AND2 C3660 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[36]), .Z(N1830)
         );
  GTECH_AND2 C3661 ( .A(N1), .B(a2stg_shr_tmp2[20]), .Z(N1831) );
  GTECH_OR2 C3662 ( .A(N1832), .B(N1833), .Z(a2stg_shr_tmp4[19]) );
  GTECH_AND2 C3663 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[35]), .Z(N1832)
         );
  GTECH_AND2 C3664 ( .A(N1), .B(a2stg_shr_tmp2[19]), .Z(N1833) );
  GTECH_OR2 C3665 ( .A(N1834), .B(N1835), .Z(a2stg_shr_tmp4[18]) );
  GTECH_AND2 C3666 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[34]), .Z(N1834)
         );
  GTECH_AND2 C3667 ( .A(N1), .B(a2stg_shr_tmp2[18]), .Z(N1835) );
  GTECH_OR2 C3668 ( .A(N1836), .B(N1837), .Z(a2stg_shr_tmp4[17]) );
  GTECH_AND2 C3669 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[33]), .Z(N1836)
         );
  GTECH_AND2 C3670 ( .A(N1), .B(a2stg_shr_tmp2[17]), .Z(N1837) );
  GTECH_OR2 C3671 ( .A(N1838), .B(N1839), .Z(a2stg_shr_tmp4[16]) );
  GTECH_AND2 C3672 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[32]), .Z(N1838)
         );
  GTECH_AND2 C3673 ( .A(N1), .B(a2stg_shr_tmp2[16]), .Z(N1839) );
  GTECH_OR2 C3674 ( .A(N1840), .B(N1841), .Z(a2stg_shr_tmp4[15]) );
  GTECH_AND2 C3675 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[31]), .Z(N1840)
         );
  GTECH_AND2 C3676 ( .A(N1), .B(a2stg_shr_tmp2[15]), .Z(N1841) );
  GTECH_OR2 C3677 ( .A(N1842), .B(N1843), .Z(a2stg_shr_tmp4[14]) );
  GTECH_AND2 C3678 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[30]), .Z(N1842)
         );
  GTECH_AND2 C3679 ( .A(N1), .B(a2stg_shr_tmp2[14]), .Z(N1843) );
  GTECH_OR2 C3680 ( .A(N1844), .B(N1845), .Z(a2stg_shr_tmp4[13]) );
  GTECH_AND2 C3681 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[29]), .Z(N1844)
         );
  GTECH_AND2 C3682 ( .A(N1), .B(a2stg_shr_tmp2[13]), .Z(N1845) );
  GTECH_OR2 C3683 ( .A(N1846), .B(N1847), .Z(a2stg_shr_tmp4[12]) );
  GTECH_AND2 C3684 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[28]), .Z(N1846)
         );
  GTECH_AND2 C3685 ( .A(N1), .B(a2stg_shr_tmp2[12]), .Z(N1847) );
  GTECH_OR2 C3686 ( .A(N1848), .B(N1849), .Z(a2stg_shr_tmp4[11]) );
  GTECH_AND2 C3687 ( .A(a2stg_shr_cnt_4[2]), .B(a2stg_shr_tmp2[27]), .Z(N1848)
         );
  GTECH_AND2 C3688 ( .A(N1), .B(a2stg_shr_tmp2[11]), .Z(N1849) );
  GTECH_OR2 C3689 ( .A(N1850), .B(N1851), .Z(a2stg_shr_tmp4[10]) );
  GTECH_AND2 C3690 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[26]), .Z(N1850)
         );
  GTECH_AND2 C3691 ( .A(N1), .B(a2stg_shr_tmp2[10]), .Z(N1851) );
  GTECH_OR2 C3692 ( .A(N1852), .B(N1853), .Z(a2stg_shr_tmp4[9]) );
  GTECH_AND2 C3693 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[25]), .Z(N1852)
         );
  GTECH_AND2 C3694 ( .A(N1), .B(a2stg_shr_tmp2[9]), .Z(N1853) );
  GTECH_OR2 C3695 ( .A(N1854), .B(N1855), .Z(a2stg_shr_tmp4[8]) );
  GTECH_AND2 C3696 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[24]), .Z(N1854)
         );
  GTECH_AND2 C3697 ( .A(N1), .B(a2stg_shr_tmp2[8]), .Z(N1855) );
  GTECH_OR2 C3698 ( .A(N1856), .B(N1857), .Z(a2stg_shr_tmp4[7]) );
  GTECH_AND2 C3699 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[23]), .Z(N1856)
         );
  GTECH_AND2 C3700 ( .A(N1), .B(a2stg_shr_tmp2[7]), .Z(N1857) );
  GTECH_OR2 C3701 ( .A(N1858), .B(N1859), .Z(a2stg_shr_tmp4[6]) );
  GTECH_AND2 C3702 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[22]), .Z(N1858)
         );
  GTECH_AND2 C3703 ( .A(N1), .B(a2stg_shr_tmp2[6]), .Z(N1859) );
  GTECH_OR2 C3704 ( .A(N1860), .B(N1861), .Z(a2stg_shr_tmp4[5]) );
  GTECH_AND2 C3705 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[21]), .Z(N1860)
         );
  GTECH_AND2 C3706 ( .A(N1), .B(a2stg_shr_tmp2[5]), .Z(N1861) );
  GTECH_OR2 C3707 ( .A(N1862), .B(N1863), .Z(a2stg_shr_tmp4[4]) );
  GTECH_AND2 C3708 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[20]), .Z(N1862)
         );
  GTECH_AND2 C3709 ( .A(N1), .B(a2stg_shr_tmp2[4]), .Z(N1863) );
  GTECH_OR2 C3710 ( .A(N1864), .B(N1865), .Z(a2stg_shr_tmp4[3]) );
  GTECH_AND2 C3711 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[19]), .Z(N1864)
         );
  GTECH_AND2 C3712 ( .A(N1), .B(a2stg_shr_tmp2[3]), .Z(N1865) );
  GTECH_OR2 C3713 ( .A(N1866), .B(N1867), .Z(a2stg_shr_tmp4[2]) );
  GTECH_AND2 C3714 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[18]), .Z(N1866)
         );
  GTECH_AND2 C3715 ( .A(N1), .B(a2stg_shr_tmp2[2]), .Z(N1867) );
  GTECH_OR2 C3716 ( .A(N1868), .B(N1869), .Z(a2stg_shr_tmp4[1]) );
  GTECH_AND2 C3717 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[17]), .Z(N1868)
         );
  GTECH_AND2 C3718 ( .A(N1), .B(a2stg_shr_tmp2[1]), .Z(N1869) );
  GTECH_OR2 C3719 ( .A(N1870), .B(N1871), .Z(a2stg_shr_tmp4[0]) );
  GTECH_AND2 C3720 ( .A(a2stg_shr_cnt_4[3]), .B(a2stg_shr_tmp2[16]), .Z(N1870)
         );
  GTECH_AND2 C3721 ( .A(N1), .B(a2stg_shr_tmp2[0]), .Z(N1871) );
  GTECH_NOT I_78 ( .A(N1873), .Z(a2stg_shr_tmp6[63]) );
  GTECH_AND2 C3723 ( .A(N1872), .B(a2stg_shr_tmp4[63]), .Z(N1873) );
  GTECH_NOT I_79 ( .A(a2stg_shr_cnt_3[4]), .Z(N1872) );
  GTECH_NOT I_80 ( .A(N1874), .Z(a2stg_shr_tmp6[62]) );
  GTECH_AND2 C3726 ( .A(N1872), .B(a2stg_shr_tmp4[62]), .Z(N1874) );
  GTECH_NOT I_81 ( .A(N1875), .Z(a2stg_shr_tmp6[61]) );
  GTECH_AND2 C3729 ( .A(N1872), .B(a2stg_shr_tmp4[61]), .Z(N1875) );
  GTECH_NOT I_82 ( .A(N1876), .Z(a2stg_shr_tmp6[60]) );
  GTECH_AND2 C3732 ( .A(N1872), .B(a2stg_shr_tmp4[60]), .Z(N1876) );
  GTECH_NOT I_83 ( .A(N1877), .Z(a2stg_shr_tmp6[59]) );
  GTECH_AND2 C3735 ( .A(N1872), .B(a2stg_shr_tmp4[59]), .Z(N1877) );
  GTECH_NOT I_84 ( .A(N1878), .Z(a2stg_shr_tmp6[58]) );
  GTECH_AND2 C3738 ( .A(N1872), .B(a2stg_shr_tmp4[58]), .Z(N1878) );
  GTECH_NOT I_85 ( .A(N1879), .Z(a2stg_shr_tmp6[57]) );
  GTECH_AND2 C3741 ( .A(N1872), .B(a2stg_shr_tmp4[57]), .Z(N1879) );
  GTECH_NOT I_86 ( .A(N1880), .Z(a2stg_shr_tmp6[56]) );
  GTECH_AND2 C3744 ( .A(N1872), .B(a2stg_shr_tmp4[56]), .Z(N1880) );
  GTECH_NOT I_87 ( .A(N1883), .Z(a2stg_shr_tmp6[55]) );
  GTECH_OR2 C3747 ( .A(N1881), .B(N1882), .Z(N1883) );
  GTECH_AND2 C3748 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[63]), .Z(N1881)
         );
  GTECH_AND2 C3749 ( .A(N1872), .B(a2stg_shr_tmp4[55]), .Z(N1882) );
  GTECH_NOT I_88 ( .A(N1886), .Z(a2stg_shr_tmp6[54]) );
  GTECH_OR2 C3752 ( .A(N1884), .B(N1885), .Z(N1886) );
  GTECH_AND2 C3753 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[62]), .Z(N1884)
         );
  GTECH_AND2 C3754 ( .A(N1872), .B(a2stg_shr_tmp4[54]), .Z(N1885) );
  GTECH_NOT I_89 ( .A(N1889), .Z(a2stg_shr_tmp6[53]) );
  GTECH_OR2 C3757 ( .A(N1887), .B(N1888), .Z(N1889) );
  GTECH_AND2 C3758 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[61]), .Z(N1887)
         );
  GTECH_AND2 C3759 ( .A(N1872), .B(a2stg_shr_tmp4[53]), .Z(N1888) );
  GTECH_NOT I_90 ( .A(N1892), .Z(a2stg_shr_tmp6[52]) );
  GTECH_OR2 C3762 ( .A(N1890), .B(N1891), .Z(N1892) );
  GTECH_AND2 C3763 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[60]), .Z(N1890)
         );
  GTECH_AND2 C3764 ( .A(N1872), .B(a2stg_shr_tmp4[52]), .Z(N1891) );
  GTECH_NOT I_91 ( .A(N1895), .Z(a2stg_shr_tmp6[51]) );
  GTECH_OR2 C3767 ( .A(N1893), .B(N1894), .Z(N1895) );
  GTECH_AND2 C3768 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[59]), .Z(N1893)
         );
  GTECH_AND2 C3769 ( .A(N1872), .B(a2stg_shr_tmp4[51]), .Z(N1894) );
  GTECH_NOT I_92 ( .A(N1898), .Z(a2stg_shr_tmp6[50]) );
  GTECH_OR2 C3772 ( .A(N1896), .B(N1897), .Z(N1898) );
  GTECH_AND2 C3773 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[58]), .Z(N1896)
         );
  GTECH_AND2 C3774 ( .A(N1872), .B(a2stg_shr_tmp4[50]), .Z(N1897) );
  GTECH_NOT I_93 ( .A(N1901), .Z(a2stg_shr_tmp6[49]) );
  GTECH_OR2 C3777 ( .A(N1899), .B(N1900), .Z(N1901) );
  GTECH_AND2 C3778 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[57]), .Z(N1899)
         );
  GTECH_AND2 C3779 ( .A(N1872), .B(a2stg_shr_tmp4[49]), .Z(N1900) );
  GTECH_NOT I_94 ( .A(N1904), .Z(a2stg_shr_tmp6[48]) );
  GTECH_OR2 C3782 ( .A(N1902), .B(N1903), .Z(N1904) );
  GTECH_AND2 C3783 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[56]), .Z(N1902)
         );
  GTECH_AND2 C3784 ( .A(N1872), .B(a2stg_shr_tmp4[48]), .Z(N1903) );
  GTECH_NOT I_95 ( .A(N1907), .Z(a2stg_shr_tmp6[47]) );
  GTECH_OR2 C3787 ( .A(N1905), .B(N1906), .Z(N1907) );
  GTECH_AND2 C3788 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[55]), .Z(N1905)
         );
  GTECH_AND2 C3789 ( .A(N1872), .B(a2stg_shr_tmp4[47]), .Z(N1906) );
  GTECH_NOT I_96 ( .A(N1910), .Z(a2stg_shr_tmp6[46]) );
  GTECH_OR2 C3792 ( .A(N1908), .B(N1909), .Z(N1910) );
  GTECH_AND2 C3793 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[54]), .Z(N1908)
         );
  GTECH_AND2 C3794 ( .A(N1872), .B(a2stg_shr_tmp4[46]), .Z(N1909) );
  GTECH_NOT I_97 ( .A(N1913), .Z(a2stg_shr_tmp6[45]) );
  GTECH_OR2 C3797 ( .A(N1911), .B(N1912), .Z(N1913) );
  GTECH_AND2 C3798 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[53]), .Z(N1911)
         );
  GTECH_AND2 C3799 ( .A(N1872), .B(a2stg_shr_tmp4[45]), .Z(N1912) );
  GTECH_NOT I_98 ( .A(N1916), .Z(a2stg_shr_tmp6[44]) );
  GTECH_OR2 C3802 ( .A(N1914), .B(N1915), .Z(N1916) );
  GTECH_AND2 C3803 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[52]), .Z(N1914)
         );
  GTECH_AND2 C3804 ( .A(N1872), .B(a2stg_shr_tmp4[44]), .Z(N1915) );
  GTECH_NOT I_99 ( .A(N1919), .Z(a2stg_shr_tmp6[43]) );
  GTECH_OR2 C3807 ( .A(N1917), .B(N1918), .Z(N1919) );
  GTECH_AND2 C3808 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[51]), .Z(N1917)
         );
  GTECH_AND2 C3809 ( .A(N1872), .B(a2stg_shr_tmp4[43]), .Z(N1918) );
  GTECH_NOT I_100 ( .A(N1922), .Z(a2stg_shr_tmp6[42]) );
  GTECH_OR2 C3812 ( .A(N1920), .B(N1921), .Z(N1922) );
  GTECH_AND2 C3813 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[50]), .Z(N1920)
         );
  GTECH_AND2 C3814 ( .A(N1872), .B(a2stg_shr_tmp4[42]), .Z(N1921) );
  GTECH_NOT I_101 ( .A(N1925), .Z(a2stg_shr_tmp6[41]) );
  GTECH_OR2 C3817 ( .A(N1923), .B(N1924), .Z(N1925) );
  GTECH_AND2 C3818 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[49]), .Z(N1923)
         );
  GTECH_AND2 C3819 ( .A(N1872), .B(a2stg_shr_tmp4[41]), .Z(N1924) );
  GTECH_NOT I_102 ( .A(N1928), .Z(a2stg_shr_tmp6[40]) );
  GTECH_OR2 C3822 ( .A(N1926), .B(N1927), .Z(N1928) );
  GTECH_AND2 C3823 ( .A(a2stg_shr_cnt_3[0]), .B(a2stg_shr_tmp4[48]), .Z(N1926)
         );
  GTECH_AND2 C3824 ( .A(N1872), .B(a2stg_shr_tmp4[40]), .Z(N1927) );
  GTECH_NOT I_103 ( .A(N1931), .Z(a2stg_shr_tmp6[39]) );
  GTECH_OR2 C3827 ( .A(N1929), .B(N1930), .Z(N1931) );
  GTECH_AND2 C3828 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[47]), .Z(N1929)
         );
  GTECH_AND2 C3829 ( .A(N1872), .B(a2stg_shr_tmp4[39]), .Z(N1930) );
  GTECH_NOT I_104 ( .A(N1934), .Z(a2stg_shr_tmp6[38]) );
  GTECH_OR2 C3832 ( .A(N1932), .B(N1933), .Z(N1934) );
  GTECH_AND2 C3833 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[46]), .Z(N1932)
         );
  GTECH_AND2 C3834 ( .A(N1872), .B(a2stg_shr_tmp4[38]), .Z(N1933) );
  GTECH_NOT I_105 ( .A(N1937), .Z(a2stg_shr_tmp6[37]) );
  GTECH_OR2 C3837 ( .A(N1935), .B(N1936), .Z(N1937) );
  GTECH_AND2 C3838 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[45]), .Z(N1935)
         );
  GTECH_AND2 C3839 ( .A(N1872), .B(a2stg_shr_tmp4[37]), .Z(N1936) );
  GTECH_NOT I_106 ( .A(N1940), .Z(a2stg_shr_tmp6[36]) );
  GTECH_OR2 C3842 ( .A(N1938), .B(N1939), .Z(N1940) );
  GTECH_AND2 C3843 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[44]), .Z(N1938)
         );
  GTECH_AND2 C3844 ( .A(N1872), .B(a2stg_shr_tmp4[36]), .Z(N1939) );
  GTECH_NOT I_107 ( .A(N1943), .Z(a2stg_shr_tmp6[35]) );
  GTECH_OR2 C3847 ( .A(N1941), .B(N1942), .Z(N1943) );
  GTECH_AND2 C3848 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[43]), .Z(N1941)
         );
  GTECH_AND2 C3849 ( .A(N1872), .B(a2stg_shr_tmp4[35]), .Z(N1942) );
  GTECH_NOT I_108 ( .A(N1946), .Z(a2stg_shr_tmp6[34]) );
  GTECH_OR2 C3852 ( .A(N1944), .B(N1945), .Z(N1946) );
  GTECH_AND2 C3853 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[42]), .Z(N1944)
         );
  GTECH_AND2 C3854 ( .A(N1872), .B(a2stg_shr_tmp4[34]), .Z(N1945) );
  GTECH_NOT I_109 ( .A(N1949), .Z(a2stg_shr_tmp6[33]) );
  GTECH_OR2 C3857 ( .A(N1947), .B(N1948), .Z(N1949) );
  GTECH_AND2 C3858 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[41]), .Z(N1947)
         );
  GTECH_AND2 C3859 ( .A(N1872), .B(a2stg_shr_tmp4[33]), .Z(N1948) );
  GTECH_NOT I_110 ( .A(N1952), .Z(a2stg_shr_tmp6[32]) );
  GTECH_OR2 C3862 ( .A(N1950), .B(N1951), .Z(N1952) );
  GTECH_AND2 C3863 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[40]), .Z(N1950)
         );
  GTECH_AND2 C3864 ( .A(N1872), .B(a2stg_shr_tmp4[32]), .Z(N1951) );
  GTECH_NOT I_111 ( .A(N1955), .Z(a2stg_shr_tmp6[31]) );
  GTECH_OR2 C3867 ( .A(N1953), .B(N1954), .Z(N1955) );
  GTECH_AND2 C3868 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[39]), .Z(N1953)
         );
  GTECH_AND2 C3869 ( .A(N1872), .B(a2stg_shr_tmp4[31]), .Z(N1954) );
  GTECH_NOT I_112 ( .A(N1958), .Z(a2stg_shr_tmp6[30]) );
  GTECH_OR2 C3872 ( .A(N1956), .B(N1957), .Z(N1958) );
  GTECH_AND2 C3873 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[38]), .Z(N1956)
         );
  GTECH_AND2 C3874 ( .A(N1872), .B(a2stg_shr_tmp4[30]), .Z(N1957) );
  GTECH_NOT I_113 ( .A(N1961), .Z(a2stg_shr_tmp6[29]) );
  GTECH_OR2 C3877 ( .A(N1959), .B(N1960), .Z(N1961) );
  GTECH_AND2 C3878 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[37]), .Z(N1959)
         );
  GTECH_AND2 C3879 ( .A(N1872), .B(a2stg_shr_tmp4[29]), .Z(N1960) );
  GTECH_NOT I_114 ( .A(N1964), .Z(a2stg_shr_tmp6[28]) );
  GTECH_OR2 C3882 ( .A(N1962), .B(N1963), .Z(N1964) );
  GTECH_AND2 C3883 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[36]), .Z(N1962)
         );
  GTECH_AND2 C3884 ( .A(N1872), .B(a2stg_shr_tmp4[28]), .Z(N1963) );
  GTECH_NOT I_115 ( .A(N1967), .Z(a2stg_shr_tmp6[27]) );
  GTECH_OR2 C3887 ( .A(N1965), .B(N1966), .Z(N1967) );
  GTECH_AND2 C3888 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[35]), .Z(N1965)
         );
  GTECH_AND2 C3889 ( .A(N1872), .B(a2stg_shr_tmp4[27]), .Z(N1966) );
  GTECH_NOT I_116 ( .A(N1970), .Z(a2stg_shr_tmp6[26]) );
  GTECH_OR2 C3892 ( .A(N1968), .B(N1969), .Z(N1970) );
  GTECH_AND2 C3893 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[34]), .Z(N1968)
         );
  GTECH_AND2 C3894 ( .A(N1872), .B(a2stg_shr_tmp4[26]), .Z(N1969) );
  GTECH_NOT I_117 ( .A(N1973), .Z(a2stg_shr_tmp6[25]) );
  GTECH_OR2 C3897 ( .A(N1971), .B(N1972), .Z(N1973) );
  GTECH_AND2 C3898 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[33]), .Z(N1971)
         );
  GTECH_AND2 C3899 ( .A(N1872), .B(a2stg_shr_tmp4[25]), .Z(N1972) );
  GTECH_NOT I_118 ( .A(N1976), .Z(a2stg_shr_tmp6[24]) );
  GTECH_OR2 C3902 ( .A(N1974), .B(N1975), .Z(N1976) );
  GTECH_AND2 C3903 ( .A(a2stg_shr_cnt_3[1]), .B(a2stg_shr_tmp4[32]), .Z(N1974)
         );
  GTECH_AND2 C3904 ( .A(N1872), .B(a2stg_shr_tmp4[24]), .Z(N1975) );
  GTECH_NOT I_119 ( .A(N1979), .Z(a2stg_shr_tmp6[23]) );
  GTECH_OR2 C3907 ( .A(N1977), .B(N1978), .Z(N1979) );
  GTECH_AND2 C3908 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[31]), .Z(N1977)
         );
  GTECH_AND2 C3909 ( .A(N1872), .B(a2stg_shr_tmp4[23]), .Z(N1978) );
  GTECH_NOT I_120 ( .A(N1982), .Z(a2stg_shr_tmp6[22]) );
  GTECH_OR2 C3912 ( .A(N1980), .B(N1981), .Z(N1982) );
  GTECH_AND2 C3913 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[30]), .Z(N1980)
         );
  GTECH_AND2 C3914 ( .A(N1872), .B(a2stg_shr_tmp4[22]), .Z(N1981) );
  GTECH_NOT I_121 ( .A(N1985), .Z(a2stg_shr_tmp6[21]) );
  GTECH_OR2 C3917 ( .A(N1983), .B(N1984), .Z(N1985) );
  GTECH_AND2 C3918 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[29]), .Z(N1983)
         );
  GTECH_AND2 C3919 ( .A(N1872), .B(a2stg_shr_tmp4[21]), .Z(N1984) );
  GTECH_NOT I_122 ( .A(N1988), .Z(a2stg_shr_tmp6[20]) );
  GTECH_OR2 C3922 ( .A(N1986), .B(N1987), .Z(N1988) );
  GTECH_AND2 C3923 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[28]), .Z(N1986)
         );
  GTECH_AND2 C3924 ( .A(N1872), .B(a2stg_shr_tmp4[20]), .Z(N1987) );
  GTECH_NOT I_123 ( .A(N1991), .Z(a2stg_shr_tmp6[19]) );
  GTECH_OR2 C3927 ( .A(N1989), .B(N1990), .Z(N1991) );
  GTECH_AND2 C3928 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[27]), .Z(N1989)
         );
  GTECH_AND2 C3929 ( .A(N1872), .B(a2stg_shr_tmp4[19]), .Z(N1990) );
  GTECH_NOT I_124 ( .A(N1994), .Z(a2stg_shr_tmp6[18]) );
  GTECH_OR2 C3932 ( .A(N1992), .B(N1993), .Z(N1994) );
  GTECH_AND2 C3933 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[26]), .Z(N1992)
         );
  GTECH_AND2 C3934 ( .A(N1872), .B(a2stg_shr_tmp4[18]), .Z(N1993) );
  GTECH_NOT I_125 ( .A(N1997), .Z(a2stg_shr_tmp6[17]) );
  GTECH_OR2 C3937 ( .A(N1995), .B(N1996), .Z(N1997) );
  GTECH_AND2 C3938 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[25]), .Z(N1995)
         );
  GTECH_AND2 C3939 ( .A(N1872), .B(a2stg_shr_tmp4[17]), .Z(N1996) );
  GTECH_NOT I_126 ( .A(N2000), .Z(a2stg_shr_tmp6[16]) );
  GTECH_OR2 C3942 ( .A(N1998), .B(N1999), .Z(N2000) );
  GTECH_AND2 C3943 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[24]), .Z(N1998)
         );
  GTECH_AND2 C3944 ( .A(N1872), .B(a2stg_shr_tmp4[16]), .Z(N1999) );
  GTECH_NOT I_127 ( .A(N2003), .Z(a2stg_shr_tmp6[15]) );
  GTECH_OR2 C3947 ( .A(N2001), .B(N2002), .Z(N2003) );
  GTECH_AND2 C3948 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[23]), .Z(N2001)
         );
  GTECH_AND2 C3949 ( .A(N1872), .B(a2stg_shr_tmp4[15]), .Z(N2002) );
  GTECH_NOT I_128 ( .A(N2006), .Z(a2stg_shr_tmp6[14]) );
  GTECH_OR2 C3952 ( .A(N2004), .B(N2005), .Z(N2006) );
  GTECH_AND2 C3953 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[22]), .Z(N2004)
         );
  GTECH_AND2 C3954 ( .A(N1872), .B(a2stg_shr_tmp4[14]), .Z(N2005) );
  GTECH_NOT I_129 ( .A(N2009), .Z(a2stg_shr_tmp6[13]) );
  GTECH_OR2 C3957 ( .A(N2007), .B(N2008), .Z(N2009) );
  GTECH_AND2 C3958 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[21]), .Z(N2007)
         );
  GTECH_AND2 C3959 ( .A(N1872), .B(a2stg_shr_tmp4[13]), .Z(N2008) );
  GTECH_NOT I_130 ( .A(N2012), .Z(a2stg_shr_tmp6[12]) );
  GTECH_OR2 C3962 ( .A(N2010), .B(N2011), .Z(N2012) );
  GTECH_AND2 C3963 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[20]), .Z(N2010)
         );
  GTECH_AND2 C3964 ( .A(N1872), .B(a2stg_shr_tmp4[12]), .Z(N2011) );
  GTECH_NOT I_131 ( .A(N2015), .Z(a2stg_shr_tmp6[11]) );
  GTECH_OR2 C3967 ( .A(N2013), .B(N2014), .Z(N2015) );
  GTECH_AND2 C3968 ( .A(a2stg_shr_cnt_3[2]), .B(a2stg_shr_tmp4[19]), .Z(N2013)
         );
  GTECH_AND2 C3969 ( .A(N1872), .B(a2stg_shr_tmp4[11]), .Z(N2014) );
  GTECH_NOT I_132 ( .A(N2018), .Z(a2stg_shr_tmp6[10]) );
  GTECH_OR2 C3972 ( .A(N2016), .B(N2017), .Z(N2018) );
  GTECH_AND2 C3973 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[18]), .Z(N2016)
         );
  GTECH_AND2 C3974 ( .A(N1872), .B(a2stg_shr_tmp4[10]), .Z(N2017) );
  GTECH_NOT I_133 ( .A(N2021), .Z(a2stg_shr_tmp6[9]) );
  GTECH_OR2 C3977 ( .A(N2019), .B(N2020), .Z(N2021) );
  GTECH_AND2 C3978 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[17]), .Z(N2019)
         );
  GTECH_AND2 C3979 ( .A(N1872), .B(a2stg_shr_tmp4[9]), .Z(N2020) );
  GTECH_NOT I_134 ( .A(N2024), .Z(a2stg_shr_tmp6[8]) );
  GTECH_OR2 C3982 ( .A(N2022), .B(N2023), .Z(N2024) );
  GTECH_AND2 C3983 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[16]), .Z(N2022)
         );
  GTECH_AND2 C3984 ( .A(N1872), .B(a2stg_shr_tmp4[8]), .Z(N2023) );
  GTECH_NOT I_135 ( .A(N2027), .Z(a2stg_shr_tmp6[7]) );
  GTECH_OR2 C3987 ( .A(N2025), .B(N2026), .Z(N2027) );
  GTECH_AND2 C3988 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[15]), .Z(N2025)
         );
  GTECH_AND2 C3989 ( .A(N1872), .B(a2stg_shr_tmp4[7]), .Z(N2026) );
  GTECH_NOT I_136 ( .A(N2030), .Z(a2stg_shr_tmp6[6]) );
  GTECH_OR2 C3992 ( .A(N2028), .B(N2029), .Z(N2030) );
  GTECH_AND2 C3993 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[14]), .Z(N2028)
         );
  GTECH_AND2 C3994 ( .A(N1872), .B(a2stg_shr_tmp4[6]), .Z(N2029) );
  GTECH_NOT I_137 ( .A(N2033), .Z(a2stg_shr_tmp6[5]) );
  GTECH_OR2 C3997 ( .A(N2031), .B(N2032), .Z(N2033) );
  GTECH_AND2 C3998 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[13]), .Z(N2031)
         );
  GTECH_AND2 C3999 ( .A(N1872), .B(a2stg_shr_tmp4[5]), .Z(N2032) );
  GTECH_NOT I_138 ( .A(N2036), .Z(a2stg_shr_tmp6[4]) );
  GTECH_OR2 C4002 ( .A(N2034), .B(N2035), .Z(N2036) );
  GTECH_AND2 C4003 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[12]), .Z(N2034)
         );
  GTECH_AND2 C4004 ( .A(N1872), .B(a2stg_shr_tmp4[4]), .Z(N2035) );
  GTECH_NOT I_139 ( .A(N2039), .Z(a2stg_shr_tmp6[3]) );
  GTECH_OR2 C4007 ( .A(N2037), .B(N2038), .Z(N2039) );
  GTECH_AND2 C4008 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[11]), .Z(N2037)
         );
  GTECH_AND2 C4009 ( .A(N1872), .B(a2stg_shr_tmp4[3]), .Z(N2038) );
  GTECH_NOT I_140 ( .A(N2042), .Z(a2stg_shr_tmp6[2]) );
  GTECH_OR2 C4012 ( .A(N2040), .B(N2041), .Z(N2042) );
  GTECH_AND2 C4013 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[10]), .Z(N2040)
         );
  GTECH_AND2 C4014 ( .A(N1872), .B(a2stg_shr_tmp4[2]), .Z(N2041) );
  GTECH_NOT I_141 ( .A(N2045), .Z(a2stg_shr_tmp6[1]) );
  GTECH_OR2 C4017 ( .A(N2043), .B(N2044), .Z(N2045) );
  GTECH_AND2 C4018 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[9]), .Z(N2043)
         );
  GTECH_AND2 C4019 ( .A(N1872), .B(a2stg_shr_tmp4[1]), .Z(N2044) );
  GTECH_NOT I_142 ( .A(N2048), .Z(a2stg_shr_tmp6[0]) );
  GTECH_OR2 C4022 ( .A(N2046), .B(N2047), .Z(N2048) );
  GTECH_AND2 C4023 ( .A(a2stg_shr_cnt_3[3]), .B(a2stg_shr_tmp4[8]), .Z(N2046)
         );
  GTECH_AND2 C4024 ( .A(N1872), .B(a2stg_shr_tmp4[0]), .Z(N2047) );
  GTECH_NOT I_143 ( .A(N2049), .Z(a2stg_shr_tmp8[63]) );
  GTECH_OR2 C4027 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[63]), .Z(N2049)
         );
  GTECH_NOT I_144 ( .A(N2050), .Z(a2stg_shr_tmp8[62]) );
  GTECH_OR2 C4029 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[62]), .Z(N2050)
         );
  GTECH_NOT I_145 ( .A(N2051), .Z(a2stg_shr_tmp8[61]) );
  GTECH_OR2 C4031 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[61]), .Z(N2051)
         );
  GTECH_NOT I_146 ( .A(N2052), .Z(a2stg_shr_tmp8[60]) );
  GTECH_OR2 C4033 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[60]), .Z(N2052)
         );
  GTECH_NOT I_147 ( .A(N2056), .Z(a2stg_shr_tmp8[59]) );
  GTECH_AND2 C4035 ( .A(N2053), .B(N2055), .Z(N2056) );
  GTECH_OR2 C4036 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[59]), .Z(N2053)
         );
  GTECH_OR2 C4037 ( .A(N2054), .B(a2stg_shr_tmp6[63]), .Z(N2055) );
  GTECH_NOT I_148 ( .A(a2stg_shr_cnt_2[1]), .Z(N2054) );
  GTECH_NOT I_149 ( .A(N2059), .Z(a2stg_shr_tmp8[58]) );
  GTECH_AND2 C4040 ( .A(N2057), .B(N2058), .Z(N2059) );
  GTECH_OR2 C4041 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[58]), .Z(N2057)
         );
  GTECH_OR2 C4042 ( .A(N2054), .B(a2stg_shr_tmp6[62]), .Z(N2058) );
  GTECH_NOT I_150 ( .A(N2062), .Z(a2stg_shr_tmp8[57]) );
  GTECH_AND2 C4045 ( .A(N2060), .B(N2061), .Z(N2062) );
  GTECH_OR2 C4046 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[57]), .Z(N2060)
         );
  GTECH_OR2 C4047 ( .A(N2054), .B(a2stg_shr_tmp6[61]), .Z(N2061) );
  GTECH_NOT I_151 ( .A(N2065), .Z(a2stg_shr_tmp8[56]) );
  GTECH_AND2 C4050 ( .A(N2063), .B(N2064), .Z(N2065) );
  GTECH_OR2 C4051 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[56]), .Z(N2063)
         );
  GTECH_OR2 C4052 ( .A(N2054), .B(a2stg_shr_tmp6[60]), .Z(N2064) );
  GTECH_NOT I_152 ( .A(N2068), .Z(a2stg_shr_tmp8[55]) );
  GTECH_AND2 C4055 ( .A(N2066), .B(N2067), .Z(N2068) );
  GTECH_OR2 C4056 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[55]), .Z(N2066)
         );
  GTECH_OR2 C4057 ( .A(N2054), .B(a2stg_shr_tmp6[59]), .Z(N2067) );
  GTECH_NOT I_153 ( .A(N2071), .Z(a2stg_shr_tmp8[54]) );
  GTECH_AND2 C4060 ( .A(N2069), .B(N2070), .Z(N2071) );
  GTECH_OR2 C4061 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[54]), .Z(N2069)
         );
  GTECH_OR2 C4062 ( .A(N2054), .B(a2stg_shr_tmp6[58]), .Z(N2070) );
  GTECH_NOT I_154 ( .A(N2074), .Z(a2stg_shr_tmp8[53]) );
  GTECH_AND2 C4065 ( .A(N2072), .B(N2073), .Z(N2074) );
  GTECH_OR2 C4066 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[53]), .Z(N2072)
         );
  GTECH_OR2 C4067 ( .A(N2054), .B(a2stg_shr_tmp6[57]), .Z(N2073) );
  GTECH_NOT I_155 ( .A(N2077), .Z(a2stg_shr_tmp8[52]) );
  GTECH_AND2 C4070 ( .A(N2075), .B(N2076), .Z(N2077) );
  GTECH_OR2 C4071 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[52]), .Z(N2075)
         );
  GTECH_OR2 C4072 ( .A(N2054), .B(a2stg_shr_tmp6[56]), .Z(N2076) );
  GTECH_NOT I_156 ( .A(N2080), .Z(a2stg_shr_tmp8[51]) );
  GTECH_AND2 C4075 ( .A(N2078), .B(N2079), .Z(N2080) );
  GTECH_OR2 C4076 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[51]), .Z(N2078)
         );
  GTECH_OR2 C4077 ( .A(N2054), .B(a2stg_shr_tmp6[55]), .Z(N2079) );
  GTECH_NOT I_157 ( .A(N2083), .Z(a2stg_shr_tmp8[50]) );
  GTECH_AND2 C4080 ( .A(N2081), .B(N2082), .Z(N2083) );
  GTECH_OR2 C4081 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[50]), .Z(N2081)
         );
  GTECH_OR2 C4082 ( .A(N2054), .B(a2stg_shr_tmp6[54]), .Z(N2082) );
  GTECH_NOT I_158 ( .A(N2086), .Z(a2stg_shr_tmp8[49]) );
  GTECH_AND2 C4085 ( .A(N2084), .B(N2085), .Z(N2086) );
  GTECH_OR2 C4086 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[49]), .Z(N2084)
         );
  GTECH_OR2 C4087 ( .A(N2054), .B(a2stg_shr_tmp6[53]), .Z(N2085) );
  GTECH_NOT I_159 ( .A(N2089), .Z(a2stg_shr_tmp8[48]) );
  GTECH_AND2 C4090 ( .A(N2087), .B(N2088), .Z(N2089) );
  GTECH_OR2 C4091 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[48]), .Z(N2087)
         );
  GTECH_OR2 C4092 ( .A(N2054), .B(a2stg_shr_tmp6[52]), .Z(N2088) );
  GTECH_NOT I_160 ( .A(N2092), .Z(a2stg_shr_tmp8[47]) );
  GTECH_AND2 C4095 ( .A(N2090), .B(N2091), .Z(N2092) );
  GTECH_OR2 C4096 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[47]), .Z(N2090)
         );
  GTECH_OR2 C4097 ( .A(N2054), .B(a2stg_shr_tmp6[51]), .Z(N2091) );
  GTECH_NOT I_161 ( .A(N2095), .Z(a2stg_shr_tmp8[46]) );
  GTECH_AND2 C4100 ( .A(N2093), .B(N2094), .Z(N2095) );
  GTECH_OR2 C4101 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[46]), .Z(N2093)
         );
  GTECH_OR2 C4102 ( .A(N2054), .B(a2stg_shr_tmp6[50]), .Z(N2094) );
  GTECH_NOT I_162 ( .A(N2098), .Z(a2stg_shr_tmp8[45]) );
  GTECH_AND2 C4105 ( .A(N2096), .B(N2097), .Z(N2098) );
  GTECH_OR2 C4106 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[45]), .Z(N2096)
         );
  GTECH_OR2 C4107 ( .A(N2054), .B(a2stg_shr_tmp6[49]), .Z(N2097) );
  GTECH_NOT I_163 ( .A(N2101), .Z(a2stg_shr_tmp8[44]) );
  GTECH_AND2 C4110 ( .A(N2099), .B(N2100), .Z(N2101) );
  GTECH_OR2 C4111 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[44]), .Z(N2099)
         );
  GTECH_OR2 C4112 ( .A(N2054), .B(a2stg_shr_tmp6[48]), .Z(N2100) );
  GTECH_NOT I_164 ( .A(N2104), .Z(a2stg_shr_tmp8[43]) );
  GTECH_AND2 C4115 ( .A(N2102), .B(N2103), .Z(N2104) );
  GTECH_OR2 C4116 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[43]), .Z(N2102)
         );
  GTECH_OR2 C4117 ( .A(N2054), .B(a2stg_shr_tmp6[47]), .Z(N2103) );
  GTECH_NOT I_165 ( .A(N2107), .Z(a2stg_shr_tmp8[42]) );
  GTECH_AND2 C4120 ( .A(N2105), .B(N2106), .Z(N2107) );
  GTECH_OR2 C4121 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[42]), .Z(N2105)
         );
  GTECH_OR2 C4122 ( .A(N2054), .B(a2stg_shr_tmp6[46]), .Z(N2106) );
  GTECH_NOT I_166 ( .A(N2110), .Z(a2stg_shr_tmp8[41]) );
  GTECH_AND2 C4125 ( .A(N2108), .B(N2109), .Z(N2110) );
  GTECH_OR2 C4126 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[41]), .Z(N2108)
         );
  GTECH_OR2 C4127 ( .A(N2054), .B(a2stg_shr_tmp6[45]), .Z(N2109) );
  GTECH_NOT I_167 ( .A(N2113), .Z(a2stg_shr_tmp8[40]) );
  GTECH_AND2 C4130 ( .A(N2111), .B(N2112), .Z(N2113) );
  GTECH_OR2 C4131 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[40]), .Z(N2111)
         );
  GTECH_OR2 C4132 ( .A(N2054), .B(a2stg_shr_tmp6[44]), .Z(N2112) );
  GTECH_NOT I_168 ( .A(N2116), .Z(a2stg_shr_tmp8[39]) );
  GTECH_AND2 C4135 ( .A(N2114), .B(N2115), .Z(N2116) );
  GTECH_OR2 C4136 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[39]), .Z(N2114)
         );
  GTECH_OR2 C4137 ( .A(N2054), .B(a2stg_shr_tmp6[43]), .Z(N2115) );
  GTECH_NOT I_169 ( .A(N2119), .Z(a2stg_shr_tmp8[38]) );
  GTECH_AND2 C4140 ( .A(N2117), .B(N2118), .Z(N2119) );
  GTECH_OR2 C4141 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[38]), .Z(N2117)
         );
  GTECH_OR2 C4142 ( .A(N2054), .B(a2stg_shr_tmp6[42]), .Z(N2118) );
  GTECH_NOT I_170 ( .A(N2122), .Z(a2stg_shr_tmp8[37]) );
  GTECH_AND2 C4145 ( .A(N2120), .B(N2121), .Z(N2122) );
  GTECH_OR2 C4146 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[37]), .Z(N2120)
         );
  GTECH_OR2 C4147 ( .A(N2054), .B(a2stg_shr_tmp6[41]), .Z(N2121) );
  GTECH_NOT I_171 ( .A(N2125), .Z(a2stg_shr_tmp8[36]) );
  GTECH_AND2 C4150 ( .A(N2123), .B(N2124), .Z(N2125) );
  GTECH_OR2 C4151 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[36]), .Z(N2123)
         );
  GTECH_OR2 C4152 ( .A(N2054), .B(a2stg_shr_tmp6[40]), .Z(N2124) );
  GTECH_NOT I_172 ( .A(N2128), .Z(a2stg_shr_tmp8[35]) );
  GTECH_AND2 C4155 ( .A(N2126), .B(N2127), .Z(N2128) );
  GTECH_OR2 C4156 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[35]), .Z(N2126)
         );
  GTECH_OR2 C4157 ( .A(N2054), .B(a2stg_shr_tmp6[39]), .Z(N2127) );
  GTECH_NOT I_173 ( .A(N2131), .Z(a2stg_shr_tmp8[34]) );
  GTECH_AND2 C4160 ( .A(N2129), .B(N2130), .Z(N2131) );
  GTECH_OR2 C4161 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[34]), .Z(N2129)
         );
  GTECH_OR2 C4162 ( .A(N2054), .B(a2stg_shr_tmp6[38]), .Z(N2130) );
  GTECH_NOT I_174 ( .A(N2134), .Z(a2stg_shr_tmp8[33]) );
  GTECH_AND2 C4165 ( .A(N2132), .B(N2133), .Z(N2134) );
  GTECH_OR2 C4166 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[33]), .Z(N2132)
         );
  GTECH_OR2 C4167 ( .A(N2054), .B(a2stg_shr_tmp6[37]), .Z(N2133) );
  GTECH_NOT I_175 ( .A(N2137), .Z(a2stg_shr_tmp8[32]) );
  GTECH_AND2 C4170 ( .A(N2135), .B(N2136), .Z(N2137) );
  GTECH_OR2 C4171 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[32]), .Z(N2135)
         );
  GTECH_OR2 C4172 ( .A(N2054), .B(a2stg_shr_tmp6[36]), .Z(N2136) );
  GTECH_NOT I_176 ( .A(N2140), .Z(a2stg_shr_tmp8[31]) );
  GTECH_AND2 C4175 ( .A(N2138), .B(N2139), .Z(N2140) );
  GTECH_OR2 C4176 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[31]), .Z(N2138)
         );
  GTECH_OR2 C4177 ( .A(N2054), .B(a2stg_shr_tmp6[35]), .Z(N2139) );
  GTECH_NOT I_177 ( .A(N2143), .Z(a2stg_shr_tmp8[30]) );
  GTECH_AND2 C4180 ( .A(N2141), .B(N2142), .Z(N2143) );
  GTECH_OR2 C4181 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[30]), .Z(N2141)
         );
  GTECH_OR2 C4182 ( .A(N2054), .B(a2stg_shr_tmp6[34]), .Z(N2142) );
  GTECH_NOT I_178 ( .A(N2146), .Z(a2stg_shr_tmp8[29]) );
  GTECH_AND2 C4185 ( .A(N2144), .B(N2145), .Z(N2146) );
  GTECH_OR2 C4186 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[29]), .Z(N2144)
         );
  GTECH_OR2 C4187 ( .A(N2054), .B(a2stg_shr_tmp6[33]), .Z(N2145) );
  GTECH_NOT I_179 ( .A(N2149), .Z(a2stg_shr_tmp8[28]) );
  GTECH_AND2 C4190 ( .A(N2147), .B(N2148), .Z(N2149) );
  GTECH_OR2 C4191 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[28]), .Z(N2147)
         );
  GTECH_OR2 C4192 ( .A(N2054), .B(a2stg_shr_tmp6[32]), .Z(N2148) );
  GTECH_NOT I_180 ( .A(N2152), .Z(a2stg_shr_tmp8[27]) );
  GTECH_AND2 C4195 ( .A(N2150), .B(N2151), .Z(N2152) );
  GTECH_OR2 C4196 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[27]), .Z(N2150)
         );
  GTECH_OR2 C4197 ( .A(N2054), .B(a2stg_shr_tmp6[31]), .Z(N2151) );
  GTECH_NOT I_181 ( .A(N2155), .Z(a2stg_shr_tmp8[26]) );
  GTECH_AND2 C4200 ( .A(N2153), .B(N2154), .Z(N2155) );
  GTECH_OR2 C4201 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[26]), .Z(N2153)
         );
  GTECH_OR2 C4202 ( .A(N2054), .B(a2stg_shr_tmp6[30]), .Z(N2154) );
  GTECH_NOT I_182 ( .A(N2158), .Z(a2stg_shr_tmp8[25]) );
  GTECH_AND2 C4205 ( .A(N2156), .B(N2157), .Z(N2158) );
  GTECH_OR2 C4206 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[25]), .Z(N2156)
         );
  GTECH_OR2 C4207 ( .A(N2054), .B(a2stg_shr_tmp6[29]), .Z(N2157) );
  GTECH_NOT I_183 ( .A(N2161), .Z(a2stg_shr_tmp8[24]) );
  GTECH_AND2 C4210 ( .A(N2159), .B(N2160), .Z(N2161) );
  GTECH_OR2 C4211 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[24]), .Z(N2159)
         );
  GTECH_OR2 C4212 ( .A(N2054), .B(a2stg_shr_tmp6[28]), .Z(N2160) );
  GTECH_NOT I_184 ( .A(N2164), .Z(a2stg_shr_tmp8[23]) );
  GTECH_AND2 C4215 ( .A(N2162), .B(N2163), .Z(N2164) );
  GTECH_OR2 C4216 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[23]), .Z(N2162)
         );
  GTECH_OR2 C4217 ( .A(N2054), .B(a2stg_shr_tmp6[27]), .Z(N2163) );
  GTECH_NOT I_185 ( .A(N2167), .Z(a2stg_shr_tmp8[22]) );
  GTECH_AND2 C4220 ( .A(N2165), .B(N2166), .Z(N2167) );
  GTECH_OR2 C4221 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[22]), .Z(N2165)
         );
  GTECH_OR2 C4222 ( .A(N2054), .B(a2stg_shr_tmp6[26]), .Z(N2166) );
  GTECH_NOT I_186 ( .A(N2170), .Z(a2stg_shr_tmp8[21]) );
  GTECH_AND2 C4225 ( .A(N2168), .B(N2169), .Z(N2170) );
  GTECH_OR2 C4226 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[21]), .Z(N2168)
         );
  GTECH_OR2 C4227 ( .A(N2054), .B(a2stg_shr_tmp6[25]), .Z(N2169) );
  GTECH_NOT I_187 ( .A(N2173), .Z(a2stg_shr_tmp8[20]) );
  GTECH_AND2 C4230 ( .A(N2171), .B(N2172), .Z(N2173) );
  GTECH_OR2 C4231 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[20]), .Z(N2171)
         );
  GTECH_OR2 C4232 ( .A(N2054), .B(a2stg_shr_tmp6[24]), .Z(N2172) );
  GTECH_NOT I_188 ( .A(N2176), .Z(a2stg_shr_tmp8[19]) );
  GTECH_AND2 C4235 ( .A(N2174), .B(N2175), .Z(N2176) );
  GTECH_OR2 C4236 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[19]), .Z(N2174)
         );
  GTECH_OR2 C4237 ( .A(N2054), .B(a2stg_shr_tmp6[23]), .Z(N2175) );
  GTECH_NOT I_189 ( .A(N2179), .Z(a2stg_shr_tmp8[18]) );
  GTECH_AND2 C4240 ( .A(N2177), .B(N2178), .Z(N2179) );
  GTECH_OR2 C4241 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[18]), .Z(N2177)
         );
  GTECH_OR2 C4242 ( .A(N2054), .B(a2stg_shr_tmp6[22]), .Z(N2178) );
  GTECH_NOT I_190 ( .A(N2182), .Z(a2stg_shr_tmp8[17]) );
  GTECH_AND2 C4245 ( .A(N2180), .B(N2181), .Z(N2182) );
  GTECH_OR2 C4246 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[17]), .Z(N2180)
         );
  GTECH_OR2 C4247 ( .A(N2054), .B(a2stg_shr_tmp6[21]), .Z(N2181) );
  GTECH_NOT I_191 ( .A(N2185), .Z(a2stg_shr_tmp8[16]) );
  GTECH_AND2 C4250 ( .A(N2183), .B(N2184), .Z(N2185) );
  GTECH_OR2 C4251 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[16]), .Z(N2183)
         );
  GTECH_OR2 C4252 ( .A(N2054), .B(a2stg_shr_tmp6[20]), .Z(N2184) );
  GTECH_NOT I_192 ( .A(N2188), .Z(a2stg_shr_tmp8[15]) );
  GTECH_AND2 C4255 ( .A(N2186), .B(N2187), .Z(N2188) );
  GTECH_OR2 C4256 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[15]), .Z(N2186)
         );
  GTECH_OR2 C4257 ( .A(N2054), .B(a2stg_shr_tmp6[19]), .Z(N2187) );
  GTECH_NOT I_193 ( .A(N2191), .Z(a2stg_shr_tmp8[14]) );
  GTECH_AND2 C4260 ( .A(N2189), .B(N2190), .Z(N2191) );
  GTECH_OR2 C4261 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[14]), .Z(N2189)
         );
  GTECH_OR2 C4262 ( .A(N2054), .B(a2stg_shr_tmp6[18]), .Z(N2190) );
  GTECH_NOT I_194 ( .A(N2194), .Z(a2stg_shr_tmp8[13]) );
  GTECH_AND2 C4265 ( .A(N2192), .B(N2193), .Z(N2194) );
  GTECH_OR2 C4266 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[13]), .Z(N2192)
         );
  GTECH_OR2 C4267 ( .A(N2054), .B(a2stg_shr_tmp6[17]), .Z(N2193) );
  GTECH_NOT I_195 ( .A(N2197), .Z(a2stg_shr_tmp8[12]) );
  GTECH_AND2 C4270 ( .A(N2195), .B(N2196), .Z(N2197) );
  GTECH_OR2 C4271 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[12]), .Z(N2195)
         );
  GTECH_OR2 C4272 ( .A(N2054), .B(a2stg_shr_tmp6[16]), .Z(N2196) );
  GTECH_NOT I_196 ( .A(N2200), .Z(a2stg_shr_tmp8[11]) );
  GTECH_AND2 C4275 ( .A(N2198), .B(N2199), .Z(N2200) );
  GTECH_OR2 C4276 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[11]), .Z(N2198)
         );
  GTECH_OR2 C4277 ( .A(N2054), .B(a2stg_shr_tmp6[15]), .Z(N2199) );
  GTECH_NOT I_197 ( .A(N2203), .Z(a2stg_shr_tmp8[10]) );
  GTECH_AND2 C4280 ( .A(N2201), .B(N2202), .Z(N2203) );
  GTECH_OR2 C4281 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[10]), .Z(N2201)
         );
  GTECH_OR2 C4282 ( .A(N2054), .B(a2stg_shr_tmp6[14]), .Z(N2202) );
  GTECH_NOT I_198 ( .A(N2206), .Z(a2stg_shr_tmp8[9]) );
  GTECH_AND2 C4285 ( .A(N2204), .B(N2205), .Z(N2206) );
  GTECH_OR2 C4286 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[9]), .Z(N2204)
         );
  GTECH_OR2 C4287 ( .A(N2054), .B(a2stg_shr_tmp6[13]), .Z(N2205) );
  GTECH_NOT I_199 ( .A(N2209), .Z(a2stg_shr_tmp8[8]) );
  GTECH_AND2 C4290 ( .A(N2207), .B(N2208), .Z(N2209) );
  GTECH_OR2 C4291 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[8]), .Z(N2207)
         );
  GTECH_OR2 C4292 ( .A(N2054), .B(a2stg_shr_tmp6[12]), .Z(N2208) );
  GTECH_NOT I_200 ( .A(N2212), .Z(a2stg_shr_tmp8[7]) );
  GTECH_AND2 C4295 ( .A(N2210), .B(N2211), .Z(N2212) );
  GTECH_OR2 C4296 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[7]), .Z(N2210)
         );
  GTECH_OR2 C4297 ( .A(N2054), .B(a2stg_shr_tmp6[11]), .Z(N2211) );
  GTECH_NOT I_201 ( .A(N2215), .Z(a2stg_shr_tmp8[6]) );
  GTECH_AND2 C4300 ( .A(N2213), .B(N2214), .Z(N2215) );
  GTECH_OR2 C4301 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[6]), .Z(N2213)
         );
  GTECH_OR2 C4302 ( .A(N2054), .B(a2stg_shr_tmp6[10]), .Z(N2214) );
  GTECH_NOT I_202 ( .A(N2218), .Z(a2stg_shr_tmp8[5]) );
  GTECH_AND2 C4305 ( .A(N2216), .B(N2217), .Z(N2218) );
  GTECH_OR2 C4306 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[5]), .Z(N2216)
         );
  GTECH_OR2 C4307 ( .A(N2054), .B(a2stg_shr_tmp6[9]), .Z(N2217) );
  GTECH_NOT I_203 ( .A(N2221), .Z(a2stg_shr_tmp8[4]) );
  GTECH_AND2 C4310 ( .A(N2219), .B(N2220), .Z(N2221) );
  GTECH_OR2 C4311 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[4]), .Z(N2219)
         );
  GTECH_OR2 C4312 ( .A(N2054), .B(a2stg_shr_tmp6[8]), .Z(N2220) );
  GTECH_NOT I_204 ( .A(N2224), .Z(a2stg_shr_tmp8[3]) );
  GTECH_AND2 C4315 ( .A(N2222), .B(N2223), .Z(N2224) );
  GTECH_OR2 C4316 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[3]), .Z(N2222)
         );
  GTECH_OR2 C4317 ( .A(N2054), .B(a2stg_shr_tmp6[7]), .Z(N2223) );
  GTECH_NOT I_205 ( .A(N2227), .Z(a2stg_shr_tmp8[2]) );
  GTECH_AND2 C4320 ( .A(N2225), .B(N2226), .Z(N2227) );
  GTECH_OR2 C4321 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[2]), .Z(N2225)
         );
  GTECH_OR2 C4322 ( .A(N2054), .B(a2stg_shr_tmp6[6]), .Z(N2226) );
  GTECH_NOT I_206 ( .A(N2230), .Z(a2stg_shr_tmp8[1]) );
  GTECH_AND2 C4325 ( .A(N2228), .B(N2229), .Z(N2230) );
  GTECH_OR2 C4326 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[1]), .Z(N2228)
         );
  GTECH_OR2 C4327 ( .A(N2054), .B(a2stg_shr_tmp6[5]), .Z(N2229) );
  GTECH_NOT I_207 ( .A(N2233), .Z(a2stg_shr_tmp8[0]) );
  GTECH_AND2 C4330 ( .A(N2231), .B(N2232), .Z(N2233) );
  GTECH_OR2 C4331 ( .A(a2stg_shr_cnt_2[0]), .B(a2stg_shr_tmp6[0]), .Z(N2231)
         );
  GTECH_OR2 C4332 ( .A(N2054), .B(a2stg_shr_tmp6[4]), .Z(N2232) );
  GTECH_NOT I_208 ( .A(N2235), .Z(a2stg_shr_tmp10[63]) );
  GTECH_AND2 C4335 ( .A(N2234), .B(a2stg_shr_tmp8[63]), .Z(N2235) );
  GTECH_NOT I_209 ( .A(a2stg_shr_cnt_1[1]), .Z(N2234) );
  GTECH_NOT I_210 ( .A(N2236), .Z(a2stg_shr_tmp10[62]) );
  GTECH_AND2 C4338 ( .A(N2234), .B(a2stg_shr_tmp8[62]), .Z(N2236) );
  GTECH_NOT I_211 ( .A(N2239), .Z(a2stg_shr_tmp10[61]) );
  GTECH_OR2 C4341 ( .A(N2237), .B(N2238), .Z(N2239) );
  GTECH_AND2 C4342 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[63]), .Z(N2237)
         );
  GTECH_AND2 C4343 ( .A(N2234), .B(a2stg_shr_tmp8[61]), .Z(N2238) );
  GTECH_NOT I_212 ( .A(N2242), .Z(a2stg_shr_tmp10[60]) );
  GTECH_OR2 C4346 ( .A(N2240), .B(N2241), .Z(N2242) );
  GTECH_AND2 C4347 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[62]), .Z(N2240)
         );
  GTECH_AND2 C4348 ( .A(N2234), .B(a2stg_shr_tmp8[60]), .Z(N2241) );
  GTECH_NOT I_213 ( .A(N2245), .Z(a2stg_shr_tmp10[59]) );
  GTECH_OR2 C4351 ( .A(N2243), .B(N2244), .Z(N2245) );
  GTECH_AND2 C4352 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[61]), .Z(N2243)
         );
  GTECH_AND2 C4353 ( .A(N2234), .B(a2stg_shr_tmp8[59]), .Z(N2244) );
  GTECH_NOT I_214 ( .A(N2248), .Z(a2stg_shr_tmp10[58]) );
  GTECH_OR2 C4356 ( .A(N2246), .B(N2247), .Z(N2248) );
  GTECH_AND2 C4357 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[60]), .Z(N2246)
         );
  GTECH_AND2 C4358 ( .A(N2234), .B(a2stg_shr_tmp8[58]), .Z(N2247) );
  GTECH_NOT I_215 ( .A(N2251), .Z(a2stg_shr_tmp10[57]) );
  GTECH_OR2 C4361 ( .A(N2249), .B(N2250), .Z(N2251) );
  GTECH_AND2 C4362 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[59]), .Z(N2249)
         );
  GTECH_AND2 C4363 ( .A(N2234), .B(a2stg_shr_tmp8[57]), .Z(N2250) );
  GTECH_NOT I_216 ( .A(N2254), .Z(a2stg_shr_tmp10[56]) );
  GTECH_OR2 C4366 ( .A(N2252), .B(N2253), .Z(N2254) );
  GTECH_AND2 C4367 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[58]), .Z(N2252)
         );
  GTECH_AND2 C4368 ( .A(N2234), .B(a2stg_shr_tmp8[56]), .Z(N2253) );
  GTECH_NOT I_217 ( .A(N2257), .Z(a2stg_shr_tmp10[55]) );
  GTECH_OR2 C4371 ( .A(N2255), .B(N2256), .Z(N2257) );
  GTECH_AND2 C4372 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[57]), .Z(N2255)
         );
  GTECH_AND2 C4373 ( .A(N2234), .B(a2stg_shr_tmp8[55]), .Z(N2256) );
  GTECH_NOT I_218 ( .A(N2260), .Z(a2stg_shr_tmp10[54]) );
  GTECH_OR2 C4376 ( .A(N2258), .B(N2259), .Z(N2260) );
  GTECH_AND2 C4377 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[56]), .Z(N2258)
         );
  GTECH_AND2 C4378 ( .A(N2234), .B(a2stg_shr_tmp8[54]), .Z(N2259) );
  GTECH_NOT I_219 ( .A(N2263), .Z(a2stg_shr_tmp10[53]) );
  GTECH_OR2 C4381 ( .A(N2261), .B(N2262), .Z(N2263) );
  GTECH_AND2 C4382 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[55]), .Z(N2261)
         );
  GTECH_AND2 C4383 ( .A(N2234), .B(a2stg_shr_tmp8[53]), .Z(N2262) );
  GTECH_NOT I_220 ( .A(N2266), .Z(a2stg_shr_tmp10[52]) );
  GTECH_OR2 C4386 ( .A(N2264), .B(N2265), .Z(N2266) );
  GTECH_AND2 C4387 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[54]), .Z(N2264)
         );
  GTECH_AND2 C4388 ( .A(N2234), .B(a2stg_shr_tmp8[52]), .Z(N2265) );
  GTECH_NOT I_221 ( .A(N2269), .Z(a2stg_shr_tmp10[51]) );
  GTECH_OR2 C4391 ( .A(N2267), .B(N2268), .Z(N2269) );
  GTECH_AND2 C4392 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[53]), .Z(N2267)
         );
  GTECH_AND2 C4393 ( .A(N2234), .B(a2stg_shr_tmp8[51]), .Z(N2268) );
  GTECH_NOT I_222 ( .A(N2272), .Z(a2stg_shr_tmp10[50]) );
  GTECH_OR2 C4396 ( .A(N2270), .B(N2271), .Z(N2272) );
  GTECH_AND2 C4397 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[52]), .Z(N2270)
         );
  GTECH_AND2 C4398 ( .A(N2234), .B(a2stg_shr_tmp8[50]), .Z(N2271) );
  GTECH_NOT I_223 ( .A(N2275), .Z(a2stg_shr_tmp10[49]) );
  GTECH_OR2 C4401 ( .A(N2273), .B(N2274), .Z(N2275) );
  GTECH_AND2 C4402 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[51]), .Z(N2273)
         );
  GTECH_AND2 C4403 ( .A(N2234), .B(a2stg_shr_tmp8[49]), .Z(N2274) );
  GTECH_NOT I_224 ( .A(N2278), .Z(a2stg_shr_tmp10[48]) );
  GTECH_OR2 C4406 ( .A(N2276), .B(N2277), .Z(N2278) );
  GTECH_AND2 C4407 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[50]), .Z(N2276)
         );
  GTECH_AND2 C4408 ( .A(N2234), .B(a2stg_shr_tmp8[48]), .Z(N2277) );
  GTECH_NOT I_225 ( .A(N2281), .Z(a2stg_shr_tmp10[47]) );
  GTECH_OR2 C4411 ( .A(N2279), .B(N2280), .Z(N2281) );
  GTECH_AND2 C4412 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[49]), .Z(N2279)
         );
  GTECH_AND2 C4413 ( .A(N2234), .B(a2stg_shr_tmp8[47]), .Z(N2280) );
  GTECH_NOT I_226 ( .A(N2284), .Z(a2stg_shr_tmp10[46]) );
  GTECH_OR2 C4416 ( .A(N2282), .B(N2283), .Z(N2284) );
  GTECH_AND2 C4417 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[48]), .Z(N2282)
         );
  GTECH_AND2 C4418 ( .A(N2234), .B(a2stg_shr_tmp8[46]), .Z(N2283) );
  GTECH_NOT I_227 ( .A(N2287), .Z(a2stg_shr_tmp10[45]) );
  GTECH_OR2 C4421 ( .A(N2285), .B(N2286), .Z(N2287) );
  GTECH_AND2 C4422 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[47]), .Z(N2285)
         );
  GTECH_AND2 C4423 ( .A(N2234), .B(a2stg_shr_tmp8[45]), .Z(N2286) );
  GTECH_NOT I_228 ( .A(N2290), .Z(a2stg_shr_tmp10[44]) );
  GTECH_OR2 C4426 ( .A(N2288), .B(N2289), .Z(N2290) );
  GTECH_AND2 C4427 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[46]), .Z(N2288)
         );
  GTECH_AND2 C4428 ( .A(N2234), .B(a2stg_shr_tmp8[44]), .Z(N2289) );
  GTECH_NOT I_229 ( .A(N2293), .Z(a2stg_shr_tmp10[43]) );
  GTECH_OR2 C4431 ( .A(N2291), .B(N2292), .Z(N2293) );
  GTECH_AND2 C4432 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[45]), .Z(N2291)
         );
  GTECH_AND2 C4433 ( .A(N2234), .B(a2stg_shr_tmp8[43]), .Z(N2292) );
  GTECH_NOT I_230 ( .A(N2296), .Z(a2stg_shr_tmp10[42]) );
  GTECH_OR2 C4436 ( .A(N2294), .B(N2295), .Z(N2296) );
  GTECH_AND2 C4437 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[44]), .Z(N2294)
         );
  GTECH_AND2 C4438 ( .A(N2234), .B(a2stg_shr_tmp8[42]), .Z(N2295) );
  GTECH_NOT I_231 ( .A(N2299), .Z(a2stg_shr_tmp10[41]) );
  GTECH_OR2 C4441 ( .A(N2297), .B(N2298), .Z(N2299) );
  GTECH_AND2 C4442 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[43]), .Z(N2297)
         );
  GTECH_AND2 C4443 ( .A(N2234), .B(a2stg_shr_tmp8[41]), .Z(N2298) );
  GTECH_NOT I_232 ( .A(N2302), .Z(a2stg_shr_tmp10[40]) );
  GTECH_OR2 C4446 ( .A(N2300), .B(N2301), .Z(N2302) );
  GTECH_AND2 C4447 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[42]), .Z(N2300)
         );
  GTECH_AND2 C4448 ( .A(N2234), .B(a2stg_shr_tmp8[40]), .Z(N2301) );
  GTECH_NOT I_233 ( .A(N2305), .Z(a2stg_shr_tmp10[39]) );
  GTECH_OR2 C4451 ( .A(N2303), .B(N2304), .Z(N2305) );
  GTECH_AND2 C4452 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[41]), .Z(N2303)
         );
  GTECH_AND2 C4453 ( .A(N2234), .B(a2stg_shr_tmp8[39]), .Z(N2304) );
  GTECH_NOT I_234 ( .A(N2308), .Z(a2stg_shr_tmp10[38]) );
  GTECH_OR2 C4456 ( .A(N2306), .B(N2307), .Z(N2308) );
  GTECH_AND2 C4457 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[40]), .Z(N2306)
         );
  GTECH_AND2 C4458 ( .A(N2234), .B(a2stg_shr_tmp8[38]), .Z(N2307) );
  GTECH_NOT I_235 ( .A(N2311), .Z(a2stg_shr_tmp10[37]) );
  GTECH_OR2 C4461 ( .A(N2309), .B(N2310), .Z(N2311) );
  GTECH_AND2 C4462 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[39]), .Z(N2309)
         );
  GTECH_AND2 C4463 ( .A(N2234), .B(a2stg_shr_tmp8[37]), .Z(N2310) );
  GTECH_NOT I_236 ( .A(N2314), .Z(a2stg_shr_tmp10[36]) );
  GTECH_OR2 C4466 ( .A(N2312), .B(N2313), .Z(N2314) );
  GTECH_AND2 C4467 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[38]), .Z(N2312)
         );
  GTECH_AND2 C4468 ( .A(N2234), .B(a2stg_shr_tmp8[36]), .Z(N2313) );
  GTECH_NOT I_237 ( .A(N2317), .Z(a2stg_shr_tmp10[35]) );
  GTECH_OR2 C4471 ( .A(N2315), .B(N2316), .Z(N2317) );
  GTECH_AND2 C4472 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[37]), .Z(N2315)
         );
  GTECH_AND2 C4473 ( .A(N2234), .B(a2stg_shr_tmp8[35]), .Z(N2316) );
  GTECH_NOT I_238 ( .A(N2320), .Z(a2stg_shr_tmp10[34]) );
  GTECH_OR2 C4476 ( .A(N2318), .B(N2319), .Z(N2320) );
  GTECH_AND2 C4477 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[36]), .Z(N2318)
         );
  GTECH_AND2 C4478 ( .A(N2234), .B(a2stg_shr_tmp8[34]), .Z(N2319) );
  GTECH_NOT I_239 ( .A(N2323), .Z(a2stg_shr_tmp10[33]) );
  GTECH_OR2 C4481 ( .A(N2321), .B(N2322), .Z(N2323) );
  GTECH_AND2 C4482 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[35]), .Z(N2321)
         );
  GTECH_AND2 C4483 ( .A(N2234), .B(a2stg_shr_tmp8[33]), .Z(N2322) );
  GTECH_NOT I_240 ( .A(N2326), .Z(a2stg_shr_tmp10[32]) );
  GTECH_OR2 C4486 ( .A(N2324), .B(N2325), .Z(N2326) );
  GTECH_AND2 C4487 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[34]), .Z(N2324)
         );
  GTECH_AND2 C4488 ( .A(N2234), .B(a2stg_shr_tmp8[32]), .Z(N2325) );
  GTECH_NOT I_241 ( .A(N2329), .Z(a2stg_shr_tmp10[31]) );
  GTECH_OR2 C4491 ( .A(N2327), .B(N2328), .Z(N2329) );
  GTECH_AND2 C4492 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[33]), .Z(N2327)
         );
  GTECH_AND2 C4493 ( .A(N2234), .B(a2stg_shr_tmp8[31]), .Z(N2328) );
  GTECH_NOT I_242 ( .A(N2332), .Z(a2stg_shr_tmp10[30]) );
  GTECH_OR2 C4496 ( .A(N2330), .B(N2331), .Z(N2332) );
  GTECH_AND2 C4497 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[32]), .Z(N2330)
         );
  GTECH_AND2 C4498 ( .A(N2234), .B(a2stg_shr_tmp8[30]), .Z(N2331) );
  GTECH_NOT I_243 ( .A(N2335), .Z(a2stg_shr_tmp10[29]) );
  GTECH_OR2 C4501 ( .A(N2333), .B(N2334), .Z(N2335) );
  GTECH_AND2 C4502 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[31]), .Z(N2333)
         );
  GTECH_AND2 C4503 ( .A(N2234), .B(a2stg_shr_tmp8[29]), .Z(N2334) );
  GTECH_NOT I_244 ( .A(N2338), .Z(a2stg_shr_tmp10[28]) );
  GTECH_OR2 C4506 ( .A(N2336), .B(N2337), .Z(N2338) );
  GTECH_AND2 C4507 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[30]), .Z(N2336)
         );
  GTECH_AND2 C4508 ( .A(N2234), .B(a2stg_shr_tmp8[28]), .Z(N2337) );
  GTECH_NOT I_245 ( .A(N2341), .Z(a2stg_shr_tmp10[27]) );
  GTECH_OR2 C4511 ( .A(N2339), .B(N2340), .Z(N2341) );
  GTECH_AND2 C4512 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[29]), .Z(N2339)
         );
  GTECH_AND2 C4513 ( .A(N2234), .B(a2stg_shr_tmp8[27]), .Z(N2340) );
  GTECH_NOT I_246 ( .A(N2344), .Z(a2stg_shr_tmp10[26]) );
  GTECH_OR2 C4516 ( .A(N2342), .B(N2343), .Z(N2344) );
  GTECH_AND2 C4517 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[28]), .Z(N2342)
         );
  GTECH_AND2 C4518 ( .A(N2234), .B(a2stg_shr_tmp8[26]), .Z(N2343) );
  GTECH_NOT I_247 ( .A(N2347), .Z(a2stg_shr_tmp10[25]) );
  GTECH_OR2 C4521 ( .A(N2345), .B(N2346), .Z(N2347) );
  GTECH_AND2 C4522 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[27]), .Z(N2345)
         );
  GTECH_AND2 C4523 ( .A(N2234), .B(a2stg_shr_tmp8[25]), .Z(N2346) );
  GTECH_NOT I_248 ( .A(N2350), .Z(a2stg_shr_tmp10[24]) );
  GTECH_OR2 C4526 ( .A(N2348), .B(N2349), .Z(N2350) );
  GTECH_AND2 C4527 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[26]), .Z(N2348)
         );
  GTECH_AND2 C4528 ( .A(N2234), .B(a2stg_shr_tmp8[24]), .Z(N2349) );
  GTECH_NOT I_249 ( .A(N2353), .Z(a2stg_shr_tmp10[23]) );
  GTECH_OR2 C4531 ( .A(N2351), .B(N2352), .Z(N2353) );
  GTECH_AND2 C4532 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[25]), .Z(N2351)
         );
  GTECH_AND2 C4533 ( .A(N2234), .B(a2stg_shr_tmp8[23]), .Z(N2352) );
  GTECH_NOT I_250 ( .A(N2356), .Z(a2stg_shr_tmp10[22]) );
  GTECH_OR2 C4536 ( .A(N2354), .B(N2355), .Z(N2356) );
  GTECH_AND2 C4537 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[24]), .Z(N2354)
         );
  GTECH_AND2 C4538 ( .A(N2234), .B(a2stg_shr_tmp8[22]), .Z(N2355) );
  GTECH_NOT I_251 ( .A(N2359), .Z(a2stg_shr_tmp10[21]) );
  GTECH_OR2 C4541 ( .A(N2357), .B(N2358), .Z(N2359) );
  GTECH_AND2 C4542 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[23]), .Z(N2357)
         );
  GTECH_AND2 C4543 ( .A(N2234), .B(a2stg_shr_tmp8[21]), .Z(N2358) );
  GTECH_NOT I_252 ( .A(N2362), .Z(a2stg_shr_tmp10[20]) );
  GTECH_OR2 C4546 ( .A(N2360), .B(N2361), .Z(N2362) );
  GTECH_AND2 C4547 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[22]), .Z(N2360)
         );
  GTECH_AND2 C4548 ( .A(N2234), .B(a2stg_shr_tmp8[20]), .Z(N2361) );
  GTECH_NOT I_253 ( .A(N2365), .Z(a2stg_shr_tmp10[19]) );
  GTECH_OR2 C4551 ( .A(N2363), .B(N2364), .Z(N2365) );
  GTECH_AND2 C4552 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[21]), .Z(N2363)
         );
  GTECH_AND2 C4553 ( .A(N2234), .B(a2stg_shr_tmp8[19]), .Z(N2364) );
  GTECH_NOT I_254 ( .A(N2368), .Z(a2stg_shr_tmp10[18]) );
  GTECH_OR2 C4556 ( .A(N2366), .B(N2367), .Z(N2368) );
  GTECH_AND2 C4557 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[20]), .Z(N2366)
         );
  GTECH_AND2 C4558 ( .A(N2234), .B(a2stg_shr_tmp8[18]), .Z(N2367) );
  GTECH_NOT I_255 ( .A(N2371), .Z(a2stg_shr_tmp10[17]) );
  GTECH_OR2 C4561 ( .A(N2369), .B(N2370), .Z(N2371) );
  GTECH_AND2 C4562 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[19]), .Z(N2369)
         );
  GTECH_AND2 C4563 ( .A(N2234), .B(a2stg_shr_tmp8[17]), .Z(N2370) );
  GTECH_NOT I_256 ( .A(N2374), .Z(a2stg_shr_tmp10[16]) );
  GTECH_OR2 C4566 ( .A(N2372), .B(N2373), .Z(N2374) );
  GTECH_AND2 C4567 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[18]), .Z(N2372)
         );
  GTECH_AND2 C4568 ( .A(N2234), .B(a2stg_shr_tmp8[16]), .Z(N2373) );
  GTECH_NOT I_257 ( .A(N2377), .Z(a2stg_shr_tmp10[15]) );
  GTECH_OR2 C4571 ( .A(N2375), .B(N2376), .Z(N2377) );
  GTECH_AND2 C4572 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[17]), .Z(N2375)
         );
  GTECH_AND2 C4573 ( .A(N2234), .B(a2stg_shr_tmp8[15]), .Z(N2376) );
  GTECH_NOT I_258 ( .A(N2380), .Z(a2stg_shr_tmp10[14]) );
  GTECH_OR2 C4576 ( .A(N2378), .B(N2379), .Z(N2380) );
  GTECH_AND2 C4577 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[16]), .Z(N2378)
         );
  GTECH_AND2 C4578 ( .A(N2234), .B(a2stg_shr_tmp8[14]), .Z(N2379) );
  GTECH_NOT I_259 ( .A(N2383), .Z(a2stg_shr_tmp10[13]) );
  GTECH_OR2 C4581 ( .A(N2381), .B(N2382), .Z(N2383) );
  GTECH_AND2 C4582 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[15]), .Z(N2381)
         );
  GTECH_AND2 C4583 ( .A(N2234), .B(a2stg_shr_tmp8[13]), .Z(N2382) );
  GTECH_NOT I_260 ( .A(N2386), .Z(a2stg_shr_tmp10[12]) );
  GTECH_OR2 C4586 ( .A(N2384), .B(N2385), .Z(N2386) );
  GTECH_AND2 C4587 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[14]), .Z(N2384)
         );
  GTECH_AND2 C4588 ( .A(N2234), .B(a2stg_shr_tmp8[12]), .Z(N2385) );
  GTECH_NOT I_261 ( .A(N2389), .Z(a2stg_shr_tmp10[11]) );
  GTECH_OR2 C4591 ( .A(N2387), .B(N2388), .Z(N2389) );
  GTECH_AND2 C4592 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[13]), .Z(N2387)
         );
  GTECH_AND2 C4593 ( .A(N2234), .B(a2stg_shr_tmp8[11]), .Z(N2388) );
  GTECH_NOT I_262 ( .A(N2392), .Z(a2stg_shr_tmp10[10]) );
  GTECH_OR2 C4596 ( .A(N2390), .B(N2391), .Z(N2392) );
  GTECH_AND2 C4597 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[12]), .Z(N2390)
         );
  GTECH_AND2 C4598 ( .A(N2234), .B(a2stg_shr_tmp8[10]), .Z(N2391) );
  GTECH_NOT I_263 ( .A(N2395), .Z(a2stg_shr_tmp10[9]) );
  GTECH_OR2 C4601 ( .A(N2393), .B(N2394), .Z(N2395) );
  GTECH_AND2 C4602 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[11]), .Z(N2393)
         );
  GTECH_AND2 C4603 ( .A(N2234), .B(a2stg_shr_tmp8[9]), .Z(N2394) );
  GTECH_NOT I_264 ( .A(N2398), .Z(a2stg_shr_tmp10[8]) );
  GTECH_OR2 C4606 ( .A(N2396), .B(N2397), .Z(N2398) );
  GTECH_AND2 C4607 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[10]), .Z(N2396)
         );
  GTECH_AND2 C4608 ( .A(N2234), .B(a2stg_shr_tmp8[8]), .Z(N2397) );
  GTECH_NOT I_265 ( .A(N2401), .Z(a2stg_shr_tmp10[7]) );
  GTECH_OR2 C4611 ( .A(N2399), .B(N2400), .Z(N2401) );
  GTECH_AND2 C4612 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[9]), .Z(N2399)
         );
  GTECH_AND2 C4613 ( .A(N2234), .B(a2stg_shr_tmp8[7]), .Z(N2400) );
  GTECH_NOT I_266 ( .A(N2404), .Z(a2stg_shr_tmp10[6]) );
  GTECH_OR2 C4616 ( .A(N2402), .B(N2403), .Z(N2404) );
  GTECH_AND2 C4617 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[8]), .Z(N2402)
         );
  GTECH_AND2 C4618 ( .A(N2234), .B(a2stg_shr_tmp8[6]), .Z(N2403) );
  GTECH_NOT I_267 ( .A(N2407), .Z(a2stg_shr_tmp10[5]) );
  GTECH_OR2 C4621 ( .A(N2405), .B(N2406), .Z(N2407) );
  GTECH_AND2 C4622 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[7]), .Z(N2405)
         );
  GTECH_AND2 C4623 ( .A(N2234), .B(a2stg_shr_tmp8[5]), .Z(N2406) );
  GTECH_NOT I_268 ( .A(N2410), .Z(a2stg_shr_tmp10[4]) );
  GTECH_OR2 C4626 ( .A(N2408), .B(N2409), .Z(N2410) );
  GTECH_AND2 C4627 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[6]), .Z(N2408)
         );
  GTECH_AND2 C4628 ( .A(N2234), .B(a2stg_shr_tmp8[4]), .Z(N2409) );
  GTECH_NOT I_269 ( .A(N2413), .Z(a2stg_shr_tmp10[3]) );
  GTECH_OR2 C4631 ( .A(N2411), .B(N2412), .Z(N2413) );
  GTECH_AND2 C4632 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[5]), .Z(N2411)
         );
  GTECH_AND2 C4633 ( .A(N2234), .B(a2stg_shr_tmp8[3]), .Z(N2412) );
  GTECH_NOT I_270 ( .A(N2416), .Z(a2stg_shr_tmp10[2]) );
  GTECH_OR2 C4636 ( .A(N2414), .B(N2415), .Z(N2416) );
  GTECH_AND2 C4637 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[4]), .Z(N2414)
         );
  GTECH_AND2 C4638 ( .A(N2234), .B(a2stg_shr_tmp8[2]), .Z(N2415) );
  GTECH_NOT I_271 ( .A(N2419), .Z(a2stg_shr_tmp10[1]) );
  GTECH_OR2 C4641 ( .A(N2417), .B(N2418), .Z(N2419) );
  GTECH_AND2 C4642 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[3]), .Z(N2417)
         );
  GTECH_AND2 C4643 ( .A(N2234), .B(a2stg_shr_tmp8[1]), .Z(N2418) );
  GTECH_NOT I_272 ( .A(N2422), .Z(a2stg_shr_tmp10[0]) );
  GTECH_OR2 C4646 ( .A(N2420), .B(N2421), .Z(N2422) );
  GTECH_AND2 C4647 ( .A(a2stg_shr_cnt_1[0]), .B(a2stg_shr_tmp8[2]), .Z(N2420)
         );
  GTECH_AND2 C4648 ( .A(N2234), .B(a2stg_shr_tmp8[0]), .Z(N2421) );
  GTECH_NOT I_273 ( .A(N2423), .Z(a2stg_shr[115]) );
  GTECH_OR2 C4651 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[63]), .Z(N2423)
         );
  GTECH_NOT I_274 ( .A(N2427), .Z(a2stg_shr[114]) );
  GTECH_AND2 C4653 ( .A(N2424), .B(N2426), .Z(N2427) );
  GTECH_OR2 C4654 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[62]), .Z(N2424)
         );
  GTECH_OR2 C4655 ( .A(N2425), .B(a2stg_shr_tmp10[63]), .Z(N2426) );
  GTECH_NOT I_275 ( .A(a2stg_shr_cnt_0[1]), .Z(N2425) );
  GTECH_NOT I_276 ( .A(N2430), .Z(a2stg_shr[113]) );
  GTECH_AND2 C4658 ( .A(N2428), .B(N2429), .Z(N2430) );
  GTECH_OR2 C4659 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[61]), .Z(N2428)
         );
  GTECH_OR2 C4660 ( .A(N2425), .B(a2stg_shr_tmp10[62]), .Z(N2429) );
  GTECH_NOT I_277 ( .A(N2433), .Z(a2stg_shr[112]) );
  GTECH_AND2 C4663 ( .A(N2431), .B(N2432), .Z(N2433) );
  GTECH_OR2 C4664 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[60]), .Z(N2431)
         );
  GTECH_OR2 C4665 ( .A(N2425), .B(a2stg_shr_tmp10[61]), .Z(N2432) );
  GTECH_NOT I_278 ( .A(N2436), .Z(a2stg_shr[111]) );
  GTECH_AND2 C4668 ( .A(N2434), .B(N2435), .Z(N2436) );
  GTECH_OR2 C4669 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[59]), .Z(N2434)
         );
  GTECH_OR2 C4670 ( .A(N2425), .B(a2stg_shr_tmp10[60]), .Z(N2435) );
  GTECH_NOT I_279 ( .A(N2439), .Z(a2stg_shr[110]) );
  GTECH_AND2 C4673 ( .A(N2437), .B(N2438), .Z(N2439) );
  GTECH_OR2 C4674 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[58]), .Z(N2437)
         );
  GTECH_OR2 C4675 ( .A(N2425), .B(a2stg_shr_tmp10[59]), .Z(N2438) );
  GTECH_NOT I_280 ( .A(N2442), .Z(a2stg_shr[109]) );
  GTECH_AND2 C4678 ( .A(N2440), .B(N2441), .Z(N2442) );
  GTECH_OR2 C4679 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[57]), .Z(N2440)
         );
  GTECH_OR2 C4680 ( .A(N2425), .B(a2stg_shr_tmp10[58]), .Z(N2441) );
  GTECH_NOT I_281 ( .A(N2445), .Z(a2stg_shr[108]) );
  GTECH_AND2 C4683 ( .A(N2443), .B(N2444), .Z(N2445) );
  GTECH_OR2 C4684 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[56]), .Z(N2443)
         );
  GTECH_OR2 C4685 ( .A(N2425), .B(a2stg_shr_tmp10[57]), .Z(N2444) );
  GTECH_NOT I_282 ( .A(N2448), .Z(a2stg_shr[107]) );
  GTECH_AND2 C4688 ( .A(N2446), .B(N2447), .Z(N2448) );
  GTECH_OR2 C4689 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[55]), .Z(N2446)
         );
  GTECH_OR2 C4690 ( .A(N2425), .B(a2stg_shr_tmp10[56]), .Z(N2447) );
  GTECH_NOT I_283 ( .A(N2451), .Z(a2stg_shr[106]) );
  GTECH_AND2 C4693 ( .A(N2449), .B(N2450), .Z(N2451) );
  GTECH_OR2 C4694 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[54]), .Z(N2449)
         );
  GTECH_OR2 C4695 ( .A(N2425), .B(a2stg_shr_tmp10[55]), .Z(N2450) );
  GTECH_NOT I_284 ( .A(N2454), .Z(a2stg_shr[105]) );
  GTECH_AND2 C4698 ( .A(N2452), .B(N2453), .Z(N2454) );
  GTECH_OR2 C4699 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[53]), .Z(N2452)
         );
  GTECH_OR2 C4700 ( .A(N2425), .B(a2stg_shr_tmp10[54]), .Z(N2453) );
  GTECH_NOT I_285 ( .A(N2457), .Z(a2stg_shr[104]) );
  GTECH_AND2 C4703 ( .A(N2455), .B(N2456), .Z(N2457) );
  GTECH_OR2 C4704 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[52]), .Z(N2455)
         );
  GTECH_OR2 C4705 ( .A(N2425), .B(a2stg_shr_tmp10[53]), .Z(N2456) );
  GTECH_NOT I_286 ( .A(N2460), .Z(a2stg_shr[103]) );
  GTECH_AND2 C4708 ( .A(N2458), .B(N2459), .Z(N2460) );
  GTECH_OR2 C4709 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[51]), .Z(N2458)
         );
  GTECH_OR2 C4710 ( .A(N2425), .B(a2stg_shr_tmp10[52]), .Z(N2459) );
  GTECH_NOT I_287 ( .A(N2463), .Z(a2stg_shr[102]) );
  GTECH_AND2 C4713 ( .A(N2461), .B(N2462), .Z(N2463) );
  GTECH_OR2 C4714 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[50]), .Z(N2461)
         );
  GTECH_OR2 C4715 ( .A(N2425), .B(a2stg_shr_tmp10[51]), .Z(N2462) );
  GTECH_NOT I_288 ( .A(N2466), .Z(a2stg_shr[101]) );
  GTECH_AND2 C4718 ( .A(N2464), .B(N2465), .Z(N2466) );
  GTECH_OR2 C4719 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[49]), .Z(N2464)
         );
  GTECH_OR2 C4720 ( .A(N2425), .B(a2stg_shr_tmp10[50]), .Z(N2465) );
  GTECH_NOT I_289 ( .A(N2469), .Z(a2stg_shr[100]) );
  GTECH_AND2 C4723 ( .A(N2467), .B(N2468), .Z(N2469) );
  GTECH_OR2 C4724 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[48]), .Z(N2467)
         );
  GTECH_OR2 C4725 ( .A(N2425), .B(a2stg_shr_tmp10[49]), .Z(N2468) );
  GTECH_NOT I_290 ( .A(N2472), .Z(a2stg_shr[99]) );
  GTECH_AND2 C4728 ( .A(N2470), .B(N2471), .Z(N2472) );
  GTECH_OR2 C4729 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[47]), .Z(N2470)
         );
  GTECH_OR2 C4730 ( .A(N2425), .B(a2stg_shr_tmp10[48]), .Z(N2471) );
  GTECH_NOT I_291 ( .A(N2475), .Z(a2stg_shr[98]) );
  GTECH_AND2 C4733 ( .A(N2473), .B(N2474), .Z(N2475) );
  GTECH_OR2 C4734 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[46]), .Z(N2473)
         );
  GTECH_OR2 C4735 ( .A(N2425), .B(a2stg_shr_tmp10[47]), .Z(N2474) );
  GTECH_NOT I_292 ( .A(N2478), .Z(a2stg_shr[97]) );
  GTECH_AND2 C4738 ( .A(N2476), .B(N2477), .Z(N2478) );
  GTECH_OR2 C4739 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[45]), .Z(N2476)
         );
  GTECH_OR2 C4740 ( .A(N2425), .B(a2stg_shr_tmp10[46]), .Z(N2477) );
  GTECH_NOT I_293 ( .A(N2481), .Z(a2stg_shr[96]) );
  GTECH_AND2 C4743 ( .A(N2479), .B(N2480), .Z(N2481) );
  GTECH_OR2 C4744 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[44]), .Z(N2479)
         );
  GTECH_OR2 C4745 ( .A(N2425), .B(a2stg_shr_tmp10[45]), .Z(N2480) );
  GTECH_NOT I_294 ( .A(N2484), .Z(a2stg_shr[95]) );
  GTECH_AND2 C4748 ( .A(N2482), .B(N2483), .Z(N2484) );
  GTECH_OR2 C4749 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[43]), .Z(N2482)
         );
  GTECH_OR2 C4750 ( .A(N2425), .B(a2stg_shr_tmp10[44]), .Z(N2483) );
  GTECH_NOT I_295 ( .A(N2487), .Z(a2stg_shr[94]) );
  GTECH_AND2 C4753 ( .A(N2485), .B(N2486), .Z(N2487) );
  GTECH_OR2 C4754 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[42]), .Z(N2485)
         );
  GTECH_OR2 C4755 ( .A(N2425), .B(a2stg_shr_tmp10[43]), .Z(N2486) );
  GTECH_NOT I_296 ( .A(N2490), .Z(a2stg_shr[93]) );
  GTECH_AND2 C4758 ( .A(N2488), .B(N2489), .Z(N2490) );
  GTECH_OR2 C4759 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[41]), .Z(N2488)
         );
  GTECH_OR2 C4760 ( .A(N2425), .B(a2stg_shr_tmp10[42]), .Z(N2489) );
  GTECH_NOT I_297 ( .A(N2493), .Z(a2stg_shr[92]) );
  GTECH_AND2 C4763 ( .A(N2491), .B(N2492), .Z(N2493) );
  GTECH_OR2 C4764 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[40]), .Z(N2491)
         );
  GTECH_OR2 C4765 ( .A(N2425), .B(a2stg_shr_tmp10[41]), .Z(N2492) );
  GTECH_NOT I_298 ( .A(N2496), .Z(a2stg_shr[91]) );
  GTECH_AND2 C4768 ( .A(N2494), .B(N2495), .Z(N2496) );
  GTECH_OR2 C4769 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[39]), .Z(N2494)
         );
  GTECH_OR2 C4770 ( .A(N2425), .B(a2stg_shr_tmp10[40]), .Z(N2495) );
  GTECH_NOT I_299 ( .A(N2499), .Z(a2stg_shr[90]) );
  GTECH_AND2 C4773 ( .A(N2497), .B(N2498), .Z(N2499) );
  GTECH_OR2 C4774 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[38]), .Z(N2497)
         );
  GTECH_OR2 C4775 ( .A(N2425), .B(a2stg_shr_tmp10[39]), .Z(N2498) );
  GTECH_NOT I_300 ( .A(N2502), .Z(a2stg_shr[89]) );
  GTECH_AND2 C4778 ( .A(N2500), .B(N2501), .Z(N2502) );
  GTECH_OR2 C4779 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[37]), .Z(N2500)
         );
  GTECH_OR2 C4780 ( .A(N2425), .B(a2stg_shr_tmp10[38]), .Z(N2501) );
  GTECH_NOT I_301 ( .A(N2505), .Z(a2stg_shr[88]) );
  GTECH_AND2 C4783 ( .A(N2503), .B(N2504), .Z(N2505) );
  GTECH_OR2 C4784 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[36]), .Z(N2503)
         );
  GTECH_OR2 C4785 ( .A(N2425), .B(a2stg_shr_tmp10[37]), .Z(N2504) );
  GTECH_NOT I_302 ( .A(N2508), .Z(a2stg_shr[87]) );
  GTECH_AND2 C4788 ( .A(N2506), .B(N2507), .Z(N2508) );
  GTECH_OR2 C4789 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[35]), .Z(N2506)
         );
  GTECH_OR2 C4790 ( .A(N2425), .B(a2stg_shr_tmp10[36]), .Z(N2507) );
  GTECH_NOT I_303 ( .A(N2511), .Z(a2stg_shr[86]) );
  GTECH_AND2 C4793 ( .A(N2509), .B(N2510), .Z(N2511) );
  GTECH_OR2 C4794 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[34]), .Z(N2509)
         );
  GTECH_OR2 C4795 ( .A(N2425), .B(a2stg_shr_tmp10[35]), .Z(N2510) );
  GTECH_NOT I_304 ( .A(N2514), .Z(a2stg_shr[85]) );
  GTECH_AND2 C4798 ( .A(N2512), .B(N2513), .Z(N2514) );
  GTECH_OR2 C4799 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[33]), .Z(N2512)
         );
  GTECH_OR2 C4800 ( .A(N2425), .B(a2stg_shr_tmp10[34]), .Z(N2513) );
  GTECH_NOT I_305 ( .A(N2517), .Z(a2stg_shr[84]) );
  GTECH_AND2 C4803 ( .A(N2515), .B(N2516), .Z(N2517) );
  GTECH_OR2 C4804 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[32]), .Z(N2515)
         );
  GTECH_OR2 C4805 ( .A(N2425), .B(a2stg_shr_tmp10[33]), .Z(N2516) );
  GTECH_NOT I_306 ( .A(N2520), .Z(a2stg_shr[83]) );
  GTECH_AND2 C4808 ( .A(N2518), .B(N2519), .Z(N2520) );
  GTECH_OR2 C4809 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[31]), .Z(N2518)
         );
  GTECH_OR2 C4810 ( .A(N2425), .B(a2stg_shr_tmp10[32]), .Z(N2519) );
  GTECH_NOT I_307 ( .A(N2523), .Z(a2stg_shr[82]) );
  GTECH_AND2 C4813 ( .A(N2521), .B(N2522), .Z(N2523) );
  GTECH_OR2 C4814 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[30]), .Z(N2521)
         );
  GTECH_OR2 C4815 ( .A(N2425), .B(a2stg_shr_tmp10[31]), .Z(N2522) );
  GTECH_NOT I_308 ( .A(N2526), .Z(a2stg_shr[81]) );
  GTECH_AND2 C4818 ( .A(N2524), .B(N2525), .Z(N2526) );
  GTECH_OR2 C4819 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[29]), .Z(N2524)
         );
  GTECH_OR2 C4820 ( .A(N2425), .B(a2stg_shr_tmp10[30]), .Z(N2525) );
  GTECH_NOT I_309 ( .A(N2529), .Z(a2stg_shr[80]) );
  GTECH_AND2 C4823 ( .A(N2527), .B(N2528), .Z(N2529) );
  GTECH_OR2 C4824 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[28]), .Z(N2527)
         );
  GTECH_OR2 C4825 ( .A(N2425), .B(a2stg_shr_tmp10[29]), .Z(N2528) );
  GTECH_NOT I_310 ( .A(N2532), .Z(a2stg_shr[79]) );
  GTECH_AND2 C4828 ( .A(N2530), .B(N2531), .Z(N2532) );
  GTECH_OR2 C4829 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[27]), .Z(N2530)
         );
  GTECH_OR2 C4830 ( .A(N2425), .B(a2stg_shr_tmp10[28]), .Z(N2531) );
  GTECH_NOT I_311 ( .A(N2535), .Z(a2stg_shr[78]) );
  GTECH_AND2 C4833 ( .A(N2533), .B(N2534), .Z(N2535) );
  GTECH_OR2 C4834 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[26]), .Z(N2533)
         );
  GTECH_OR2 C4835 ( .A(N2425), .B(a2stg_shr_tmp10[27]), .Z(N2534) );
  GTECH_NOT I_312 ( .A(N2538), .Z(a2stg_shr[77]) );
  GTECH_AND2 C4838 ( .A(N2536), .B(N2537), .Z(N2538) );
  GTECH_OR2 C4839 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[25]), .Z(N2536)
         );
  GTECH_OR2 C4840 ( .A(N2425), .B(a2stg_shr_tmp10[26]), .Z(N2537) );
  GTECH_NOT I_313 ( .A(N2541), .Z(a2stg_shr[76]) );
  GTECH_AND2 C4843 ( .A(N2539), .B(N2540), .Z(N2541) );
  GTECH_OR2 C4844 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[24]), .Z(N2539)
         );
  GTECH_OR2 C4845 ( .A(N2425), .B(a2stg_shr_tmp10[25]), .Z(N2540) );
  GTECH_NOT I_314 ( .A(N2544), .Z(a2stg_shr[75]) );
  GTECH_AND2 C4848 ( .A(N2542), .B(N2543), .Z(N2544) );
  GTECH_OR2 C4849 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[23]), .Z(N2542)
         );
  GTECH_OR2 C4850 ( .A(N2425), .B(a2stg_shr_tmp10[24]), .Z(N2543) );
  GTECH_NOT I_315 ( .A(N2547), .Z(a2stg_shr[74]) );
  GTECH_AND2 C4853 ( .A(N2545), .B(N2546), .Z(N2547) );
  GTECH_OR2 C4854 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[22]), .Z(N2545)
         );
  GTECH_OR2 C4855 ( .A(N2425), .B(a2stg_shr_tmp10[23]), .Z(N2546) );
  GTECH_NOT I_316 ( .A(N2550), .Z(a2stg_shr[73]) );
  GTECH_AND2 C4858 ( .A(N2548), .B(N2549), .Z(N2550) );
  GTECH_OR2 C4859 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[21]), .Z(N2548)
         );
  GTECH_OR2 C4860 ( .A(N2425), .B(a2stg_shr_tmp10[22]), .Z(N2549) );
  GTECH_NOT I_317 ( .A(N2553), .Z(a2stg_shr[72]) );
  GTECH_AND2 C4863 ( .A(N2551), .B(N2552), .Z(N2553) );
  GTECH_OR2 C4864 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[20]), .Z(N2551)
         );
  GTECH_OR2 C4865 ( .A(N2425), .B(a2stg_shr_tmp10[21]), .Z(N2552) );
  GTECH_NOT I_318 ( .A(N2556), .Z(a2stg_shr[71]) );
  GTECH_AND2 C4868 ( .A(N2554), .B(N2555), .Z(N2556) );
  GTECH_OR2 C4869 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[19]), .Z(N2554)
         );
  GTECH_OR2 C4870 ( .A(N2425), .B(a2stg_shr_tmp10[20]), .Z(N2555) );
  GTECH_NOT I_319 ( .A(N2559), .Z(a2stg_shr[70]) );
  GTECH_AND2 C4873 ( .A(N2557), .B(N2558), .Z(N2559) );
  GTECH_OR2 C4874 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[18]), .Z(N2557)
         );
  GTECH_OR2 C4875 ( .A(N2425), .B(a2stg_shr_tmp10[19]), .Z(N2558) );
  GTECH_NOT I_320 ( .A(N2562), .Z(a2stg_shr[69]) );
  GTECH_AND2 C4878 ( .A(N2560), .B(N2561), .Z(N2562) );
  GTECH_OR2 C4879 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[17]), .Z(N2560)
         );
  GTECH_OR2 C4880 ( .A(N2425), .B(a2stg_shr_tmp10[18]), .Z(N2561) );
  GTECH_NOT I_321 ( .A(N2565), .Z(a2stg_shr[68]) );
  GTECH_AND2 C4883 ( .A(N2563), .B(N2564), .Z(N2565) );
  GTECH_OR2 C4884 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[16]), .Z(N2563)
         );
  GTECH_OR2 C4885 ( .A(N2425), .B(a2stg_shr_tmp10[17]), .Z(N2564) );
  GTECH_NOT I_322 ( .A(N2568), .Z(a2stg_shr[67]) );
  GTECH_AND2 C4888 ( .A(N2566), .B(N2567), .Z(N2568) );
  GTECH_OR2 C4889 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[15]), .Z(N2566)
         );
  GTECH_OR2 C4890 ( .A(N2425), .B(a2stg_shr_tmp10[16]), .Z(N2567) );
  GTECH_NOT I_323 ( .A(N2571), .Z(a2stg_shr[66]) );
  GTECH_AND2 C4893 ( .A(N2569), .B(N2570), .Z(N2571) );
  GTECH_OR2 C4894 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[14]), .Z(N2569)
         );
  GTECH_OR2 C4895 ( .A(N2425), .B(a2stg_shr_tmp10[15]), .Z(N2570) );
  GTECH_NOT I_324 ( .A(N2574), .Z(a2stg_shr[65]) );
  GTECH_AND2 C4898 ( .A(N2572), .B(N2573), .Z(N2574) );
  GTECH_OR2 C4899 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[13]), .Z(N2572)
         );
  GTECH_OR2 C4900 ( .A(N2425), .B(a2stg_shr_tmp10[14]), .Z(N2573) );
  GTECH_NOT I_325 ( .A(N2577), .Z(a2stg_shr[64]) );
  GTECH_AND2 C4903 ( .A(N2575), .B(N2576), .Z(N2577) );
  GTECH_OR2 C4904 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[12]), .Z(N2575)
         );
  GTECH_OR2 C4905 ( .A(N2425), .B(a2stg_shr_tmp10[13]), .Z(N2576) );
  GTECH_NOT I_326 ( .A(N2580), .Z(a2stg_shr[63]) );
  GTECH_AND2 C4908 ( .A(N2578), .B(N2579), .Z(N2580) );
  GTECH_OR2 C4909 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[11]), .Z(N2578)
         );
  GTECH_OR2 C4910 ( .A(N2425), .B(a2stg_shr_tmp10[12]), .Z(N2579) );
  GTECH_NOT I_327 ( .A(N2583), .Z(a2stg_shr[62]) );
  GTECH_AND2 C4913 ( .A(N2581), .B(N2582), .Z(N2583) );
  GTECH_OR2 C4914 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[10]), .Z(N2581)
         );
  GTECH_OR2 C4915 ( .A(N2425), .B(a2stg_shr_tmp10[11]), .Z(N2582) );
  GTECH_NOT I_328 ( .A(N2586), .Z(a2stg_shr[61]) );
  GTECH_AND2 C4918 ( .A(N2584), .B(N2585), .Z(N2586) );
  GTECH_OR2 C4919 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[9]), .Z(N2584)
         );
  GTECH_OR2 C4920 ( .A(N2425), .B(a2stg_shr_tmp10[10]), .Z(N2585) );
  GTECH_NOT I_329 ( .A(N2589), .Z(a2stg_shr[60]) );
  GTECH_AND2 C4923 ( .A(N2587), .B(N2588), .Z(N2589) );
  GTECH_OR2 C4924 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[8]), .Z(N2587)
         );
  GTECH_OR2 C4925 ( .A(N2425), .B(a2stg_shr_tmp10[9]), .Z(N2588) );
  GTECH_NOT I_330 ( .A(N2592), .Z(a2stg_shr[59]) );
  GTECH_AND2 C4928 ( .A(N2590), .B(N2591), .Z(N2592) );
  GTECH_OR2 C4929 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[7]), .Z(N2590)
         );
  GTECH_OR2 C4930 ( .A(N2425), .B(a2stg_shr_tmp10[8]), .Z(N2591) );
  GTECH_NOT I_331 ( .A(N2595), .Z(a2stg_shr[58]) );
  GTECH_AND2 C4933 ( .A(N2593), .B(N2594), .Z(N2595) );
  GTECH_OR2 C4934 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[6]), .Z(N2593)
         );
  GTECH_OR2 C4935 ( .A(N2425), .B(a2stg_shr_tmp10[7]), .Z(N2594) );
  GTECH_NOT I_332 ( .A(N2598), .Z(a2stg_shr[57]) );
  GTECH_AND2 C4938 ( .A(N2596), .B(N2597), .Z(N2598) );
  GTECH_OR2 C4939 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[5]), .Z(N2596)
         );
  GTECH_OR2 C4940 ( .A(N2425), .B(a2stg_shr_tmp10[6]), .Z(N2597) );
  GTECH_NOT I_333 ( .A(N2601), .Z(a2stg_shr[56]) );
  GTECH_AND2 C4943 ( .A(N2599), .B(N2600), .Z(N2601) );
  GTECH_OR2 C4944 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[4]), .Z(N2599)
         );
  GTECH_OR2 C4945 ( .A(N2425), .B(a2stg_shr_tmp10[5]), .Z(N2600) );
  GTECH_NOT I_334 ( .A(N2604), .Z(a2stg_shr[55]) );
  GTECH_AND2 C4948 ( .A(N2602), .B(N2603), .Z(N2604) );
  GTECH_OR2 C4949 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[3]), .Z(N2602)
         );
  GTECH_OR2 C4950 ( .A(N2425), .B(a2stg_shr_tmp10[4]), .Z(N2603) );
  GTECH_NOT I_335 ( .A(N2607), .Z(a2stg_shr[54]) );
  GTECH_AND2 C4953 ( .A(N2605), .B(N2606), .Z(N2607) );
  GTECH_OR2 C4954 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[2]), .Z(N2605)
         );
  GTECH_OR2 C4955 ( .A(N2425), .B(a2stg_shr_tmp10[3]), .Z(N2606) );
  GTECH_NOT I_336 ( .A(N2610), .Z(a2stg_shr[53]) );
  GTECH_AND2 C4958 ( .A(N2608), .B(N2609), .Z(N2610) );
  GTECH_OR2 C4959 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[1]), .Z(N2608)
         );
  GTECH_OR2 C4960 ( .A(N2425), .B(a2stg_shr_tmp10[2]), .Z(N2609) );
  GTECH_NOT I_337 ( .A(N2613), .Z(a2stg_shr[52]) );
  GTECH_AND2 C4963 ( .A(N2611), .B(N2612), .Z(N2613) );
  GTECH_OR2 C4964 ( .A(a2stg_shr_cnt_0[0]), .B(a2stg_shr_tmp10[0]), .Z(N2611)
         );
  GTECH_OR2 C4965 ( .A(N2425), .B(a2stg_shr_tmp10[1]), .Z(N2612) );
  GTECH_NOT I_338 ( .A(a2stg_shr_tmp2[27]), .Z(a2stg_shr_tmp18[27]) );
  GTECH_NOT I_339 ( .A(a2stg_shr_tmp2[26]), .Z(a2stg_shr_tmp18[26]) );
  GTECH_NOT I_340 ( .A(a2stg_shr_tmp2[25]), .Z(a2stg_shr_tmp18[25]) );
  GTECH_NOT I_341 ( .A(a2stg_shr_tmp2[24]), .Z(a2stg_shr_tmp18[24]) );
  GTECH_NOT I_342 ( .A(a2stg_shr_tmp2[23]), .Z(a2stg_shr_tmp18[23]) );
  GTECH_NOT I_343 ( .A(a2stg_shr_tmp2[22]), .Z(a2stg_shr_tmp18[22]) );
  GTECH_NOT I_344 ( .A(a2stg_shr_tmp2[21]), .Z(a2stg_shr_tmp18[21]) );
  GTECH_NOT I_345 ( .A(a2stg_shr_tmp2[20]), .Z(a2stg_shr_tmp18[20]) );
  GTECH_NOT I_346 ( .A(a2stg_shr_tmp2[19]), .Z(a2stg_shr_tmp18[19]) );
  GTECH_NOT I_347 ( .A(a2stg_shr_tmp2[18]), .Z(a2stg_shr_tmp18[18]) );
  GTECH_NOT I_348 ( .A(a2stg_shr_tmp2[17]), .Z(a2stg_shr_tmp18[17]) );
  GTECH_NOT I_349 ( .A(a2stg_shr_tmp2[16]), .Z(a2stg_shr_tmp18[16]) );
  GTECH_NOT I_350 ( .A(a2stg_shr_tmp2[15]), .Z(a2stg_shr_tmp18[15]) );
  GTECH_NOT I_351 ( .A(a2stg_shr_tmp2[14]), .Z(a2stg_shr_tmp18[14]) );
  GTECH_NOT I_352 ( .A(a2stg_shr_tmp2[13]), .Z(a2stg_shr_tmp18[13]) );
  GTECH_NOT I_353 ( .A(a2stg_shr_tmp2[12]), .Z(a2stg_shr_tmp18[12]) );
  GTECH_OR2 C4983 ( .A(N2660), .B(a2stg_shr[83]), .Z(a2stg_fsdtoi_nx) );
  GTECH_OR2 C4984 ( .A(N2657), .B(N2659), .Z(N2660) );
  GTECH_OR2 C4985 ( .A(N2653), .B(N2656), .Z(N2657) );
  GTECH_OR2 C4986 ( .A(N2644), .B(N2652), .Z(N2653) );
  GTECH_OR2 C4987 ( .A(N2643), .B(a2stg_shr_tmp4[0]), .Z(N2644) );
  GTECH_OR2 C4988 ( .A(N2642), .B(a2stg_shr_tmp4[1]), .Z(N2643) );
  GTECH_OR2 C4989 ( .A(N2641), .B(a2stg_shr_tmp4[2]), .Z(N2642) );
  GTECH_OR2 C4990 ( .A(N2640), .B(a2stg_shr_tmp4[3]), .Z(N2641) );
  GTECH_OR2 C4991 ( .A(N2639), .B(a2stg_shr_tmp4[4]), .Z(N2640) );
  GTECH_OR2 C4992 ( .A(N2638), .B(a2stg_shr_tmp4[5]), .Z(N2639) );
  GTECH_OR2 C4993 ( .A(N2637), .B(a2stg_shr_tmp4[6]), .Z(N2638) );
  GTECH_OR2 C4994 ( .A(N2636), .B(a2stg_shr_tmp4[7]), .Z(N2637) );
  GTECH_OR2 C4995 ( .A(N2635), .B(a2stg_shr_tmp4[8]), .Z(N2636) );
  GTECH_OR2 C4996 ( .A(N2634), .B(a2stg_shr_tmp4[9]), .Z(N2635) );
  GTECH_OR2 C4997 ( .A(N2633), .B(a2stg_shr_tmp4[10]), .Z(N2634) );
  GTECH_OR2 C4998 ( .A(N2632), .B(a2stg_shr_tmp4[11]), .Z(N2633) );
  GTECH_OR2 C4999 ( .A(N2631), .B(a2stg_shr_tmp4[12]), .Z(N2632) );
  GTECH_OR2 C5000 ( .A(N2630), .B(a2stg_shr_tmp4[13]), .Z(N2631) );
  GTECH_OR2 C5001 ( .A(N2629), .B(a2stg_shr_tmp4[14]), .Z(N2630) );
  GTECH_OR2 C5002 ( .A(N2628), .B(a2stg_shr_tmp4[15]), .Z(N2629) );
  GTECH_OR2 C5003 ( .A(N2627), .B(a2stg_shr_tmp4[16]), .Z(N2628) );
  GTECH_OR2 C5004 ( .A(N2626), .B(a2stg_shr_tmp4[17]), .Z(N2627) );
  GTECH_OR2 C5005 ( .A(N2625), .B(a2stg_shr_tmp4[18]), .Z(N2626) );
  GTECH_OR2 C5006 ( .A(N2624), .B(a2stg_shr_tmp4[19]), .Z(N2625) );
  GTECH_OR2 C5007 ( .A(N2623), .B(a2stg_shr_tmp4[20]), .Z(N2624) );
  GTECH_OR2 C5008 ( .A(N2622), .B(a2stg_shr_tmp4[21]), .Z(N2623) );
  GTECH_OR2 C5009 ( .A(N2621), .B(a2stg_shr_tmp4[22]), .Z(N2622) );
  GTECH_OR2 C5010 ( .A(N2620), .B(a2stg_shr_tmp4[23]), .Z(N2621) );
  GTECH_OR2 C5011 ( .A(N2619), .B(a2stg_shr_tmp4[24]), .Z(N2620) );
  GTECH_OR2 C5012 ( .A(N2618), .B(a2stg_shr_tmp4[25]), .Z(N2619) );
  GTECH_OR2 C5013 ( .A(N2617), .B(a2stg_shr_tmp4[26]), .Z(N2618) );
  GTECH_OR2 C5014 ( .A(N2616), .B(a2stg_shr_tmp4[27]), .Z(N2617) );
  GTECH_OR2 C5015 ( .A(N2615), .B(a2stg_shr_tmp4[28]), .Z(N2616) );
  GTECH_OR2 C5016 ( .A(N2614), .B(a2stg_shr_tmp4[29]), .Z(N2615) );
  GTECH_OR2 C5017 ( .A(a2stg_shr_tmp4[31]), .B(a2stg_shr_tmp4[30]), .Z(N2614)
         );
  GTECH_NOT I_354 ( .A(N2651), .Z(N2652) );
  GTECH_AND2 C5019 ( .A(N2650), .B(a2stg_shr_tmp6[24]), .Z(N2651) );
  GTECH_AND2 C5020 ( .A(N2649), .B(a2stg_shr_tmp6[25]), .Z(N2650) );
  GTECH_AND2 C5021 ( .A(N2648), .B(a2stg_shr_tmp6[26]), .Z(N2649) );
  GTECH_AND2 C5022 ( .A(N2647), .B(a2stg_shr_tmp6[27]), .Z(N2648) );
  GTECH_AND2 C5023 ( .A(N2646), .B(a2stg_shr_tmp6[28]), .Z(N2647) );
  GTECH_AND2 C5024 ( .A(N2645), .B(a2stg_shr_tmp6[29]), .Z(N2646) );
  GTECH_AND2 C5025 ( .A(a2stg_shr_tmp6[31]), .B(a2stg_shr_tmp6[30]), .Z(N2645)
         );
  GTECH_OR2 C5026 ( .A(N2655), .B(a2stg_shr_tmp8[28]), .Z(N2656) );
  GTECH_OR2 C5027 ( .A(N2654), .B(a2stg_shr_tmp8[29]), .Z(N2655) );
  GTECH_OR2 C5028 ( .A(a2stg_shr_tmp8[31]), .B(a2stg_shr_tmp8[30]), .Z(N2654)
         );
  GTECH_NOT I_355 ( .A(N2658), .Z(N2659) );
  GTECH_AND2 C5030 ( .A(a2stg_shr_tmp10[31]), .B(a2stg_shr_tmp10[30]), .Z(
        N2658) );
  GTECH_NOT I_356 ( .A(N2664), .Z(a2stg_nx_neq0_84_tmp_1[63]) );
  GTECH_OR2 C5032 ( .A(N2661), .B(N2663), .Z(N2664) );
  GTECH_AND2 C5033 ( .A(a2stg_frac2a[43]), .B(a2stg_shr_cnt[5]), .Z(N2661) );
  GTECH_AND2 C5034 ( .A(a2stg_frac2a[11]), .B(N2662), .Z(N2663) );
  GTECH_NOT I_357 ( .A(a2stg_shr_cnt[5]), .Z(N2662) );
  GTECH_NOT I_358 ( .A(N2667), .Z(a2stg_nx_neq0_84_tmp_1[62]) );
  GTECH_OR2 C5037 ( .A(N2665), .B(N2666), .Z(N2667) );
  GTECH_AND2 C5038 ( .A(a2stg_frac2a[42]), .B(a2stg_shr_cnt[5]), .Z(N2665) );
  GTECH_AND2 C5039 ( .A(a2stg_frac2a[10]), .B(N2662), .Z(N2666) );
  GTECH_NOT I_359 ( .A(N2670), .Z(a2stg_nx_neq0_84_tmp_1[61]) );
  GTECH_OR2 C5042 ( .A(N2668), .B(N2669), .Z(N2670) );
  GTECH_AND2 C5043 ( .A(a2stg_frac2a[41]), .B(a2stg_shr_cnt[5]), .Z(N2668) );
  GTECH_AND2 C5044 ( .A(a2stg_frac2a[9]), .B(N2662), .Z(N2669) );
  GTECH_NOT I_360 ( .A(N2673), .Z(a2stg_nx_neq0_84_tmp_1[60]) );
  GTECH_OR2 C5047 ( .A(N2671), .B(N2672), .Z(N2673) );
  GTECH_AND2 C5048 ( .A(a2stg_frac2a[40]), .B(a2stg_shr_cnt[5]), .Z(N2671) );
  GTECH_AND2 C5049 ( .A(a2stg_frac2a[8]), .B(N2662), .Z(N2672) );
  GTECH_NOT I_361 ( .A(N2676), .Z(a2stg_nx_neq0_84_tmp_1[59]) );
  GTECH_OR2 C5052 ( .A(N2674), .B(N2675), .Z(N2676) );
  GTECH_AND2 C5053 ( .A(a2stg_frac2a[39]), .B(a2stg_shr_cnt[5]), .Z(N2674) );
  GTECH_AND2 C5054 ( .A(a2stg_frac2a[7]), .B(N2662), .Z(N2675) );
  GTECH_NOT I_362 ( .A(N2679), .Z(a2stg_nx_neq0_84_tmp_1[58]) );
  GTECH_OR2 C5057 ( .A(N2677), .B(N2678), .Z(N2679) );
  GTECH_AND2 C5058 ( .A(a2stg_frac2a[38]), .B(a2stg_shr_cnt[5]), .Z(N2677) );
  GTECH_AND2 C5059 ( .A(a2stg_frac2a[6]), .B(N2662), .Z(N2678) );
  GTECH_NOT I_363 ( .A(N2682), .Z(a2stg_nx_neq0_84_tmp_1[57]) );
  GTECH_OR2 C5062 ( .A(N2680), .B(N2681), .Z(N2682) );
  GTECH_AND2 C5063 ( .A(a2stg_frac2a[37]), .B(a2stg_shr_cnt[5]), .Z(N2680) );
  GTECH_AND2 C5064 ( .A(a2stg_frac2a[5]), .B(N2662), .Z(N2681) );
  GTECH_NOT I_364 ( .A(N2685), .Z(a2stg_nx_neq0_84_tmp_1[56]) );
  GTECH_OR2 C5067 ( .A(N2683), .B(N2684), .Z(N2685) );
  GTECH_AND2 C5068 ( .A(a2stg_frac2a[36]), .B(a2stg_shr_cnt[5]), .Z(N2683) );
  GTECH_AND2 C5069 ( .A(a2stg_frac2a[4]), .B(N2662), .Z(N2684) );
  GTECH_NOT I_365 ( .A(N2688), .Z(a2stg_nx_neq0_84_tmp_1[55]) );
  GTECH_OR2 C5072 ( .A(N2686), .B(N2687), .Z(N2688) );
  GTECH_AND2 C5073 ( .A(a2stg_frac2a[35]), .B(a2stg_shr_cnt[5]), .Z(N2686) );
  GTECH_AND2 C5074 ( .A(a2stg_frac2a[3]), .B(N2662), .Z(N2687) );
  GTECH_NOT I_366 ( .A(N2691), .Z(a2stg_nx_neq0_84_tmp_1[54]) );
  GTECH_OR2 C5077 ( .A(N2689), .B(N2690), .Z(N2691) );
  GTECH_AND2 C5078 ( .A(a2stg_frac2a[34]), .B(a2stg_shr_cnt[5]), .Z(N2689) );
  GTECH_AND2 C5079 ( .A(a2stg_frac2a[2]), .B(N2662), .Z(N2690) );
  GTECH_NOT I_367 ( .A(N2694), .Z(a2stg_nx_neq0_84_tmp_1[53]) );
  GTECH_OR2 C5082 ( .A(N2692), .B(N2693), .Z(N2694) );
  GTECH_AND2 C5083 ( .A(a2stg_frac2a[33]), .B(a2stg_shr_cnt[5]), .Z(N2692) );
  GTECH_AND2 C5084 ( .A(a2stg_frac2a[1]), .B(N2662), .Z(N2693) );
  GTECH_NOT I_368 ( .A(N2697), .Z(a2stg_nx_neq0_84_tmp_1[52]) );
  GTECH_OR2 C5087 ( .A(N2695), .B(N2696), .Z(N2697) );
  GTECH_AND2 C5088 ( .A(a2stg_frac2a[32]), .B(a2stg_shr_cnt[5]), .Z(N2695) );
  GTECH_AND2 C5089 ( .A(a2stg_frac2a[0]), .B(N2662), .Z(N2696) );
  GTECH_NOT I_369 ( .A(N2698), .Z(a2stg_nx_neq0_84_tmp_1[51]) );
  GTECH_AND2 C5092 ( .A(a2stg_frac2a[31]), .B(a2stg_shr_cnt[5]), .Z(N2698) );
  GTECH_NOT I_370 ( .A(N2699), .Z(a2stg_nx_neq0_84_tmp_1[50]) );
  GTECH_AND2 C5094 ( .A(a2stg_frac2a[30]), .B(a2stg_shr_cnt[5]), .Z(N2699) );
  GTECH_NOT I_371 ( .A(N2700), .Z(a2stg_nx_neq0_84_tmp_1[49]) );
  GTECH_AND2 C5096 ( .A(a2stg_frac2a[29]), .B(a2stg_shr_cnt[5]), .Z(N2700) );
  GTECH_NOT I_372 ( .A(N2701), .Z(a2stg_nx_neq0_84_tmp_1[48]) );
  GTECH_AND2 C5098 ( .A(a2stg_frac2a[28]), .B(a2stg_shr_cnt[5]), .Z(N2701) );
  GTECH_NOT I_373 ( .A(N2702), .Z(a2stg_nx_neq0_84_tmp_1[47]) );
  GTECH_AND2 C5100 ( .A(a2stg_frac2a[27]), .B(a2stg_shr_cnt[5]), .Z(N2702) );
  GTECH_NOT I_374 ( .A(N2703), .Z(a2stg_nx_neq0_84_tmp_1[46]) );
  GTECH_AND2 C5102 ( .A(a2stg_frac2a[26]), .B(a2stg_shr_cnt[5]), .Z(N2703) );
  GTECH_NOT I_375 ( .A(N2704), .Z(a2stg_nx_neq0_84_tmp_1[45]) );
  GTECH_AND2 C5104 ( .A(a2stg_frac2a[25]), .B(a2stg_shr_cnt[5]), .Z(N2704) );
  GTECH_NOT I_376 ( .A(N2705), .Z(a2stg_nx_neq0_84_tmp_1[44]) );
  GTECH_AND2 C5106 ( .A(a2stg_frac2a[24]), .B(a2stg_shr_cnt[5]), .Z(N2705) );
  GTECH_NOT I_377 ( .A(N2706), .Z(a2stg_nx_neq0_84_tmp_1[43]) );
  GTECH_AND2 C5108 ( .A(a2stg_frac2a[23]), .B(a2stg_shr_cnt[5]), .Z(N2706) );
  GTECH_NOT I_378 ( .A(N2707), .Z(a2stg_nx_neq0_84_tmp_1[42]) );
  GTECH_AND2 C5110 ( .A(a2stg_frac2a[22]), .B(a2stg_shr_cnt[5]), .Z(N2707) );
  GTECH_NOT I_379 ( .A(N2708), .Z(a2stg_nx_neq0_84_tmp_1[41]) );
  GTECH_AND2 C5112 ( .A(a2stg_frac2a[21]), .B(a2stg_shr_cnt[5]), .Z(N2708) );
  GTECH_NOT I_380 ( .A(N2709), .Z(a2stg_nx_neq0_84_tmp_1[40]) );
  GTECH_AND2 C5114 ( .A(a2stg_frac2a[20]), .B(a2stg_shr_cnt[5]), .Z(N2709) );
  GTECH_NOT I_381 ( .A(N2710), .Z(a2stg_nx_neq0_84_tmp_1[39]) );
  GTECH_AND2 C5116 ( .A(a2stg_frac2a[19]), .B(a2stg_shr_cnt[5]), .Z(N2710) );
  GTECH_NOT I_382 ( .A(N2711), .Z(a2stg_nx_neq0_84_tmp_1[38]) );
  GTECH_AND2 C5118 ( .A(a2stg_frac2a[18]), .B(a2stg_shr_cnt[5]), .Z(N2711) );
  GTECH_NOT I_383 ( .A(N2712), .Z(a2stg_nx_neq0_84_tmp_1[37]) );
  GTECH_AND2 C5120 ( .A(a2stg_frac2a[17]), .B(a2stg_shr_cnt[5]), .Z(N2712) );
  GTECH_NOT I_384 ( .A(N2713), .Z(a2stg_nx_neq0_84_tmp_1[36]) );
  GTECH_AND2 C5122 ( .A(a2stg_frac2a[16]), .B(a2stg_shr_cnt[5]), .Z(N2713) );
  GTECH_NOT I_385 ( .A(N2714), .Z(a2stg_nx_neq0_84_tmp_1[35]) );
  GTECH_AND2 C5124 ( .A(a2stg_frac2a[15]), .B(a2stg_shr_cnt[5]), .Z(N2714) );
  GTECH_NOT I_386 ( .A(N2715), .Z(a2stg_nx_neq0_84_tmp_1[34]) );
  GTECH_AND2 C5126 ( .A(a2stg_frac2a[14]), .B(a2stg_shr_cnt[5]), .Z(N2715) );
  GTECH_NOT I_387 ( .A(N2716), .Z(a2stg_nx_neq0_84_tmp_1[33]) );
  GTECH_AND2 C5128 ( .A(a2stg_frac2a[13]), .B(a2stg_shr_cnt[5]), .Z(N2716) );
  GTECH_NOT I_388 ( .A(N2717), .Z(a2stg_nx_neq0_84_tmp_1[32]) );
  GTECH_AND2 C5130 ( .A(a2stg_frac2a[12]), .B(a2stg_shr_cnt[5]), .Z(N2717) );
  GTECH_NOT I_389 ( .A(N2718), .Z(a2stg_nx_neq0_84_tmp_1[31]) );
  GTECH_AND2 C5132 ( .A(a2stg_frac2a[11]), .B(a2stg_shr_cnt[5]), .Z(N2718) );
  GTECH_NOT I_390 ( .A(N2719), .Z(a2stg_nx_neq0_84_tmp_1[30]) );
  GTECH_AND2 C5134 ( .A(a2stg_frac2a[10]), .B(a2stg_shr_cnt[5]), .Z(N2719) );
  GTECH_NOT I_391 ( .A(N2720), .Z(a2stg_nx_neq0_84_tmp_1[29]) );
  GTECH_AND2 C5136 ( .A(a2stg_frac2a[9]), .B(a2stg_shr_cnt[5]), .Z(N2720) );
  GTECH_NOT I_392 ( .A(N2721), .Z(a2stg_nx_neq0_84_tmp_1[28]) );
  GTECH_AND2 C5138 ( .A(a2stg_frac2a[8]), .B(a2stg_shr_cnt[5]), .Z(N2721) );
  GTECH_NOT I_393 ( .A(N2722), .Z(a2stg_nx_neq0_84_tmp_1[27]) );
  GTECH_AND2 C5140 ( .A(a2stg_frac2a[7]), .B(a2stg_shr_cnt[5]), .Z(N2722) );
  GTECH_NOT I_394 ( .A(N2723), .Z(a2stg_nx_neq0_84_tmp_1[26]) );
  GTECH_AND2 C5142 ( .A(a2stg_frac2a[6]), .B(a2stg_shr_cnt[5]), .Z(N2723) );
  GTECH_NOT I_395 ( .A(N2724), .Z(a2stg_nx_neq0_84_tmp_1[25]) );
  GTECH_AND2 C5144 ( .A(a2stg_frac2a[5]), .B(a2stg_shr_cnt[5]), .Z(N2724) );
  GTECH_NOT I_396 ( .A(N2725), .Z(a2stg_nx_neq0_84_tmp_1[24]) );
  GTECH_AND2 C5146 ( .A(a2stg_frac2a[4]), .B(a2stg_shr_cnt[5]), .Z(N2725) );
  GTECH_NOT I_397 ( .A(N2726), .Z(a2stg_nx_neq0_84_tmp_1[23]) );
  GTECH_AND2 C5148 ( .A(a2stg_frac2a[3]), .B(a2stg_shr_cnt[5]), .Z(N2726) );
  GTECH_NOT I_398 ( .A(N2727), .Z(a2stg_nx_neq0_84_tmp_1[22]) );
  GTECH_AND2 C5150 ( .A(a2stg_frac2a[2]), .B(a2stg_shr_cnt[5]), .Z(N2727) );
  GTECH_NOT I_399 ( .A(N2728), .Z(a2stg_nx_neq0_84_tmp_1[21]) );
  GTECH_AND2 C5152 ( .A(a2stg_frac2a[1]), .B(a2stg_shr_cnt[5]), .Z(N2728) );
  GTECH_NOT I_400 ( .A(N2729), .Z(a2stg_nx_neq0_84_tmp_1[20]) );
  GTECH_AND2 C5154 ( .A(a2stg_frac2a[0]), .B(a2stg_shr_cnt[5]), .Z(N2729) );
  GTECH_NOT I_401 ( .A(N2733), .Z(a2stg_nx_neq0_84_tmp_2[63]) );
  GTECH_AND2 C5156 ( .A(N2731), .B(N2732), .Z(N2733) );
  GTECH_OR2 C5157 ( .A(a2stg_shr_tmp18[27]), .B(N2730), .Z(N2731) );
  GTECH_NOT I_402 ( .A(a2stg_shr_cnt[4]), .Z(N2730) );
  GTECH_OR2 C5159 ( .A(a2stg_nx_neq0_84_tmp_1[63]), .B(a2stg_shr_cnt[4]), .Z(
        N2732) );
  GTECH_NOT I_403 ( .A(N2736), .Z(a2stg_nx_neq0_84_tmp_2[62]) );
  GTECH_AND2 C5161 ( .A(N2734), .B(N2735), .Z(N2736) );
  GTECH_OR2 C5162 ( .A(a2stg_shr_tmp18[26]), .B(N2730), .Z(N2734) );
  GTECH_OR2 C5164 ( .A(a2stg_nx_neq0_84_tmp_1[62]), .B(a2stg_shr_cnt[4]), .Z(
        N2735) );
  GTECH_NOT I_404 ( .A(N2739), .Z(a2stg_nx_neq0_84_tmp_2[61]) );
  GTECH_AND2 C5166 ( .A(N2737), .B(N2738), .Z(N2739) );
  GTECH_OR2 C5167 ( .A(a2stg_shr_tmp18[25]), .B(N2730), .Z(N2737) );
  GTECH_OR2 C5169 ( .A(a2stg_nx_neq0_84_tmp_1[61]), .B(a2stg_shr_cnt[4]), .Z(
        N2738) );
  GTECH_NOT I_405 ( .A(N2742), .Z(a2stg_nx_neq0_84_tmp_2[60]) );
  GTECH_AND2 C5171 ( .A(N2740), .B(N2741), .Z(N2742) );
  GTECH_OR2 C5172 ( .A(a2stg_shr_tmp18[24]), .B(N2730), .Z(N2740) );
  GTECH_OR2 C5174 ( .A(a2stg_nx_neq0_84_tmp_1[60]), .B(a2stg_shr_cnt[4]), .Z(
        N2741) );
  GTECH_NOT I_406 ( .A(N2745), .Z(a2stg_nx_neq0_84_tmp_2[59]) );
  GTECH_AND2 C5176 ( .A(N2743), .B(N2744), .Z(N2745) );
  GTECH_OR2 C5177 ( .A(a2stg_shr_tmp18[23]), .B(N2730), .Z(N2743) );
  GTECH_OR2 C5179 ( .A(a2stg_nx_neq0_84_tmp_1[59]), .B(a2stg_shr_cnt[4]), .Z(
        N2744) );
  GTECH_NOT I_407 ( .A(N2748), .Z(a2stg_nx_neq0_84_tmp_2[58]) );
  GTECH_AND2 C5181 ( .A(N2746), .B(N2747), .Z(N2748) );
  GTECH_OR2 C5182 ( .A(a2stg_shr_tmp18[22]), .B(N2730), .Z(N2746) );
  GTECH_OR2 C5184 ( .A(a2stg_nx_neq0_84_tmp_1[58]), .B(a2stg_shr_cnt[4]), .Z(
        N2747) );
  GTECH_NOT I_408 ( .A(N2751), .Z(a2stg_nx_neq0_84_tmp_2[57]) );
  GTECH_AND2 C5186 ( .A(N2749), .B(N2750), .Z(N2751) );
  GTECH_OR2 C5187 ( .A(a2stg_shr_tmp18[21]), .B(N2730), .Z(N2749) );
  GTECH_OR2 C5189 ( .A(a2stg_nx_neq0_84_tmp_1[57]), .B(a2stg_shr_cnt[4]), .Z(
        N2750) );
  GTECH_NOT I_409 ( .A(N2754), .Z(a2stg_nx_neq0_84_tmp_2[56]) );
  GTECH_AND2 C5191 ( .A(N2752), .B(N2753), .Z(N2754) );
  GTECH_OR2 C5192 ( .A(a2stg_shr_tmp18[20]), .B(N2730), .Z(N2752) );
  GTECH_OR2 C5194 ( .A(a2stg_nx_neq0_84_tmp_1[56]), .B(a2stg_shr_cnt[4]), .Z(
        N2753) );
  GTECH_NOT I_410 ( .A(N2757), .Z(a2stg_nx_neq0_84_tmp_2[55]) );
  GTECH_AND2 C5196 ( .A(N2755), .B(N2756), .Z(N2757) );
  GTECH_OR2 C5197 ( .A(a2stg_shr_tmp18[19]), .B(N2730), .Z(N2755) );
  GTECH_OR2 C5199 ( .A(a2stg_nx_neq0_84_tmp_1[55]), .B(a2stg_shr_cnt[4]), .Z(
        N2756) );
  GTECH_NOT I_411 ( .A(N2760), .Z(a2stg_nx_neq0_84_tmp_2[54]) );
  GTECH_AND2 C5201 ( .A(N2758), .B(N2759), .Z(N2760) );
  GTECH_OR2 C5202 ( .A(a2stg_shr_tmp18[18]), .B(N2730), .Z(N2758) );
  GTECH_OR2 C5204 ( .A(a2stg_nx_neq0_84_tmp_1[54]), .B(a2stg_shr_cnt[4]), .Z(
        N2759) );
  GTECH_NOT I_412 ( .A(N2763), .Z(a2stg_nx_neq0_84_tmp_2[53]) );
  GTECH_AND2 C5206 ( .A(N2761), .B(N2762), .Z(N2763) );
  GTECH_OR2 C5207 ( .A(a2stg_shr_tmp18[17]), .B(N2730), .Z(N2761) );
  GTECH_OR2 C5209 ( .A(a2stg_nx_neq0_84_tmp_1[53]), .B(a2stg_shr_cnt[4]), .Z(
        N2762) );
  GTECH_NOT I_413 ( .A(N2766), .Z(a2stg_nx_neq0_84_tmp_2[52]) );
  GTECH_AND2 C5211 ( .A(N2764), .B(N2765), .Z(N2766) );
  GTECH_OR2 C5212 ( .A(a2stg_shr_tmp18[16]), .B(N2730), .Z(N2764) );
  GTECH_OR2 C5214 ( .A(a2stg_nx_neq0_84_tmp_1[52]), .B(a2stg_shr_cnt[4]), .Z(
        N2765) );
  GTECH_NOT I_414 ( .A(N2769), .Z(a2stg_nx_neq0_84_tmp_2[51]) );
  GTECH_AND2 C5216 ( .A(N2767), .B(N2768), .Z(N2769) );
  GTECH_OR2 C5217 ( .A(a2stg_shr_tmp18[15]), .B(N2730), .Z(N2767) );
  GTECH_OR2 C5219 ( .A(a2stg_nx_neq0_84_tmp_1[51]), .B(a2stg_shr_cnt[4]), .Z(
        N2768) );
  GTECH_NOT I_415 ( .A(N2772), .Z(a2stg_nx_neq0_84_tmp_2[50]) );
  GTECH_AND2 C5221 ( .A(N2770), .B(N2771), .Z(N2772) );
  GTECH_OR2 C5222 ( .A(a2stg_shr_tmp18[14]), .B(N2730), .Z(N2770) );
  GTECH_OR2 C5224 ( .A(a2stg_nx_neq0_84_tmp_1[50]), .B(a2stg_shr_cnt[4]), .Z(
        N2771) );
  GTECH_NOT I_416 ( .A(N2775), .Z(a2stg_nx_neq0_84_tmp_2[49]) );
  GTECH_AND2 C5226 ( .A(N2773), .B(N2774), .Z(N2775) );
  GTECH_OR2 C5227 ( .A(a2stg_shr_tmp18[13]), .B(N2730), .Z(N2773) );
  GTECH_OR2 C5229 ( .A(a2stg_nx_neq0_84_tmp_1[49]), .B(a2stg_shr_cnt[4]), .Z(
        N2774) );
  GTECH_NOT I_417 ( .A(N2778), .Z(a2stg_nx_neq0_84_tmp_2[48]) );
  GTECH_AND2 C5231 ( .A(N2776), .B(N2777), .Z(N2778) );
  GTECH_OR2 C5232 ( .A(a2stg_shr_tmp18[12]), .B(N2730), .Z(N2776) );
  GTECH_OR2 C5234 ( .A(a2stg_nx_neq0_84_tmp_1[48]), .B(a2stg_shr_cnt[4]), .Z(
        N2777) );
  GTECH_NOT I_418 ( .A(N2781), .Z(a2stg_nx_neq0_84_tmp_2[47]) );
  GTECH_AND2 C5236 ( .A(N2779), .B(N2780), .Z(N2781) );
  GTECH_OR2 C5237 ( .A(a2stg_nx_neq0_84_tmp_1[63]), .B(N2730), .Z(N2779) );
  GTECH_OR2 C5239 ( .A(a2stg_nx_neq0_84_tmp_1[47]), .B(a2stg_shr_cnt[4]), .Z(
        N2780) );
  GTECH_NOT I_419 ( .A(N2784), .Z(a2stg_nx_neq0_84_tmp_2[46]) );
  GTECH_AND2 C5241 ( .A(N2782), .B(N2783), .Z(N2784) );
  GTECH_OR2 C5242 ( .A(a2stg_nx_neq0_84_tmp_1[62]), .B(N2730), .Z(N2782) );
  GTECH_OR2 C5244 ( .A(a2stg_nx_neq0_84_tmp_1[46]), .B(a2stg_shr_cnt[4]), .Z(
        N2783) );
  GTECH_NOT I_420 ( .A(N2787), .Z(a2stg_nx_neq0_84_tmp_2[45]) );
  GTECH_AND2 C5246 ( .A(N2785), .B(N2786), .Z(N2787) );
  GTECH_OR2 C5247 ( .A(a2stg_nx_neq0_84_tmp_1[61]), .B(N2730), .Z(N2785) );
  GTECH_OR2 C5249 ( .A(a2stg_nx_neq0_84_tmp_1[45]), .B(a2stg_shr_cnt[4]), .Z(
        N2786) );
  GTECH_NOT I_421 ( .A(N2790), .Z(a2stg_nx_neq0_84_tmp_2[44]) );
  GTECH_AND2 C5251 ( .A(N2788), .B(N2789), .Z(N2790) );
  GTECH_OR2 C5252 ( .A(a2stg_nx_neq0_84_tmp_1[60]), .B(N2730), .Z(N2788) );
  GTECH_OR2 C5254 ( .A(a2stg_nx_neq0_84_tmp_1[44]), .B(a2stg_shr_cnt[4]), .Z(
        N2789) );
  GTECH_NOT I_422 ( .A(N2793), .Z(a2stg_nx_neq0_84_tmp_2[43]) );
  GTECH_AND2 C5256 ( .A(N2791), .B(N2792), .Z(N2793) );
  GTECH_OR2 C5257 ( .A(a2stg_nx_neq0_84_tmp_1[59]), .B(N2730), .Z(N2791) );
  GTECH_OR2 C5259 ( .A(a2stg_nx_neq0_84_tmp_1[43]), .B(a2stg_shr_cnt[4]), .Z(
        N2792) );
  GTECH_NOT I_423 ( .A(N2796), .Z(a2stg_nx_neq0_84_tmp_2[42]) );
  GTECH_AND2 C5261 ( .A(N2794), .B(N2795), .Z(N2796) );
  GTECH_OR2 C5262 ( .A(a2stg_nx_neq0_84_tmp_1[58]), .B(N2730), .Z(N2794) );
  GTECH_OR2 C5264 ( .A(a2stg_nx_neq0_84_tmp_1[42]), .B(a2stg_shr_cnt[4]), .Z(
        N2795) );
  GTECH_NOT I_424 ( .A(N2799), .Z(a2stg_nx_neq0_84_tmp_2[41]) );
  GTECH_AND2 C5266 ( .A(N2797), .B(N2798), .Z(N2799) );
  GTECH_OR2 C5267 ( .A(a2stg_nx_neq0_84_tmp_1[57]), .B(N2730), .Z(N2797) );
  GTECH_OR2 C5269 ( .A(a2stg_nx_neq0_84_tmp_1[41]), .B(a2stg_shr_cnt[4]), .Z(
        N2798) );
  GTECH_NOT I_425 ( .A(N2802), .Z(a2stg_nx_neq0_84_tmp_2[40]) );
  GTECH_AND2 C5271 ( .A(N2800), .B(N2801), .Z(N2802) );
  GTECH_OR2 C5272 ( .A(a2stg_nx_neq0_84_tmp_1[56]), .B(N2730), .Z(N2800) );
  GTECH_OR2 C5274 ( .A(a2stg_nx_neq0_84_tmp_1[40]), .B(a2stg_shr_cnt[4]), .Z(
        N2801) );
  GTECH_NOT I_426 ( .A(N2805), .Z(a2stg_nx_neq0_84_tmp_2[39]) );
  GTECH_AND2 C5276 ( .A(N2803), .B(N2804), .Z(N2805) );
  GTECH_OR2 C5277 ( .A(a2stg_nx_neq0_84_tmp_1[55]), .B(N2730), .Z(N2803) );
  GTECH_OR2 C5279 ( .A(a2stg_nx_neq0_84_tmp_1[39]), .B(a2stg_shr_cnt[4]), .Z(
        N2804) );
  GTECH_NOT I_427 ( .A(N2808), .Z(a2stg_nx_neq0_84_tmp_2[38]) );
  GTECH_AND2 C5281 ( .A(N2806), .B(N2807), .Z(N2808) );
  GTECH_OR2 C5282 ( .A(a2stg_nx_neq0_84_tmp_1[54]), .B(N2730), .Z(N2806) );
  GTECH_OR2 C5284 ( .A(a2stg_nx_neq0_84_tmp_1[38]), .B(a2stg_shr_cnt[4]), .Z(
        N2807) );
  GTECH_NOT I_428 ( .A(N2811), .Z(a2stg_nx_neq0_84_tmp_2[37]) );
  GTECH_AND2 C5286 ( .A(N2809), .B(N2810), .Z(N2811) );
  GTECH_OR2 C5287 ( .A(a2stg_nx_neq0_84_tmp_1[53]), .B(N2730), .Z(N2809) );
  GTECH_OR2 C5289 ( .A(a2stg_nx_neq0_84_tmp_1[37]), .B(a2stg_shr_cnt[4]), .Z(
        N2810) );
  GTECH_NOT I_429 ( .A(N2814), .Z(a2stg_nx_neq0_84_tmp_2[36]) );
  GTECH_AND2 C5291 ( .A(N2812), .B(N2813), .Z(N2814) );
  GTECH_OR2 C5292 ( .A(a2stg_nx_neq0_84_tmp_1[52]), .B(N2730), .Z(N2812) );
  GTECH_OR2 C5294 ( .A(a2stg_nx_neq0_84_tmp_1[36]), .B(a2stg_shr_cnt[4]), .Z(
        N2813) );
  GTECH_NOT I_430 ( .A(N2818), .Z(a2stg_nx_neq0_84_tmp_3[63]) );
  GTECH_OR2 C5296 ( .A(N2815), .B(N2817), .Z(N2818) );
  GTECH_AND2 C5297 ( .A(a2stg_shr_tmp4[19]), .B(a2stg_shr_cnt[3]), .Z(N2815)
         );
  GTECH_AND2 C5298 ( .A(a2stg_nx_neq0_84_tmp_2[63]), .B(N2816), .Z(N2817) );
  GTECH_NOT I_431 ( .A(a2stg_shr_cnt[3]), .Z(N2816) );
  GTECH_NOT I_432 ( .A(N2821), .Z(a2stg_nx_neq0_84_tmp_3[62]) );
  GTECH_OR2 C5301 ( .A(N2819), .B(N2820), .Z(N2821) );
  GTECH_AND2 C5302 ( .A(a2stg_shr_tmp4[18]), .B(a2stg_shr_cnt[3]), .Z(N2819)
         );
  GTECH_AND2 C5303 ( .A(a2stg_nx_neq0_84_tmp_2[62]), .B(N2816), .Z(N2820) );
  GTECH_NOT I_433 ( .A(N2824), .Z(a2stg_nx_neq0_84_tmp_3[61]) );
  GTECH_OR2 C5306 ( .A(N2822), .B(N2823), .Z(N2824) );
  GTECH_AND2 C5307 ( .A(a2stg_shr_tmp4[17]), .B(a2stg_shr_cnt[3]), .Z(N2822)
         );
  GTECH_AND2 C5308 ( .A(a2stg_nx_neq0_84_tmp_2[61]), .B(N2816), .Z(N2823) );
  GTECH_NOT I_434 ( .A(N2827), .Z(a2stg_nx_neq0_84_tmp_3[60]) );
  GTECH_OR2 C5311 ( .A(N2825), .B(N2826), .Z(N2827) );
  GTECH_AND2 C5312 ( .A(a2stg_shr_tmp4[16]), .B(a2stg_shr_cnt[3]), .Z(N2825)
         );
  GTECH_AND2 C5313 ( .A(a2stg_nx_neq0_84_tmp_2[60]), .B(N2816), .Z(N2826) );
  GTECH_NOT I_435 ( .A(N2830), .Z(a2stg_nx_neq0_84_tmp_3[59]) );
  GTECH_OR2 C5316 ( .A(N2828), .B(N2829), .Z(N2830) );
  GTECH_AND2 C5317 ( .A(a2stg_shr_tmp4[15]), .B(a2stg_shr_cnt[3]), .Z(N2828)
         );
  GTECH_AND2 C5318 ( .A(a2stg_nx_neq0_84_tmp_2[59]), .B(N2816), .Z(N2829) );
  GTECH_NOT I_436 ( .A(N2833), .Z(a2stg_nx_neq0_84_tmp_3[58]) );
  GTECH_OR2 C5321 ( .A(N2831), .B(N2832), .Z(N2833) );
  GTECH_AND2 C5322 ( .A(a2stg_shr_tmp4[14]), .B(a2stg_shr_cnt[3]), .Z(N2831)
         );
  GTECH_AND2 C5323 ( .A(a2stg_nx_neq0_84_tmp_2[58]), .B(N2816), .Z(N2832) );
  GTECH_NOT I_437 ( .A(N2836), .Z(a2stg_nx_neq0_84_tmp_3[57]) );
  GTECH_OR2 C5326 ( .A(N2834), .B(N2835), .Z(N2836) );
  GTECH_AND2 C5327 ( .A(a2stg_shr_tmp4[13]), .B(a2stg_shr_cnt[3]), .Z(N2834)
         );
  GTECH_AND2 C5328 ( .A(a2stg_nx_neq0_84_tmp_2[57]), .B(N2816), .Z(N2835) );
  GTECH_NOT I_438 ( .A(N2839), .Z(a2stg_nx_neq0_84_tmp_3[56]) );
  GTECH_OR2 C5331 ( .A(N2837), .B(N2838), .Z(N2839) );
  GTECH_AND2 C5332 ( .A(a2stg_shr_tmp4[12]), .B(a2stg_shr_cnt[3]), .Z(N2837)
         );
  GTECH_AND2 C5333 ( .A(a2stg_nx_neq0_84_tmp_2[56]), .B(N2816), .Z(N2838) );
  GTECH_NOT I_439 ( .A(N2842), .Z(a2stg_nx_neq0_84_tmp_3[55]) );
  GTECH_OR2 C5336 ( .A(N2840), .B(N2841), .Z(N2842) );
  GTECH_AND2 C5337 ( .A(a2stg_nx_neq0_84_tmp_2[63]), .B(a2stg_shr_cnt[3]), .Z(
        N2840) );
  GTECH_AND2 C5338 ( .A(a2stg_nx_neq0_84_tmp_2[55]), .B(N2816), .Z(N2841) );
  GTECH_NOT I_440 ( .A(N2845), .Z(a2stg_nx_neq0_84_tmp_3[54]) );
  GTECH_OR2 C5341 ( .A(N2843), .B(N2844), .Z(N2845) );
  GTECH_AND2 C5342 ( .A(a2stg_nx_neq0_84_tmp_2[62]), .B(a2stg_shr_cnt[3]), .Z(
        N2843) );
  GTECH_AND2 C5343 ( .A(a2stg_nx_neq0_84_tmp_2[54]), .B(N2816), .Z(N2844) );
  GTECH_NOT I_441 ( .A(N2848), .Z(a2stg_nx_neq0_84_tmp_3[53]) );
  GTECH_OR2 C5346 ( .A(N2846), .B(N2847), .Z(N2848) );
  GTECH_AND2 C5347 ( .A(a2stg_nx_neq0_84_tmp_2[61]), .B(a2stg_shr_cnt[3]), .Z(
        N2846) );
  GTECH_AND2 C5348 ( .A(a2stg_nx_neq0_84_tmp_2[53]), .B(N2816), .Z(N2847) );
  GTECH_NOT I_442 ( .A(N2851), .Z(a2stg_nx_neq0_84_tmp_3[52]) );
  GTECH_OR2 C5351 ( .A(N2849), .B(N2850), .Z(N2851) );
  GTECH_AND2 C5352 ( .A(a2stg_nx_neq0_84_tmp_2[60]), .B(a2stg_shr_cnt[3]), .Z(
        N2849) );
  GTECH_AND2 C5353 ( .A(a2stg_nx_neq0_84_tmp_2[52]), .B(N2816), .Z(N2850) );
  GTECH_NOT I_443 ( .A(N2854), .Z(a2stg_nx_neq0_84_tmp_3[51]) );
  GTECH_OR2 C5356 ( .A(N2852), .B(N2853), .Z(N2854) );
  GTECH_AND2 C5357 ( .A(a2stg_nx_neq0_84_tmp_2[59]), .B(a2stg_shr_cnt[3]), .Z(
        N2852) );
  GTECH_AND2 C5358 ( .A(a2stg_nx_neq0_84_tmp_2[51]), .B(N2816), .Z(N2853) );
  GTECH_NOT I_444 ( .A(N2857), .Z(a2stg_nx_neq0_84_tmp_3[50]) );
  GTECH_OR2 C5361 ( .A(N2855), .B(N2856), .Z(N2857) );
  GTECH_AND2 C5362 ( .A(a2stg_nx_neq0_84_tmp_2[58]), .B(a2stg_shr_cnt[3]), .Z(
        N2855) );
  GTECH_AND2 C5363 ( .A(a2stg_nx_neq0_84_tmp_2[50]), .B(N2816), .Z(N2856) );
  GTECH_NOT I_445 ( .A(N2860), .Z(a2stg_nx_neq0_84_tmp_3[49]) );
  GTECH_OR2 C5366 ( .A(N2858), .B(N2859), .Z(N2860) );
  GTECH_AND2 C5367 ( .A(a2stg_nx_neq0_84_tmp_2[57]), .B(a2stg_shr_cnt[3]), .Z(
        N2858) );
  GTECH_AND2 C5368 ( .A(a2stg_nx_neq0_84_tmp_2[49]), .B(N2816), .Z(N2859) );
  GTECH_NOT I_446 ( .A(N2863), .Z(a2stg_nx_neq0_84_tmp_3[48]) );
  GTECH_OR2 C5371 ( .A(N2861), .B(N2862), .Z(N2863) );
  GTECH_AND2 C5372 ( .A(a2stg_nx_neq0_84_tmp_2[56]), .B(a2stg_shr_cnt[3]), .Z(
        N2861) );
  GTECH_AND2 C5373 ( .A(a2stg_nx_neq0_84_tmp_2[48]), .B(N2816), .Z(N2862) );
  GTECH_NOT I_447 ( .A(N2866), .Z(a2stg_nx_neq0_84_tmp_3[47]) );
  GTECH_OR2 C5376 ( .A(N2864), .B(N2865), .Z(N2866) );
  GTECH_AND2 C5377 ( .A(a2stg_nx_neq0_84_tmp_2[55]), .B(a2stg_shr_cnt[3]), .Z(
        N2864) );
  GTECH_AND2 C5378 ( .A(a2stg_nx_neq0_84_tmp_2[47]), .B(N2816), .Z(N2865) );
  GTECH_NOT I_448 ( .A(N2869), .Z(a2stg_nx_neq0_84_tmp_3[46]) );
  GTECH_OR2 C5381 ( .A(N2867), .B(N2868), .Z(N2869) );
  GTECH_AND2 C5382 ( .A(a2stg_nx_neq0_84_tmp_2[54]), .B(a2stg_shr_cnt[3]), .Z(
        N2867) );
  GTECH_AND2 C5383 ( .A(a2stg_nx_neq0_84_tmp_2[46]), .B(N2816), .Z(N2868) );
  GTECH_NOT I_449 ( .A(N2872), .Z(a2stg_nx_neq0_84_tmp_3[45]) );
  GTECH_OR2 C5386 ( .A(N2870), .B(N2871), .Z(N2872) );
  GTECH_AND2 C5387 ( .A(a2stg_nx_neq0_84_tmp_2[53]), .B(a2stg_shr_cnt[3]), .Z(
        N2870) );
  GTECH_AND2 C5388 ( .A(a2stg_nx_neq0_84_tmp_2[45]), .B(N2816), .Z(N2871) );
  GTECH_NOT I_450 ( .A(N2875), .Z(a2stg_nx_neq0_84_tmp_3[44]) );
  GTECH_OR2 C5391 ( .A(N2873), .B(N2874), .Z(N2875) );
  GTECH_AND2 C5392 ( .A(a2stg_nx_neq0_84_tmp_2[52]), .B(a2stg_shr_cnt[3]), .Z(
        N2873) );
  GTECH_AND2 C5393 ( .A(a2stg_nx_neq0_84_tmp_2[44]), .B(N2816), .Z(N2874) );
  GTECH_NOT I_451 ( .A(N2879), .Z(a2stg_nx_neq0_84_tmp_4[63]) );
  GTECH_AND2 C5396 ( .A(N2877), .B(N2878), .Z(N2879) );
  GTECH_OR2 C5397 ( .A(a2stg_shr_tmp6[15]), .B(N2876), .Z(N2877) );
  GTECH_NOT I_452 ( .A(a2stg_shr_cnt[2]), .Z(N2876) );
  GTECH_OR2 C5399 ( .A(a2stg_nx_neq0_84_tmp_3[63]), .B(a2stg_shr_cnt[2]), .Z(
        N2878) );
  GTECH_NOT I_453 ( .A(N2882), .Z(a2stg_nx_neq0_84_tmp_4[62]) );
  GTECH_AND2 C5401 ( .A(N2880), .B(N2881), .Z(N2882) );
  GTECH_OR2 C5402 ( .A(a2stg_shr_tmp6[14]), .B(N2876), .Z(N2880) );
  GTECH_OR2 C5404 ( .A(a2stg_nx_neq0_84_tmp_3[62]), .B(a2stg_shr_cnt[2]), .Z(
        N2881) );
  GTECH_NOT I_454 ( .A(N2885), .Z(a2stg_nx_neq0_84_tmp_4[61]) );
  GTECH_AND2 C5406 ( .A(N2883), .B(N2884), .Z(N2885) );
  GTECH_OR2 C5407 ( .A(a2stg_shr_tmp6[13]), .B(N2876), .Z(N2883) );
  GTECH_OR2 C5409 ( .A(a2stg_nx_neq0_84_tmp_3[61]), .B(a2stg_shr_cnt[2]), .Z(
        N2884) );
  GTECH_NOT I_455 ( .A(N2888), .Z(a2stg_nx_neq0_84_tmp_4[60]) );
  GTECH_AND2 C5411 ( .A(N2886), .B(N2887), .Z(N2888) );
  GTECH_OR2 C5412 ( .A(a2stg_shr_tmp6[12]), .B(N2876), .Z(N2886) );
  GTECH_OR2 C5414 ( .A(a2stg_nx_neq0_84_tmp_3[60]), .B(a2stg_shr_cnt[2]), .Z(
        N2887) );
  GTECH_NOT I_456 ( .A(N2891), .Z(a2stg_nx_neq0_84_tmp_4[59]) );
  GTECH_AND2 C5416 ( .A(N2889), .B(N2890), .Z(N2891) );
  GTECH_OR2 C5417 ( .A(a2stg_nx_neq0_84_tmp_3[63]), .B(N2876), .Z(N2889) );
  GTECH_OR2 C5419 ( .A(a2stg_nx_neq0_84_tmp_3[59]), .B(a2stg_shr_cnt[2]), .Z(
        N2890) );
  GTECH_NOT I_457 ( .A(N2894), .Z(a2stg_nx_neq0_84_tmp_4[58]) );
  GTECH_AND2 C5421 ( .A(N2892), .B(N2893), .Z(N2894) );
  GTECH_OR2 C5422 ( .A(a2stg_nx_neq0_84_tmp_3[62]), .B(N2876), .Z(N2892) );
  GTECH_OR2 C5424 ( .A(a2stg_nx_neq0_84_tmp_3[58]), .B(a2stg_shr_cnt[2]), .Z(
        N2893) );
  GTECH_NOT I_458 ( .A(N2897), .Z(a2stg_nx_neq0_84_tmp_4[57]) );
  GTECH_AND2 C5426 ( .A(N2895), .B(N2896), .Z(N2897) );
  GTECH_OR2 C5427 ( .A(a2stg_nx_neq0_84_tmp_3[61]), .B(N2876), .Z(N2895) );
  GTECH_OR2 C5429 ( .A(a2stg_nx_neq0_84_tmp_3[57]), .B(a2stg_shr_cnt[2]), .Z(
        N2896) );
  GTECH_NOT I_459 ( .A(N2900), .Z(a2stg_nx_neq0_84_tmp_4_54) );
  GTECH_AND2 C5431 ( .A(N2898), .B(N2899), .Z(N2900) );
  GTECH_OR2 C5432 ( .A(a2stg_nx_neq0_84_tmp_3[58]), .B(N2876), .Z(N2898) );
  GTECH_OR2 C5434 ( .A(a2stg_nx_neq0_84_tmp_3[54]), .B(a2stg_shr_cnt[2]), .Z(
        N2899) );
  GTECH_NOT I_460 ( .A(N2903), .Z(a2stg_nx_neq0_84_tmp_4_53) );
  GTECH_AND2 C5436 ( .A(N2901), .B(N2902), .Z(N2903) );
  GTECH_OR2 C5437 ( .A(a2stg_nx_neq0_84_tmp_3[57]), .B(N2876), .Z(N2901) );
  GTECH_OR2 C5439 ( .A(a2stg_nx_neq0_84_tmp_3[53]), .B(a2stg_shr_cnt[2]), .Z(
        N2902) );
  GTECH_NOT I_461 ( .A(N2906), .Z(a2stg_nx_neq0_84_tmp_4_52) );
  GTECH_AND2 C5441 ( .A(N2904), .B(N2905), .Z(N2906) );
  GTECH_OR2 C5442 ( .A(a2stg_nx_neq0_84_tmp_3[56]), .B(N2876), .Z(N2904) );
  GTECH_OR2 C5444 ( .A(a2stg_nx_neq0_84_tmp_3[52]), .B(a2stg_shr_cnt[2]), .Z(
        N2905) );
  GTECH_NOT I_462 ( .A(N2909), .Z(a2stg_nx_neq0_84_tmp_4_51) );
  GTECH_AND2 C5446 ( .A(N2907), .B(N2908), .Z(N2909) );
  GTECH_OR2 C5447 ( .A(a2stg_nx_neq0_84_tmp_3[55]), .B(N2876), .Z(N2907) );
  GTECH_OR2 C5449 ( .A(a2stg_nx_neq0_84_tmp_3[51]), .B(a2stg_shr_cnt[2]), .Z(
        N2908) );
  GTECH_NOT I_463 ( .A(N2912), .Z(a2stg_nx_neq0_84_tmp_4_50) );
  GTECH_AND2 C5451 ( .A(N2910), .B(N2911), .Z(N2912) );
  GTECH_OR2 C5452 ( .A(a2stg_nx_neq0_84_tmp_3[54]), .B(N2876), .Z(N2910) );
  GTECH_OR2 C5454 ( .A(a2stg_nx_neq0_84_tmp_3[50]), .B(a2stg_shr_cnt[2]), .Z(
        N2911) );
  GTECH_NOT I_464 ( .A(N2915), .Z(a2stg_nx_neq0_84_tmp_4_49) );
  GTECH_AND2 C5456 ( .A(N2913), .B(N2914), .Z(N2915) );
  GTECH_OR2 C5457 ( .A(a2stg_nx_neq0_84_tmp_3[53]), .B(N2876), .Z(N2913) );
  GTECH_OR2 C5459 ( .A(a2stg_nx_neq0_84_tmp_3[49]), .B(a2stg_shr_cnt[2]), .Z(
        N2914) );
  GTECH_NOT I_465 ( .A(N2918), .Z(a2stg_nx_neq0_84_tmp_4_48) );
  GTECH_AND2 C5461 ( .A(N2916), .B(N2917), .Z(N2918) );
  GTECH_OR2 C5462 ( .A(a2stg_nx_neq0_84_tmp_3[52]), .B(N2876), .Z(N2916) );
  GTECH_OR2 C5464 ( .A(a2stg_nx_neq0_84_tmp_3[48]), .B(a2stg_shr_cnt[2]), .Z(
        N2917) );
  GTECH_NOT I_466 ( .A(N2922), .Z(a2stg_nx_neq0_84_tmp_5[61]) );
  GTECH_OR2 C5466 ( .A(N2919), .B(N2921), .Z(N2922) );
  GTECH_AND2 C5467 ( .A(a2stg_nx_neq0_84_tmp_4[63]), .B(a2stg_shr_cnt[1]), .Z(
        N2919) );
  GTECH_AND2 C5468 ( .A(a2stg_nx_neq0_84_tmp_4[61]), .B(N2920), .Z(N2921) );
  GTECH_NOT I_467 ( .A(a2stg_shr_cnt[1]), .Z(N2920) );
  GTECH_NOT I_468 ( .A(N2925), .Z(a2stg_nx_neq0_84_tmp_5[60]) );
  GTECH_OR2 C5471 ( .A(N2923), .B(N2924), .Z(N2925) );
  GTECH_AND2 C5472 ( .A(a2stg_nx_neq0_84_tmp_4[62]), .B(a2stg_shr_cnt[1]), .Z(
        N2923) );
  GTECH_AND2 C5473 ( .A(a2stg_nx_neq0_84_tmp_4[60]), .B(N2920), .Z(N2924) );
  GTECH_NOT I_469 ( .A(N2928), .Z(a2stg_nx_neq0_84_tmp_5[59]) );
  GTECH_OR2 C5476 ( .A(N2926), .B(N2927), .Z(N2928) );
  GTECH_AND2 C5477 ( .A(a2stg_nx_neq0_84_tmp_4[61]), .B(a2stg_shr_cnt[1]), .Z(
        N2926) );
  GTECH_AND2 C5478 ( .A(a2stg_nx_neq0_84_tmp_4[59]), .B(N2920), .Z(N2927) );
  GTECH_NOT I_470 ( .A(N2931), .Z(a2stg_nx_neq0_84_tmp_5_52) );
  GTECH_OR2 C5481 ( .A(N2929), .B(N2930), .Z(N2931) );
  GTECH_AND2 C5482 ( .A(a2stg_nx_neq0_84_tmp_4_54), .B(a2stg_shr_cnt[1]), .Z(
        N2929) );
  GTECH_AND2 C5483 ( .A(a2stg_nx_neq0_84_tmp_4_52), .B(N2920), .Z(N2930) );
  GTECH_NOT I_471 ( .A(N2934), .Z(a2stg_nx_neq0_84_tmp_5_51) );
  GTECH_OR2 C5486 ( .A(N2932), .B(N2933), .Z(N2934) );
  GTECH_AND2 C5487 ( .A(a2stg_nx_neq0_84_tmp_4_53), .B(a2stg_shr_cnt[1]), .Z(
        N2932) );
  GTECH_AND2 C5488 ( .A(a2stg_nx_neq0_84_tmp_4_51), .B(N2920), .Z(N2933) );
  GTECH_NOT I_472 ( .A(N2937), .Z(a2stg_nx_neq0_84_tmp_5_50) );
  GTECH_OR2 C5491 ( .A(N2935), .B(N2936), .Z(N2937) );
  GTECH_AND2 C5492 ( .A(a2stg_nx_neq0_84_tmp_4_52), .B(a2stg_shr_cnt[1]), .Z(
        N2935) );
  GTECH_AND2 C5493 ( .A(a2stg_nx_neq0_84_tmp_4_50), .B(N2920), .Z(N2936) );
  GTECH_NOT I_473 ( .A(N2938), .Z(a2stg_nx_neq0_84_tmp_6[59]) );
  GTECH_OR2 C5496 ( .A(a2stg_shr_cnt[0]), .B(a2stg_nx_neq0_84_tmp_5[60]), .Z(
        N2938) );
  GTECH_NOT I_474 ( .A(N2940), .Z(a2stg_nx_neq0_84_tmp_6[60]) );
  GTECH_OR2 C5498 ( .A(N2939), .B(a2stg_nx_neq0_84_tmp_5[61]), .Z(N2940) );
  GTECH_NOT I_475 ( .A(a2stg_shr_cnt[0]), .Z(N2939) );
  GTECH_NOT I_476 ( .A(N2943), .Z(a2stg_nx_neq0_84_tmp_6_51) );
  GTECH_AND2 C5501 ( .A(N2941), .B(N2942), .Z(N2943) );
  GTECH_OR2 C5502 ( .A(a2stg_nx_neq0_84_tmp_5_52), .B(N2939), .Z(N2941) );
  GTECH_OR2 C5504 ( .A(a2stg_nx_neq0_84_tmp_5_51), .B(a2stg_shr_cnt[0]), .Z(
        N2942) );
  GTECH_OR2 C5505 ( .A(N3007), .B(a2stg_nx_neq0_84_tmp_6_51), .Z(
        a2stg_fsdtoix_nx) );
  GTECH_OR2 C5506 ( .A(N3004), .B(N3006), .Z(N3007) );
  GTECH_OR2 C5507 ( .A(N3000), .B(N3003), .Z(N3004) );
  GTECH_OR2 C5508 ( .A(N2991), .B(N2999), .Z(N3000) );
  GTECH_OR2 C5509 ( .A(N2975), .B(N2990), .Z(N2991) );
  GTECH_NOT I_477 ( .A(N2974), .Z(N2975) );
  GTECH_AND2 C5511 ( .A(N2973), .B(a2stg_nx_neq0_84_tmp_1[20]), .Z(N2974) );
  GTECH_AND2 C5512 ( .A(N2972), .B(a2stg_nx_neq0_84_tmp_1[21]), .Z(N2973) );
  GTECH_AND2 C5513 ( .A(N2971), .B(a2stg_nx_neq0_84_tmp_1[22]), .Z(N2972) );
  GTECH_AND2 C5514 ( .A(N2970), .B(a2stg_nx_neq0_84_tmp_1[23]), .Z(N2971) );
  GTECH_AND2 C5515 ( .A(N2969), .B(a2stg_nx_neq0_84_tmp_1[24]), .Z(N2970) );
  GTECH_AND2 C5516 ( .A(N2968), .B(a2stg_nx_neq0_84_tmp_1[25]), .Z(N2969) );
  GTECH_AND2 C5517 ( .A(N2967), .B(a2stg_nx_neq0_84_tmp_1[26]), .Z(N2968) );
  GTECH_AND2 C5518 ( .A(N2966), .B(a2stg_nx_neq0_84_tmp_1[27]), .Z(N2967) );
  GTECH_AND2 C5519 ( .A(N2965), .B(a2stg_nx_neq0_84_tmp_1[28]), .Z(N2966) );
  GTECH_AND2 C5520 ( .A(N2964), .B(a2stg_nx_neq0_84_tmp_1[29]), .Z(N2965) );
  GTECH_AND2 C5521 ( .A(N2963), .B(a2stg_nx_neq0_84_tmp_1[30]), .Z(N2964) );
  GTECH_AND2 C5522 ( .A(N2962), .B(a2stg_nx_neq0_84_tmp_1[31]), .Z(N2963) );
  GTECH_AND2 C5523 ( .A(N2961), .B(a2stg_nx_neq0_84_tmp_1[32]), .Z(N2962) );
  GTECH_AND2 C5524 ( .A(N2960), .B(a2stg_nx_neq0_84_tmp_1[33]), .Z(N2961) );
  GTECH_AND2 C5525 ( .A(N2959), .B(a2stg_nx_neq0_84_tmp_1[34]), .Z(N2960) );
  GTECH_AND2 C5526 ( .A(N2958), .B(a2stg_nx_neq0_84_tmp_1[35]), .Z(N2959) );
  GTECH_AND2 C5527 ( .A(N2957), .B(a2stg_nx_neq0_84_tmp_1[36]), .Z(N2958) );
  GTECH_AND2 C5528 ( .A(N2956), .B(a2stg_nx_neq0_84_tmp_1[37]), .Z(N2957) );
  GTECH_AND2 C5529 ( .A(N2955), .B(a2stg_nx_neq0_84_tmp_1[38]), .Z(N2956) );
  GTECH_AND2 C5530 ( .A(N2954), .B(a2stg_nx_neq0_84_tmp_1[39]), .Z(N2955) );
  GTECH_AND2 C5531 ( .A(N2953), .B(a2stg_nx_neq0_84_tmp_1[40]), .Z(N2954) );
  GTECH_AND2 C5532 ( .A(N2952), .B(a2stg_nx_neq0_84_tmp_1[41]), .Z(N2953) );
  GTECH_AND2 C5533 ( .A(N2951), .B(a2stg_nx_neq0_84_tmp_1[42]), .Z(N2952) );
  GTECH_AND2 C5534 ( .A(N2950), .B(a2stg_nx_neq0_84_tmp_1[43]), .Z(N2951) );
  GTECH_AND2 C5535 ( .A(N2949), .B(a2stg_nx_neq0_84_tmp_1[44]), .Z(N2950) );
  GTECH_AND2 C5536 ( .A(N2948), .B(a2stg_nx_neq0_84_tmp_1[45]), .Z(N2949) );
  GTECH_AND2 C5537 ( .A(N2947), .B(a2stg_nx_neq0_84_tmp_1[46]), .Z(N2948) );
  GTECH_AND2 C5538 ( .A(N2946), .B(a2stg_nx_neq0_84_tmp_1[47]), .Z(N2947) );
  GTECH_AND2 C5539 ( .A(N2945), .B(a2stg_nx_neq0_84_tmp_1[48]), .Z(N2946) );
  GTECH_AND2 C5540 ( .A(N2944), .B(a2stg_nx_neq0_84_tmp_1[49]), .Z(N2945) );
  GTECH_AND2 C5541 ( .A(a2stg_nx_neq0_84_tmp_1[51]), .B(
        a2stg_nx_neq0_84_tmp_1[50]), .Z(N2944) );
  GTECH_OR2 C5542 ( .A(N2989), .B(a2stg_nx_neq0_84_tmp_2[36]), .Z(N2990) );
  GTECH_OR2 C5543 ( .A(N2988), .B(a2stg_nx_neq0_84_tmp_2[37]), .Z(N2989) );
  GTECH_OR2 C5544 ( .A(N2987), .B(a2stg_nx_neq0_84_tmp_2[38]), .Z(N2988) );
  GTECH_OR2 C5545 ( .A(N2986), .B(a2stg_nx_neq0_84_tmp_2[39]), .Z(N2987) );
  GTECH_OR2 C5546 ( .A(N2985), .B(a2stg_nx_neq0_84_tmp_2[40]), .Z(N2986) );
  GTECH_OR2 C5547 ( .A(N2984), .B(a2stg_nx_neq0_84_tmp_2[41]), .Z(N2985) );
  GTECH_OR2 C5548 ( .A(N2983), .B(a2stg_nx_neq0_84_tmp_2[42]), .Z(N2984) );
  GTECH_OR2 C5549 ( .A(N2982), .B(a2stg_nx_neq0_84_tmp_2[43]), .Z(N2983) );
  GTECH_OR2 C5550 ( .A(N2981), .B(a2stg_nx_neq0_84_tmp_2[44]), .Z(N2982) );
  GTECH_OR2 C5551 ( .A(N2980), .B(a2stg_nx_neq0_84_tmp_2[45]), .Z(N2981) );
  GTECH_OR2 C5552 ( .A(N2979), .B(a2stg_nx_neq0_84_tmp_2[46]), .Z(N2980) );
  GTECH_OR2 C5553 ( .A(N2978), .B(a2stg_nx_neq0_84_tmp_2[47]), .Z(N2979) );
  GTECH_OR2 C5554 ( .A(N2977), .B(a2stg_nx_neq0_84_tmp_2[48]), .Z(N2978) );
  GTECH_OR2 C5555 ( .A(N2976), .B(a2stg_nx_neq0_84_tmp_2[49]), .Z(N2977) );
  GTECH_OR2 C5556 ( .A(a2stg_nx_neq0_84_tmp_2[51]), .B(
        a2stg_nx_neq0_84_tmp_2[50]), .Z(N2976) );
  GTECH_NOT I_478 ( .A(N2998), .Z(N2999) );
  GTECH_AND2 C5558 ( .A(N2997), .B(a2stg_nx_neq0_84_tmp_3[44]), .Z(N2998) );
  GTECH_AND2 C5559 ( .A(N2996), .B(a2stg_nx_neq0_84_tmp_3[45]), .Z(N2997) );
  GTECH_AND2 C5560 ( .A(N2995), .B(a2stg_nx_neq0_84_tmp_3[46]), .Z(N2996) );
  GTECH_AND2 C5561 ( .A(N2994), .B(a2stg_nx_neq0_84_tmp_3[47]), .Z(N2995) );
  GTECH_AND2 C5562 ( .A(N2993), .B(a2stg_nx_neq0_84_tmp_3[48]), .Z(N2994) );
  GTECH_AND2 C5563 ( .A(N2992), .B(a2stg_nx_neq0_84_tmp_3[49]), .Z(N2993) );
  GTECH_AND2 C5564 ( .A(a2stg_nx_neq0_84_tmp_3[51]), .B(
        a2stg_nx_neq0_84_tmp_3[50]), .Z(N2992) );
  GTECH_OR2 C5565 ( .A(N3002), .B(a2stg_nx_neq0_84_tmp_4_48), .Z(N3003) );
  GTECH_OR2 C5566 ( .A(N3001), .B(a2stg_nx_neq0_84_tmp_4_49), .Z(N3002) );
  GTECH_OR2 C5567 ( .A(a2stg_nx_neq0_84_tmp_4_51), .B(
        a2stg_nx_neq0_84_tmp_4_50), .Z(N3001) );
  GTECH_NOT I_479 ( .A(N3005), .Z(N3006) );
  GTECH_AND2 C5569 ( .A(a2stg_nx_neq0_84_tmp_5_51), .B(
        a2stg_nx_neq0_84_tmp_5_50), .Z(N3005) );
  GTECH_OR2 C5570 ( .A(N3080), .B(N3081), .Z(a2stg_shr_60_0_neq_0) );
  GTECH_OR2 C5571 ( .A(N3077), .B(N3079), .Z(N3080) );
  GTECH_OR2 C5572 ( .A(N3073), .B(N3076), .Z(N3077) );
  GTECH_OR2 C5573 ( .A(N3064), .B(N3072), .Z(N3073) );
  GTECH_OR2 C5574 ( .A(N3048), .B(N3063), .Z(N3064) );
  GTECH_NOT I_480 ( .A(N3047), .Z(N3048) );
  GTECH_AND2 C5576 ( .A(N3046), .B(a2stg_nx_neq0_84_tmp_1[20]), .Z(N3047) );
  GTECH_AND2 C5577 ( .A(N3045), .B(a2stg_nx_neq0_84_tmp_1[21]), .Z(N3046) );
  GTECH_AND2 C5578 ( .A(N3044), .B(a2stg_nx_neq0_84_tmp_1[22]), .Z(N3045) );
  GTECH_AND2 C5579 ( .A(N3043), .B(a2stg_nx_neq0_84_tmp_1[23]), .Z(N3044) );
  GTECH_AND2 C5580 ( .A(N3042), .B(a2stg_nx_neq0_84_tmp_1[24]), .Z(N3043) );
  GTECH_AND2 C5581 ( .A(N3041), .B(a2stg_nx_neq0_84_tmp_1[25]), .Z(N3042) );
  GTECH_AND2 C5582 ( .A(N3040), .B(a2stg_nx_neq0_84_tmp_1[26]), .Z(N3041) );
  GTECH_AND2 C5583 ( .A(N3039), .B(a2stg_nx_neq0_84_tmp_1[27]), .Z(N3040) );
  GTECH_AND2 C5584 ( .A(N3038), .B(a2stg_nx_neq0_84_tmp_1[28]), .Z(N3039) );
  GTECH_AND2 C5585 ( .A(N3037), .B(a2stg_nx_neq0_84_tmp_1[29]), .Z(N3038) );
  GTECH_AND2 C5586 ( .A(N3036), .B(a2stg_nx_neq0_84_tmp_1[30]), .Z(N3037) );
  GTECH_AND2 C5587 ( .A(N3035), .B(a2stg_nx_neq0_84_tmp_1[31]), .Z(N3036) );
  GTECH_AND2 C5588 ( .A(N3034), .B(a2stg_nx_neq0_84_tmp_1[32]), .Z(N3035) );
  GTECH_AND2 C5589 ( .A(N3033), .B(a2stg_nx_neq0_84_tmp_1[33]), .Z(N3034) );
  GTECH_AND2 C5590 ( .A(N3032), .B(a2stg_nx_neq0_84_tmp_1[34]), .Z(N3033) );
  GTECH_AND2 C5591 ( .A(N3031), .B(a2stg_nx_neq0_84_tmp_1[35]), .Z(N3032) );
  GTECH_AND2 C5592 ( .A(N3030), .B(a2stg_nx_neq0_84_tmp_1[36]), .Z(N3031) );
  GTECH_AND2 C5593 ( .A(N3029), .B(a2stg_nx_neq0_84_tmp_1[37]), .Z(N3030) );
  GTECH_AND2 C5594 ( .A(N3028), .B(a2stg_nx_neq0_84_tmp_1[38]), .Z(N3029) );
  GTECH_AND2 C5595 ( .A(N3027), .B(a2stg_nx_neq0_84_tmp_1[39]), .Z(N3028) );
  GTECH_AND2 C5596 ( .A(N3026), .B(a2stg_nx_neq0_84_tmp_1[40]), .Z(N3027) );
  GTECH_AND2 C5597 ( .A(N3025), .B(a2stg_nx_neq0_84_tmp_1[41]), .Z(N3026) );
  GTECH_AND2 C5598 ( .A(N3024), .B(a2stg_nx_neq0_84_tmp_1[42]), .Z(N3025) );
  GTECH_AND2 C5599 ( .A(N3023), .B(a2stg_nx_neq0_84_tmp_1[43]), .Z(N3024) );
  GTECH_AND2 C5600 ( .A(N3022), .B(a2stg_nx_neq0_84_tmp_1[44]), .Z(N3023) );
  GTECH_AND2 C5601 ( .A(N3021), .B(a2stg_nx_neq0_84_tmp_1[45]), .Z(N3022) );
  GTECH_AND2 C5602 ( .A(N3020), .B(a2stg_nx_neq0_84_tmp_1[46]), .Z(N3021) );
  GTECH_AND2 C5603 ( .A(N3019), .B(a2stg_nx_neq0_84_tmp_1[47]), .Z(N3020) );
  GTECH_AND2 C5604 ( .A(N3018), .B(a2stg_nx_neq0_84_tmp_1[48]), .Z(N3019) );
  GTECH_AND2 C5605 ( .A(N3017), .B(a2stg_nx_neq0_84_tmp_1[49]), .Z(N3018) );
  GTECH_AND2 C5606 ( .A(N3016), .B(a2stg_nx_neq0_84_tmp_1[50]), .Z(N3017) );
  GTECH_AND2 C5607 ( .A(N3015), .B(a2stg_nx_neq0_84_tmp_1[51]), .Z(N3016) );
  GTECH_AND2 C5608 ( .A(N3014), .B(a2stg_nx_neq0_84_tmp_1[52]), .Z(N3015) );
  GTECH_AND2 C5609 ( .A(N3013), .B(a2stg_nx_neq0_84_tmp_1[53]), .Z(N3014) );
  GTECH_AND2 C5610 ( .A(N3012), .B(a2stg_nx_neq0_84_tmp_1[54]), .Z(N3013) );
  GTECH_AND2 C5611 ( .A(N3011), .B(a2stg_nx_neq0_84_tmp_1[55]), .Z(N3012) );
  GTECH_AND2 C5612 ( .A(N3010), .B(a2stg_nx_neq0_84_tmp_1[56]), .Z(N3011) );
  GTECH_AND2 C5613 ( .A(N3009), .B(a2stg_nx_neq0_84_tmp_1[57]), .Z(N3010) );
  GTECH_AND2 C5614 ( .A(N3008), .B(a2stg_nx_neq0_84_tmp_1[58]), .Z(N3009) );
  GTECH_AND2 C5615 ( .A(a2stg_nx_neq0_84_tmp_1[60]), .B(
        a2stg_nx_neq0_84_tmp_1[59]), .Z(N3008) );
  GTECH_OR2 C5616 ( .A(N3062), .B(a2stg_nx_neq0_84_tmp_2[45]), .Z(N3063) );
  GTECH_OR2 C5617 ( .A(N3061), .B(a2stg_nx_neq0_84_tmp_2[46]), .Z(N3062) );
  GTECH_OR2 C5618 ( .A(N3060), .B(a2stg_nx_neq0_84_tmp_2[47]), .Z(N3061) );
  GTECH_OR2 C5619 ( .A(N3059), .B(a2stg_nx_neq0_84_tmp_2[48]), .Z(N3060) );
  GTECH_OR2 C5620 ( .A(N3058), .B(a2stg_nx_neq0_84_tmp_2[49]), .Z(N3059) );
  GTECH_OR2 C5621 ( .A(N3057), .B(a2stg_nx_neq0_84_tmp_2[50]), .Z(N3058) );
  GTECH_OR2 C5622 ( .A(N3056), .B(a2stg_nx_neq0_84_tmp_2[51]), .Z(N3057) );
  GTECH_OR2 C5623 ( .A(N3055), .B(a2stg_nx_neq0_84_tmp_2[52]), .Z(N3056) );
  GTECH_OR2 C5624 ( .A(N3054), .B(a2stg_nx_neq0_84_tmp_2[53]), .Z(N3055) );
  GTECH_OR2 C5625 ( .A(N3053), .B(a2stg_nx_neq0_84_tmp_2[54]), .Z(N3054) );
  GTECH_OR2 C5626 ( .A(N3052), .B(a2stg_nx_neq0_84_tmp_2[55]), .Z(N3053) );
  GTECH_OR2 C5627 ( .A(N3051), .B(a2stg_nx_neq0_84_tmp_2[56]), .Z(N3052) );
  GTECH_OR2 C5628 ( .A(N3050), .B(a2stg_nx_neq0_84_tmp_2[57]), .Z(N3051) );
  GTECH_OR2 C5629 ( .A(N3049), .B(a2stg_nx_neq0_84_tmp_2[58]), .Z(N3050) );
  GTECH_OR2 C5630 ( .A(a2stg_nx_neq0_84_tmp_2[60]), .B(
        a2stg_nx_neq0_84_tmp_2[59]), .Z(N3049) );
  GTECH_NOT I_481 ( .A(N3071), .Z(N3072) );
  GTECH_AND2 C5632 ( .A(N3070), .B(a2stg_nx_neq0_84_tmp_3[53]), .Z(N3071) );
  GTECH_AND2 C5633 ( .A(N3069), .B(a2stg_nx_neq0_84_tmp_3[54]), .Z(N3070) );
  GTECH_AND2 C5634 ( .A(N3068), .B(a2stg_nx_neq0_84_tmp_3[55]), .Z(N3069) );
  GTECH_AND2 C5635 ( .A(N3067), .B(a2stg_nx_neq0_84_tmp_3[56]), .Z(N3068) );
  GTECH_AND2 C5636 ( .A(N3066), .B(a2stg_nx_neq0_84_tmp_3[57]), .Z(N3067) );
  GTECH_AND2 C5637 ( .A(N3065), .B(a2stg_nx_neq0_84_tmp_3[58]), .Z(N3066) );
  GTECH_AND2 C5638 ( .A(a2stg_nx_neq0_84_tmp_3[60]), .B(
        a2stg_nx_neq0_84_tmp_3[59]), .Z(N3065) );
  GTECH_OR2 C5639 ( .A(N3075), .B(a2stg_nx_neq0_84_tmp_4[57]), .Z(N3076) );
  GTECH_OR2 C5640 ( .A(N3074), .B(a2stg_nx_neq0_84_tmp_4[58]), .Z(N3075) );
  GTECH_OR2 C5641 ( .A(a2stg_nx_neq0_84_tmp_4[60]), .B(
        a2stg_nx_neq0_84_tmp_4[59]), .Z(N3074) );
  GTECH_NOT I_482 ( .A(N3078), .Z(N3079) );
  GTECH_AND2 C5643 ( .A(a2stg_nx_neq0_84_tmp_5[60]), .B(
        a2stg_nx_neq0_84_tmp_5[59]), .Z(N3078) );
  GTECH_OR2 C5644 ( .A(a2stg_nx_neq0_84_tmp_6[60]), .B(
        a2stg_nx_neq0_84_tmp_6[59]), .Z(N3081) );
  GTECH_NOT I_483 ( .A(N3089), .Z(a2stg_shr_frac2_inv[63]) );
  GTECH_OR2 C5646 ( .A(N3086), .B(N3088), .Z(N3089) );
  GTECH_OR2 C5647 ( .A(N3083), .B(N3085), .Z(N3086) );
  GTECH_AND2 C5648 ( .A(N3082), .B(a2stg_shr[115]), .Z(N3083) );
  GTECH_AND2 C5649 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3082) );
  GTECH_AND2 C5650 ( .A(N3084), .B(a2stg_shr[115]), .Z(N3085) );
  GTECH_AND2 C5651 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3084) );
  GTECH_AND2 C5652 ( .A(N3087), .B(a3stg_frac2[63]), .Z(N3088) );
  GTECH_NOT I_484 ( .A(a6stg_step), .Z(N3087) );
  GTECH_NOT I_485 ( .A(N3102), .Z(a2stg_shr_frac2_inv[62]) );
  GTECH_OR2 C5655 ( .A(N3099), .B(N3101), .Z(N3102) );
  GTECH_OR2 C5656 ( .A(N3096), .B(N3098), .Z(N3099) );
  GTECH_OR2 C5657 ( .A(N3093), .B(N3095), .Z(N3096) );
  GTECH_OR2 C5658 ( .A(N3090), .B(N3092), .Z(N3093) );
  GTECH_AND2 C5659 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[115]), .Z(N3090) );
  GTECH_AND2 C5660 ( .A(N3091), .B(a2stg_shr[114]), .Z(N3092) );
  GTECH_AND2 C5661 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3091) );
  GTECH_AND2 C5662 ( .A(N3094), .B(a2stg_shr[114]), .Z(N3095) );
  GTECH_AND2 C5663 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3094) );
  GTECH_AND2 C5664 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3098) );
  GTECH_NOT I_486 ( .A(a2stg_expadd_11), .Z(N3097) );
  GTECH_AND2 C5666 ( .A(N3100), .B(a3stg_frac2[62]), .Z(N3101) );
  GTECH_NOT I_487 ( .A(a6stg_step), .Z(N3100) );
  GTECH_NOT I_488 ( .A(N3114), .Z(a2stg_shr_frac2_inv[61]) );
  GTECH_OR2 C5669 ( .A(N3111), .B(N3113), .Z(N3114) );
  GTECH_OR2 C5670 ( .A(N3109), .B(N3110), .Z(N3111) );
  GTECH_OR2 C5671 ( .A(N3106), .B(N3108), .Z(N3109) );
  GTECH_OR2 C5672 ( .A(N3103), .B(N3105), .Z(N3106) );
  GTECH_AND2 C5673 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[114]), .Z(N3103) );
  GTECH_AND2 C5674 ( .A(N3104), .B(a2stg_shr[113]), .Z(N3105) );
  GTECH_AND2 C5675 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3104) );
  GTECH_AND2 C5676 ( .A(N3107), .B(a2stg_shr[113]), .Z(N3108) );
  GTECH_AND2 C5677 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3107) );
  GTECH_AND2 C5678 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3110) );
  GTECH_AND2 C5680 ( .A(N3112), .B(a3stg_frac2[61]), .Z(N3113) );
  GTECH_NOT I_489 ( .A(a6stg_step), .Z(N3112) );
  GTECH_NOT I_490 ( .A(N3126), .Z(a2stg_shr_frac2_inv[60]) );
  GTECH_OR2 C5683 ( .A(N3123), .B(N3125), .Z(N3126) );
  GTECH_OR2 C5684 ( .A(N3121), .B(N3122), .Z(N3123) );
  GTECH_OR2 C5685 ( .A(N3118), .B(N3120), .Z(N3121) );
  GTECH_OR2 C5686 ( .A(N3115), .B(N3117), .Z(N3118) );
  GTECH_AND2 C5687 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[113]), .Z(N3115) );
  GTECH_AND2 C5688 ( .A(N3116), .B(a2stg_shr[112]), .Z(N3117) );
  GTECH_AND2 C5689 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3116) );
  GTECH_AND2 C5690 ( .A(N3119), .B(a2stg_shr[112]), .Z(N3120) );
  GTECH_AND2 C5691 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3119) );
  GTECH_AND2 C5692 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3122) );
  GTECH_AND2 C5694 ( .A(N3124), .B(a3stg_frac2[60]), .Z(N3125) );
  GTECH_NOT I_491 ( .A(a6stg_step), .Z(N3124) );
  GTECH_NOT I_492 ( .A(N3138), .Z(a2stg_shr_frac2_inv[59]) );
  GTECH_OR2 C5697 ( .A(N3135), .B(N3137), .Z(N3138) );
  GTECH_OR2 C5698 ( .A(N3133), .B(N3134), .Z(N3135) );
  GTECH_OR2 C5699 ( .A(N3130), .B(N3132), .Z(N3133) );
  GTECH_OR2 C5700 ( .A(N3127), .B(N3129), .Z(N3130) );
  GTECH_AND2 C5701 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[112]), .Z(N3127) );
  GTECH_AND2 C5702 ( .A(N3128), .B(a2stg_shr[111]), .Z(N3129) );
  GTECH_AND2 C5703 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3128) );
  GTECH_AND2 C5704 ( .A(N3131), .B(a2stg_shr[111]), .Z(N3132) );
  GTECH_AND2 C5705 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3131) );
  GTECH_AND2 C5706 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3134) );
  GTECH_AND2 C5708 ( .A(N3136), .B(a3stg_frac2[59]), .Z(N3137) );
  GTECH_NOT I_493 ( .A(a6stg_step), .Z(N3136) );
  GTECH_NOT I_494 ( .A(N3150), .Z(a2stg_shr_frac2_inv[58]) );
  GTECH_OR2 C5711 ( .A(N3147), .B(N3149), .Z(N3150) );
  GTECH_OR2 C5712 ( .A(N3145), .B(N3146), .Z(N3147) );
  GTECH_OR2 C5713 ( .A(N3142), .B(N3144), .Z(N3145) );
  GTECH_OR2 C5714 ( .A(N3139), .B(N3141), .Z(N3142) );
  GTECH_AND2 C5715 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[111]), .Z(N3139) );
  GTECH_AND2 C5716 ( .A(N3140), .B(a2stg_shr[110]), .Z(N3141) );
  GTECH_AND2 C5717 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3140) );
  GTECH_AND2 C5718 ( .A(N3143), .B(a2stg_shr[110]), .Z(N3144) );
  GTECH_AND2 C5719 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3143) );
  GTECH_AND2 C5720 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3146) );
  GTECH_AND2 C5722 ( .A(N3148), .B(a3stg_frac2[58]), .Z(N3149) );
  GTECH_NOT I_495 ( .A(a6stg_step), .Z(N3148) );
  GTECH_NOT I_496 ( .A(N3162), .Z(a2stg_shr_frac2_inv[57]) );
  GTECH_OR2 C5725 ( .A(N3159), .B(N3161), .Z(N3162) );
  GTECH_OR2 C5726 ( .A(N3157), .B(N3158), .Z(N3159) );
  GTECH_OR2 C5727 ( .A(N3154), .B(N3156), .Z(N3157) );
  GTECH_OR2 C5728 ( .A(N3151), .B(N3153), .Z(N3154) );
  GTECH_AND2 C5729 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[110]), .Z(N3151) );
  GTECH_AND2 C5730 ( .A(N3152), .B(a2stg_shr[109]), .Z(N3153) );
  GTECH_AND2 C5731 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3152) );
  GTECH_AND2 C5732 ( .A(N3155), .B(a2stg_shr[109]), .Z(N3156) );
  GTECH_AND2 C5733 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3155) );
  GTECH_AND2 C5734 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3158) );
  GTECH_AND2 C5736 ( .A(N3160), .B(a3stg_frac2[57]), .Z(N3161) );
  GTECH_NOT I_497 ( .A(a6stg_step), .Z(N3160) );
  GTECH_NOT I_498 ( .A(N3174), .Z(a2stg_shr_frac2_inv[56]) );
  GTECH_OR2 C5739 ( .A(N3171), .B(N3173), .Z(N3174) );
  GTECH_OR2 C5740 ( .A(N3169), .B(N3170), .Z(N3171) );
  GTECH_OR2 C5741 ( .A(N3166), .B(N3168), .Z(N3169) );
  GTECH_OR2 C5742 ( .A(N3163), .B(N3165), .Z(N3166) );
  GTECH_AND2 C5743 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[109]), .Z(N3163) );
  GTECH_AND2 C5744 ( .A(N3164), .B(a2stg_shr[108]), .Z(N3165) );
  GTECH_AND2 C5745 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3164) );
  GTECH_AND2 C5746 ( .A(N3167), .B(a2stg_shr[108]), .Z(N3168) );
  GTECH_AND2 C5747 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3167) );
  GTECH_AND2 C5748 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3170) );
  GTECH_AND2 C5750 ( .A(N3172), .B(a3stg_frac2[56]), .Z(N3173) );
  GTECH_NOT I_499 ( .A(a6stg_step), .Z(N3172) );
  GTECH_NOT I_500 ( .A(N3186), .Z(a2stg_shr_frac2_inv[55]) );
  GTECH_OR2 C5753 ( .A(N3183), .B(N3185), .Z(N3186) );
  GTECH_OR2 C5754 ( .A(N3181), .B(N3182), .Z(N3183) );
  GTECH_OR2 C5755 ( .A(N3178), .B(N3180), .Z(N3181) );
  GTECH_OR2 C5756 ( .A(N3175), .B(N3177), .Z(N3178) );
  GTECH_AND2 C5757 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[108]), .Z(N3175) );
  GTECH_AND2 C5758 ( .A(N3176), .B(a2stg_shr[107]), .Z(N3177) );
  GTECH_AND2 C5759 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3176) );
  GTECH_AND2 C5760 ( .A(N3179), .B(a2stg_shr[107]), .Z(N3180) );
  GTECH_AND2 C5761 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3179) );
  GTECH_AND2 C5762 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3182) );
  GTECH_AND2 C5764 ( .A(N3184), .B(a3stg_frac2[55]), .Z(N3185) );
  GTECH_NOT I_501 ( .A(a6stg_step), .Z(N3184) );
  GTECH_NOT I_502 ( .A(N3198), .Z(a2stg_shr_frac2_inv[54]) );
  GTECH_OR2 C5767 ( .A(N3195), .B(N3197), .Z(N3198) );
  GTECH_OR2 C5768 ( .A(N3193), .B(N3194), .Z(N3195) );
  GTECH_OR2 C5769 ( .A(N3190), .B(N3192), .Z(N3193) );
  GTECH_OR2 C5770 ( .A(N3187), .B(N3189), .Z(N3190) );
  GTECH_AND2 C5771 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[107]), .Z(N3187) );
  GTECH_AND2 C5772 ( .A(N3188), .B(a2stg_shr[106]), .Z(N3189) );
  GTECH_AND2 C5773 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3188) );
  GTECH_AND2 C5774 ( .A(N3191), .B(a2stg_shr[106]), .Z(N3192) );
  GTECH_AND2 C5775 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3191) );
  GTECH_AND2 C5776 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3194) );
  GTECH_AND2 C5778 ( .A(N3196), .B(a3stg_frac2[54]), .Z(N3197) );
  GTECH_NOT I_503 ( .A(a6stg_step), .Z(N3196) );
  GTECH_NOT I_504 ( .A(N3210), .Z(a2stg_shr_frac2_inv[53]) );
  GTECH_OR2 C5781 ( .A(N3207), .B(N3209), .Z(N3210) );
  GTECH_OR2 C5782 ( .A(N3205), .B(N3206), .Z(N3207) );
  GTECH_OR2 C5783 ( .A(N3202), .B(N3204), .Z(N3205) );
  GTECH_OR2 C5784 ( .A(N3199), .B(N3201), .Z(N3202) );
  GTECH_AND2 C5785 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[106]), .Z(N3199) );
  GTECH_AND2 C5786 ( .A(N3200), .B(a2stg_shr[105]), .Z(N3201) );
  GTECH_AND2 C5787 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3200) );
  GTECH_AND2 C5788 ( .A(N3203), .B(a2stg_shr[105]), .Z(N3204) );
  GTECH_AND2 C5789 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3203) );
  GTECH_AND2 C5790 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3206) );
  GTECH_AND2 C5792 ( .A(N3208), .B(a3stg_frac2[53]), .Z(N3209) );
  GTECH_NOT I_505 ( .A(a6stg_step), .Z(N3208) );
  GTECH_NOT I_506 ( .A(N3222), .Z(a2stg_shr_frac2_inv[52]) );
  GTECH_OR2 C5795 ( .A(N3219), .B(N3221), .Z(N3222) );
  GTECH_OR2 C5796 ( .A(N3217), .B(N3218), .Z(N3219) );
  GTECH_OR2 C5797 ( .A(N3214), .B(N3216), .Z(N3217) );
  GTECH_OR2 C5798 ( .A(N3211), .B(N3213), .Z(N3214) );
  GTECH_AND2 C5799 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[105]), .Z(N3211) );
  GTECH_AND2 C5800 ( .A(N3212), .B(a2stg_shr[104]), .Z(N3213) );
  GTECH_AND2 C5801 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3212) );
  GTECH_AND2 C5802 ( .A(N3215), .B(a2stg_shr[104]), .Z(N3216) );
  GTECH_AND2 C5803 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3215) );
  GTECH_AND2 C5804 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3218) );
  GTECH_AND2 C5806 ( .A(N3220), .B(a3stg_frac2[52]), .Z(N3221) );
  GTECH_NOT I_507 ( .A(a6stg_step), .Z(N3220) );
  GTECH_NOT I_508 ( .A(N3234), .Z(a2stg_shr_frac2_inv[51]) );
  GTECH_OR2 C5809 ( .A(N3231), .B(N3233), .Z(N3234) );
  GTECH_OR2 C5810 ( .A(N3229), .B(N3230), .Z(N3231) );
  GTECH_OR2 C5811 ( .A(N3226), .B(N3228), .Z(N3229) );
  GTECH_OR2 C5812 ( .A(N3223), .B(N3225), .Z(N3226) );
  GTECH_AND2 C5813 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[104]), .Z(N3223) );
  GTECH_AND2 C5814 ( .A(N3224), .B(a2stg_shr[103]), .Z(N3225) );
  GTECH_AND2 C5815 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3224) );
  GTECH_AND2 C5816 ( .A(N3227), .B(a2stg_shr[103]), .Z(N3228) );
  GTECH_AND2 C5817 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3227) );
  GTECH_AND2 C5818 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3230) );
  GTECH_AND2 C5820 ( .A(N3232), .B(a3stg_frac2[51]), .Z(N3233) );
  GTECH_NOT I_509 ( .A(a6stg_step), .Z(N3232) );
  GTECH_NOT I_510 ( .A(N3246), .Z(a2stg_shr_frac2_inv[50]) );
  GTECH_OR2 C5823 ( .A(N3243), .B(N3245), .Z(N3246) );
  GTECH_OR2 C5824 ( .A(N3241), .B(N3242), .Z(N3243) );
  GTECH_OR2 C5825 ( .A(N3238), .B(N3240), .Z(N3241) );
  GTECH_OR2 C5826 ( .A(N3235), .B(N3237), .Z(N3238) );
  GTECH_AND2 C5827 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[103]), .Z(N3235) );
  GTECH_AND2 C5828 ( .A(N3236), .B(a2stg_shr[102]), .Z(N3237) );
  GTECH_AND2 C5829 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3236) );
  GTECH_AND2 C5830 ( .A(N3239), .B(a2stg_shr[102]), .Z(N3240) );
  GTECH_AND2 C5831 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3239) );
  GTECH_AND2 C5832 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3242) );
  GTECH_AND2 C5834 ( .A(N3244), .B(a3stg_frac2[50]), .Z(N3245) );
  GTECH_NOT I_511 ( .A(a6stg_step), .Z(N3244) );
  GTECH_NOT I_512 ( .A(N3258), .Z(a2stg_shr_frac2_inv[49]) );
  GTECH_OR2 C5837 ( .A(N3255), .B(N3257), .Z(N3258) );
  GTECH_OR2 C5838 ( .A(N3253), .B(N3254), .Z(N3255) );
  GTECH_OR2 C5839 ( .A(N3250), .B(N3252), .Z(N3253) );
  GTECH_OR2 C5840 ( .A(N3247), .B(N3249), .Z(N3250) );
  GTECH_AND2 C5841 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[102]), .Z(N3247) );
  GTECH_AND2 C5842 ( .A(N3248), .B(a2stg_shr[101]), .Z(N3249) );
  GTECH_AND2 C5843 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3248) );
  GTECH_AND2 C5844 ( .A(N3251), .B(a2stg_shr[101]), .Z(N3252) );
  GTECH_AND2 C5845 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3251) );
  GTECH_AND2 C5846 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3254) );
  GTECH_AND2 C5848 ( .A(N3256), .B(a3stg_frac2[49]), .Z(N3257) );
  GTECH_NOT I_513 ( .A(a6stg_step), .Z(N3256) );
  GTECH_NOT I_514 ( .A(N3270), .Z(a2stg_shr_frac2_inv[48]) );
  GTECH_OR2 C5851 ( .A(N3267), .B(N3269), .Z(N3270) );
  GTECH_OR2 C5852 ( .A(N3265), .B(N3266), .Z(N3267) );
  GTECH_OR2 C5853 ( .A(N3262), .B(N3264), .Z(N3265) );
  GTECH_OR2 C5854 ( .A(N3259), .B(N3261), .Z(N3262) );
  GTECH_AND2 C5855 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[101]), .Z(N3259) );
  GTECH_AND2 C5856 ( .A(N3260), .B(a2stg_shr[100]), .Z(N3261) );
  GTECH_AND2 C5857 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3260) );
  GTECH_AND2 C5858 ( .A(N3263), .B(a2stg_shr[100]), .Z(N3264) );
  GTECH_AND2 C5859 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3263) );
  GTECH_AND2 C5860 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3266) );
  GTECH_AND2 C5862 ( .A(N3268), .B(a3stg_frac2[48]), .Z(N3269) );
  GTECH_NOT I_515 ( .A(a6stg_step), .Z(N3268) );
  GTECH_NOT I_516 ( .A(N3282), .Z(a2stg_shr_frac2_inv[47]) );
  GTECH_OR2 C5865 ( .A(N3279), .B(N3281), .Z(N3282) );
  GTECH_OR2 C5866 ( .A(N3277), .B(N3278), .Z(N3279) );
  GTECH_OR2 C5867 ( .A(N3274), .B(N3276), .Z(N3277) );
  GTECH_OR2 C5868 ( .A(N3271), .B(N3273), .Z(N3274) );
  GTECH_AND2 C5869 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[100]), .Z(N3271) );
  GTECH_AND2 C5870 ( .A(N3272), .B(a2stg_shr[99]), .Z(N3273) );
  GTECH_AND2 C5871 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3272) );
  GTECH_AND2 C5872 ( .A(N3275), .B(a2stg_shr[99]), .Z(N3276) );
  GTECH_AND2 C5873 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3275) );
  GTECH_AND2 C5874 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3278) );
  GTECH_AND2 C5876 ( .A(N3280), .B(a3stg_frac2[47]), .Z(N3281) );
  GTECH_NOT I_517 ( .A(a6stg_step), .Z(N3280) );
  GTECH_NOT I_518 ( .A(N3294), .Z(a2stg_shr_frac2_inv[46]) );
  GTECH_OR2 C5879 ( .A(N3291), .B(N3293), .Z(N3294) );
  GTECH_OR2 C5880 ( .A(N3289), .B(N3290), .Z(N3291) );
  GTECH_OR2 C5881 ( .A(N3286), .B(N3288), .Z(N3289) );
  GTECH_OR2 C5882 ( .A(N3283), .B(N3285), .Z(N3286) );
  GTECH_AND2 C5883 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[99]), .Z(N3283)
         );
  GTECH_AND2 C5884 ( .A(N3284), .B(a2stg_shr[98]), .Z(N3285) );
  GTECH_AND2 C5885 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3284) );
  GTECH_AND2 C5886 ( .A(N3287), .B(a2stg_shr[98]), .Z(N3288) );
  GTECH_AND2 C5887 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3287) );
  GTECH_AND2 C5888 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3290) );
  GTECH_AND2 C5890 ( .A(N3292), .B(a3stg_frac2[46]), .Z(N3293) );
  GTECH_NOT I_519 ( .A(a6stg_step), .Z(N3292) );
  GTECH_NOT I_520 ( .A(N3306), .Z(a2stg_shr_frac2_inv[45]) );
  GTECH_OR2 C5893 ( .A(N3303), .B(N3305), .Z(N3306) );
  GTECH_OR2 C5894 ( .A(N3301), .B(N3302), .Z(N3303) );
  GTECH_OR2 C5895 ( .A(N3298), .B(N3300), .Z(N3301) );
  GTECH_OR2 C5896 ( .A(N3295), .B(N3297), .Z(N3298) );
  GTECH_AND2 C5897 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[98]), .Z(N3295)
         );
  GTECH_AND2 C5898 ( .A(N3296), .B(a2stg_shr[97]), .Z(N3297) );
  GTECH_AND2 C5899 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3296) );
  GTECH_AND2 C5900 ( .A(N3299), .B(a2stg_shr[97]), .Z(N3300) );
  GTECH_AND2 C5901 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3299) );
  GTECH_AND2 C5902 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3302) );
  GTECH_AND2 C5904 ( .A(N3304), .B(a3stg_frac2[45]), .Z(N3305) );
  GTECH_NOT I_521 ( .A(a6stg_step), .Z(N3304) );
  GTECH_NOT I_522 ( .A(N3318), .Z(a2stg_shr_frac2_inv[44]) );
  GTECH_OR2 C5907 ( .A(N3315), .B(N3317), .Z(N3318) );
  GTECH_OR2 C5908 ( .A(N3313), .B(N3314), .Z(N3315) );
  GTECH_OR2 C5909 ( .A(N3310), .B(N3312), .Z(N3313) );
  GTECH_OR2 C5910 ( .A(N3307), .B(N3309), .Z(N3310) );
  GTECH_AND2 C5911 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[97]), .Z(N3307)
         );
  GTECH_AND2 C5912 ( .A(N3308), .B(a2stg_shr[96]), .Z(N3309) );
  GTECH_AND2 C5913 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3308) );
  GTECH_AND2 C5914 ( .A(N3311), .B(a2stg_shr[96]), .Z(N3312) );
  GTECH_AND2 C5915 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3311) );
  GTECH_AND2 C5916 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3314) );
  GTECH_AND2 C5918 ( .A(N3316), .B(a3stg_frac2[44]), .Z(N3317) );
  GTECH_NOT I_523 ( .A(a6stg_step), .Z(N3316) );
  GTECH_NOT I_524 ( .A(N3330), .Z(a2stg_shr_frac2_inv[43]) );
  GTECH_OR2 C5921 ( .A(N3327), .B(N3329), .Z(N3330) );
  GTECH_OR2 C5922 ( .A(N3325), .B(N3326), .Z(N3327) );
  GTECH_OR2 C5923 ( .A(N3322), .B(N3324), .Z(N3325) );
  GTECH_OR2 C5924 ( .A(N3319), .B(N3321), .Z(N3322) );
  GTECH_AND2 C5925 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[96]), .Z(N3319)
         );
  GTECH_AND2 C5926 ( .A(N3320), .B(a2stg_shr[95]), .Z(N3321) );
  GTECH_AND2 C5927 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3320) );
  GTECH_AND2 C5928 ( .A(N3323), .B(a2stg_shr[95]), .Z(N3324) );
  GTECH_AND2 C5929 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3323) );
  GTECH_AND2 C5930 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3326) );
  GTECH_AND2 C5932 ( .A(N3328), .B(a3stg_frac2[43]), .Z(N3329) );
  GTECH_NOT I_525 ( .A(a6stg_step), .Z(N3328) );
  GTECH_NOT I_526 ( .A(N3342), .Z(a2stg_shr_frac2_inv[42]) );
  GTECH_OR2 C5935 ( .A(N3339), .B(N3341), .Z(N3342) );
  GTECH_OR2 C5936 ( .A(N3337), .B(N3338), .Z(N3339) );
  GTECH_OR2 C5937 ( .A(N3334), .B(N3336), .Z(N3337) );
  GTECH_OR2 C5938 ( .A(N3331), .B(N3333), .Z(N3334) );
  GTECH_AND2 C5939 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[95]), .Z(N3331)
         );
  GTECH_AND2 C5940 ( .A(N3332), .B(a2stg_shr[94]), .Z(N3333) );
  GTECH_AND2 C5941 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3332) );
  GTECH_AND2 C5942 ( .A(N3335), .B(a2stg_shr[94]), .Z(N3336) );
  GTECH_AND2 C5943 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3335) );
  GTECH_AND2 C5944 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3338) );
  GTECH_AND2 C5946 ( .A(N3340), .B(a3stg_frac2[42]), .Z(N3341) );
  GTECH_NOT I_527 ( .A(a6stg_step), .Z(N3340) );
  GTECH_NOT I_528 ( .A(N3354), .Z(a2stg_shr_frac2_inv[41]) );
  GTECH_OR2 C5949 ( .A(N3351), .B(N3353), .Z(N3354) );
  GTECH_OR2 C5950 ( .A(N3349), .B(N3350), .Z(N3351) );
  GTECH_OR2 C5951 ( .A(N3346), .B(N3348), .Z(N3349) );
  GTECH_OR2 C5952 ( .A(N3343), .B(N3345), .Z(N3346) );
  GTECH_AND2 C5953 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[94]), .Z(N3343)
         );
  GTECH_AND2 C5954 ( .A(N3344), .B(a2stg_shr[93]), .Z(N3345) );
  GTECH_AND2 C5955 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3344) );
  GTECH_AND2 C5956 ( .A(N3347), .B(a2stg_shr[93]), .Z(N3348) );
  GTECH_AND2 C5957 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3347) );
  GTECH_AND2 C5958 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3350) );
  GTECH_AND2 C5960 ( .A(N3352), .B(a3stg_frac2[41]), .Z(N3353) );
  GTECH_NOT I_529 ( .A(a6stg_step), .Z(N3352) );
  GTECH_NOT I_530 ( .A(N3366), .Z(a2stg_shr_frac2_inv[40]) );
  GTECH_OR2 C5963 ( .A(N3363), .B(N3365), .Z(N3366) );
  GTECH_OR2 C5964 ( .A(N3361), .B(N3362), .Z(N3363) );
  GTECH_OR2 C5965 ( .A(N3358), .B(N3360), .Z(N3361) );
  GTECH_OR2 C5966 ( .A(N3355), .B(N3357), .Z(N3358) );
  GTECH_AND2 C5967 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[93]), .Z(N3355)
         );
  GTECH_AND2 C5968 ( .A(N3356), .B(a2stg_shr[92]), .Z(N3357) );
  GTECH_AND2 C5969 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3356) );
  GTECH_AND2 C5970 ( .A(N3359), .B(a2stg_shr[92]), .Z(N3360) );
  GTECH_AND2 C5971 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3359) );
  GTECH_AND2 C5972 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3362) );
  GTECH_AND2 C5974 ( .A(N3364), .B(a3stg_frac2[40]), .Z(N3365) );
  GTECH_NOT I_531 ( .A(a6stg_step), .Z(N3364) );
  GTECH_NOT I_532 ( .A(N3378), .Z(a2stg_shr_frac2_inv[39]) );
  GTECH_OR2 C5977 ( .A(N3375), .B(N3377), .Z(N3378) );
  GTECH_OR2 C5978 ( .A(N3373), .B(N3374), .Z(N3375) );
  GTECH_OR2 C5979 ( .A(N3370), .B(N3372), .Z(N3373) );
  GTECH_OR2 C5980 ( .A(N3367), .B(N3369), .Z(N3370) );
  GTECH_AND2 C5981 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[92]), .Z(N3367)
         );
  GTECH_AND2 C5982 ( .A(N3368), .B(a2stg_shr[91]), .Z(N3369) );
  GTECH_AND2 C5983 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3368) );
  GTECH_AND2 C5984 ( .A(N3371), .B(a2stg_shr[91]), .Z(N3372) );
  GTECH_AND2 C5985 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3371) );
  GTECH_AND2 C5986 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3374) );
  GTECH_AND2 C5988 ( .A(N3376), .B(a3stg_frac2[39]), .Z(N3377) );
  GTECH_NOT I_533 ( .A(a6stg_step), .Z(N3376) );
  GTECH_NOT I_534 ( .A(N3390), .Z(a2stg_shr_frac2_inv[38]) );
  GTECH_OR2 C5991 ( .A(N3387), .B(N3389), .Z(N3390) );
  GTECH_OR2 C5992 ( .A(N3385), .B(N3386), .Z(N3387) );
  GTECH_OR2 C5993 ( .A(N3382), .B(N3384), .Z(N3385) );
  GTECH_OR2 C5994 ( .A(N3379), .B(N3381), .Z(N3382) );
  GTECH_AND2 C5995 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[91]), .Z(N3379)
         );
  GTECH_AND2 C5996 ( .A(N3380), .B(a2stg_shr[90]), .Z(N3381) );
  GTECH_AND2 C5997 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3380) );
  GTECH_AND2 C5998 ( .A(N3383), .B(a2stg_shr[90]), .Z(N3384) );
  GTECH_AND2 C5999 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3383) );
  GTECH_AND2 C6000 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3386) );
  GTECH_AND2 C6002 ( .A(N3388), .B(a3stg_frac2[38]), .Z(N3389) );
  GTECH_NOT I_535 ( .A(a6stg_step), .Z(N3388) );
  GTECH_NOT I_536 ( .A(N3402), .Z(a2stg_shr_frac2_inv[37]) );
  GTECH_OR2 C6005 ( .A(N3399), .B(N3401), .Z(N3402) );
  GTECH_OR2 C6006 ( .A(N3397), .B(N3398), .Z(N3399) );
  GTECH_OR2 C6007 ( .A(N3394), .B(N3396), .Z(N3397) );
  GTECH_OR2 C6008 ( .A(N3391), .B(N3393), .Z(N3394) );
  GTECH_AND2 C6009 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[90]), .Z(N3391)
         );
  GTECH_AND2 C6010 ( .A(N3392), .B(a2stg_shr[89]), .Z(N3393) );
  GTECH_AND2 C6011 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3392) );
  GTECH_AND2 C6012 ( .A(N3395), .B(a2stg_shr[89]), .Z(N3396) );
  GTECH_AND2 C6013 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3395) );
  GTECH_AND2 C6014 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3398) );
  GTECH_AND2 C6016 ( .A(N3400), .B(a3stg_frac2[37]), .Z(N3401) );
  GTECH_NOT I_537 ( .A(a6stg_step), .Z(N3400) );
  GTECH_NOT I_538 ( .A(N3414), .Z(a2stg_shr_frac2_inv[36]) );
  GTECH_OR2 C6019 ( .A(N3411), .B(N3413), .Z(N3414) );
  GTECH_OR2 C6020 ( .A(N3409), .B(N3410), .Z(N3411) );
  GTECH_OR2 C6021 ( .A(N3406), .B(N3408), .Z(N3409) );
  GTECH_OR2 C6022 ( .A(N3403), .B(N3405), .Z(N3406) );
  GTECH_AND2 C6023 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[89]), .Z(N3403)
         );
  GTECH_AND2 C6024 ( .A(N3404), .B(a2stg_shr[88]), .Z(N3405) );
  GTECH_AND2 C6025 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3404) );
  GTECH_AND2 C6026 ( .A(N3407), .B(a2stg_shr[88]), .Z(N3408) );
  GTECH_AND2 C6027 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3407) );
  GTECH_AND2 C6028 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3410) );
  GTECH_AND2 C6030 ( .A(N3412), .B(a3stg_frac2[36]), .Z(N3413) );
  GTECH_NOT I_539 ( .A(a6stg_step), .Z(N3412) );
  GTECH_NOT I_540 ( .A(N3426), .Z(a2stg_shr_frac2_inv[35]) );
  GTECH_OR2 C6033 ( .A(N3423), .B(N3425), .Z(N3426) );
  GTECH_OR2 C6034 ( .A(N3421), .B(N3422), .Z(N3423) );
  GTECH_OR2 C6035 ( .A(N3418), .B(N3420), .Z(N3421) );
  GTECH_OR2 C6036 ( .A(N3415), .B(N3417), .Z(N3418) );
  GTECH_AND2 C6037 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[88]), .Z(N3415)
         );
  GTECH_AND2 C6038 ( .A(N3416), .B(a2stg_shr[87]), .Z(N3417) );
  GTECH_AND2 C6039 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3416) );
  GTECH_AND2 C6040 ( .A(N3419), .B(a2stg_shr[87]), .Z(N3420) );
  GTECH_AND2 C6041 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3419) );
  GTECH_AND2 C6042 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3422) );
  GTECH_AND2 C6044 ( .A(N3424), .B(a3stg_frac2[35]), .Z(N3425) );
  GTECH_NOT I_541 ( .A(a6stg_step), .Z(N3424) );
  GTECH_NOT I_542 ( .A(N3438), .Z(a2stg_shr_frac2_inv[34]) );
  GTECH_OR2 C6047 ( .A(N3435), .B(N3437), .Z(N3438) );
  GTECH_OR2 C6048 ( .A(N3433), .B(N3434), .Z(N3435) );
  GTECH_OR2 C6049 ( .A(N3430), .B(N3432), .Z(N3433) );
  GTECH_OR2 C6050 ( .A(N3427), .B(N3429), .Z(N3430) );
  GTECH_AND2 C6051 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[87]), .Z(N3427)
         );
  GTECH_AND2 C6052 ( .A(N3428), .B(a2stg_shr[86]), .Z(N3429) );
  GTECH_AND2 C6053 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3428) );
  GTECH_AND2 C6054 ( .A(N3431), .B(a2stg_shr[86]), .Z(N3432) );
  GTECH_AND2 C6055 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3431) );
  GTECH_AND2 C6056 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3434) );
  GTECH_AND2 C6058 ( .A(N3436), .B(a3stg_frac2[34]), .Z(N3437) );
  GTECH_NOT I_543 ( .A(a6stg_step), .Z(N3436) );
  GTECH_NOT I_544 ( .A(N3450), .Z(a2stg_shr_frac2_inv[33]) );
  GTECH_OR2 C6061 ( .A(N3447), .B(N3449), .Z(N3450) );
  GTECH_OR2 C6062 ( .A(N3445), .B(N3446), .Z(N3447) );
  GTECH_OR2 C6063 ( .A(N3442), .B(N3444), .Z(N3445) );
  GTECH_OR2 C6064 ( .A(N3439), .B(N3441), .Z(N3442) );
  GTECH_AND2 C6065 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[86]), .Z(N3439)
         );
  GTECH_AND2 C6066 ( .A(N3440), .B(a2stg_shr[85]), .Z(N3441) );
  GTECH_AND2 C6067 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3440) );
  GTECH_AND2 C6068 ( .A(N3443), .B(a2stg_shr[85]), .Z(N3444) );
  GTECH_AND2 C6069 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3443) );
  GTECH_AND2 C6070 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3446) );
  GTECH_AND2 C6072 ( .A(N3448), .B(a3stg_frac2[33]), .Z(N3449) );
  GTECH_NOT I_545 ( .A(a6stg_step), .Z(N3448) );
  GTECH_NOT I_546 ( .A(N3462), .Z(a2stg_shr_frac2_inv[32]) );
  GTECH_OR2 C6075 ( .A(N3459), .B(N3461), .Z(N3462) );
  GTECH_OR2 C6076 ( .A(N3457), .B(N3458), .Z(N3459) );
  GTECH_OR2 C6077 ( .A(N3454), .B(N3456), .Z(N3457) );
  GTECH_OR2 C6078 ( .A(N3451), .B(N3453), .Z(N3454) );
  GTECH_AND2 C6079 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[85]), .Z(N3451)
         );
  GTECH_AND2 C6080 ( .A(N3452), .B(a2stg_shr[84]), .Z(N3453) );
  GTECH_AND2 C6081 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3452) );
  GTECH_AND2 C6082 ( .A(N3455), .B(a2stg_shr[84]), .Z(N3456) );
  GTECH_AND2 C6083 ( .A(a2stg_shr_frac2_shr_sng), .B(a2stg_expadd_11), .Z(
        N3455) );
  GTECH_AND2 C6084 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3458) );
  GTECH_AND2 C6086 ( .A(N3460), .B(a3stg_frac2[32]), .Z(N3461) );
  GTECH_NOT I_547 ( .A(a6stg_step), .Z(N3460) );
  GTECH_NOT I_548 ( .A(N3471), .Z(a2stg_shr_frac2_inv[31]) );
  GTECH_OR2 C6089 ( .A(N3468), .B(N3470), .Z(N3471) );
  GTECH_OR2 C6090 ( .A(N3466), .B(N3467), .Z(N3468) );
  GTECH_OR2 C6091 ( .A(N3463), .B(N3465), .Z(N3466) );
  GTECH_AND2 C6092 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[84]), .Z(N3463)
         );
  GTECH_AND2 C6093 ( .A(N3464), .B(a2stg_shr[83]), .Z(N3465) );
  GTECH_AND2 C6094 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3464) );
  GTECH_AND2 C6095 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3467) );
  GTECH_AND2 C6097 ( .A(N3469), .B(a3stg_frac2[31]), .Z(N3470) );
  GTECH_NOT I_549 ( .A(a6stg_step), .Z(N3469) );
  GTECH_NOT I_550 ( .A(N3480), .Z(a2stg_shr_frac2_inv[30]) );
  GTECH_OR2 C6100 ( .A(N3477), .B(N3479), .Z(N3480) );
  GTECH_OR2 C6101 ( .A(N3475), .B(N3476), .Z(N3477) );
  GTECH_OR2 C6102 ( .A(N3472), .B(N3474), .Z(N3475) );
  GTECH_AND2 C6103 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[83]), .Z(N3472)
         );
  GTECH_AND2 C6104 ( .A(N3473), .B(a2stg_shr[82]), .Z(N3474) );
  GTECH_AND2 C6105 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3473) );
  GTECH_AND2 C6106 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3476) );
  GTECH_AND2 C6108 ( .A(N3478), .B(a3stg_frac2[30]), .Z(N3479) );
  GTECH_NOT I_551 ( .A(a6stg_step), .Z(N3478) );
  GTECH_NOT I_552 ( .A(N3489), .Z(a2stg_shr_frac2_inv[29]) );
  GTECH_OR2 C6111 ( .A(N3486), .B(N3488), .Z(N3489) );
  GTECH_OR2 C6112 ( .A(N3484), .B(N3485), .Z(N3486) );
  GTECH_OR2 C6113 ( .A(N3481), .B(N3483), .Z(N3484) );
  GTECH_AND2 C6114 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[82]), .Z(N3481)
         );
  GTECH_AND2 C6115 ( .A(N3482), .B(a2stg_shr[81]), .Z(N3483) );
  GTECH_AND2 C6116 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3482) );
  GTECH_AND2 C6117 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3485) );
  GTECH_AND2 C6119 ( .A(N3487), .B(a3stg_frac2[29]), .Z(N3488) );
  GTECH_NOT I_553 ( .A(a6stg_step), .Z(N3487) );
  GTECH_NOT I_554 ( .A(N3498), .Z(a2stg_shr_frac2_inv[28]) );
  GTECH_OR2 C6122 ( .A(N3495), .B(N3497), .Z(N3498) );
  GTECH_OR2 C6123 ( .A(N3493), .B(N3494), .Z(N3495) );
  GTECH_OR2 C6124 ( .A(N3490), .B(N3492), .Z(N3493) );
  GTECH_AND2 C6125 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[81]), .Z(N3490)
         );
  GTECH_AND2 C6126 ( .A(N3491), .B(a2stg_shr[80]), .Z(N3492) );
  GTECH_AND2 C6127 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3491) );
  GTECH_AND2 C6128 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3494) );
  GTECH_AND2 C6130 ( .A(N3496), .B(a3stg_frac2[28]), .Z(N3497) );
  GTECH_NOT I_555 ( .A(a6stg_step), .Z(N3496) );
  GTECH_NOT I_556 ( .A(N3507), .Z(a2stg_shr_frac2_inv[27]) );
  GTECH_OR2 C6133 ( .A(N3504), .B(N3506), .Z(N3507) );
  GTECH_OR2 C6134 ( .A(N3502), .B(N3503), .Z(N3504) );
  GTECH_OR2 C6135 ( .A(N3499), .B(N3501), .Z(N3502) );
  GTECH_AND2 C6136 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[80]), .Z(N3499)
         );
  GTECH_AND2 C6137 ( .A(N3500), .B(a2stg_shr[79]), .Z(N3501) );
  GTECH_AND2 C6138 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3500) );
  GTECH_AND2 C6139 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3503) );
  GTECH_AND2 C6141 ( .A(N3505), .B(a3stg_frac2[27]), .Z(N3506) );
  GTECH_NOT I_557 ( .A(a6stg_step), .Z(N3505) );
  GTECH_NOT I_558 ( .A(N3516), .Z(a2stg_shr_frac2_inv[26]) );
  GTECH_OR2 C6144 ( .A(N3513), .B(N3515), .Z(N3516) );
  GTECH_OR2 C6145 ( .A(N3511), .B(N3512), .Z(N3513) );
  GTECH_OR2 C6146 ( .A(N3508), .B(N3510), .Z(N3511) );
  GTECH_AND2 C6147 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[79]), .Z(N3508)
         );
  GTECH_AND2 C6148 ( .A(N3509), .B(a2stg_shr[78]), .Z(N3510) );
  GTECH_AND2 C6149 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3509) );
  GTECH_AND2 C6150 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3512) );
  GTECH_AND2 C6152 ( .A(N3514), .B(a3stg_frac2[26]), .Z(N3515) );
  GTECH_NOT I_559 ( .A(a6stg_step), .Z(N3514) );
  GTECH_NOT I_560 ( .A(N3525), .Z(a2stg_shr_frac2_inv[25]) );
  GTECH_OR2 C6155 ( .A(N3522), .B(N3524), .Z(N3525) );
  GTECH_OR2 C6156 ( .A(N3520), .B(N3521), .Z(N3522) );
  GTECH_OR2 C6157 ( .A(N3517), .B(N3519), .Z(N3520) );
  GTECH_AND2 C6158 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[78]), .Z(N3517)
         );
  GTECH_AND2 C6159 ( .A(N3518), .B(a2stg_shr[77]), .Z(N3519) );
  GTECH_AND2 C6160 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3518) );
  GTECH_AND2 C6161 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3521) );
  GTECH_AND2 C6163 ( .A(N3523), .B(a3stg_frac2[25]), .Z(N3524) );
  GTECH_NOT I_561 ( .A(a6stg_step), .Z(N3523) );
  GTECH_NOT I_562 ( .A(N3534), .Z(a2stg_shr_frac2_inv[24]) );
  GTECH_OR2 C6166 ( .A(N3531), .B(N3533), .Z(N3534) );
  GTECH_OR2 C6167 ( .A(N3529), .B(N3530), .Z(N3531) );
  GTECH_OR2 C6168 ( .A(N3526), .B(N3528), .Z(N3529) );
  GTECH_AND2 C6169 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[77]), .Z(N3526)
         );
  GTECH_AND2 C6170 ( .A(N3527), .B(a2stg_shr[76]), .Z(N3528) );
  GTECH_AND2 C6171 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3527) );
  GTECH_AND2 C6172 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3530) );
  GTECH_AND2 C6174 ( .A(N3532), .B(a3stg_frac2[24]), .Z(N3533) );
  GTECH_NOT I_563 ( .A(a6stg_step), .Z(N3532) );
  GTECH_NOT I_564 ( .A(N3543), .Z(a2stg_shr_frac2_inv[23]) );
  GTECH_OR2 C6177 ( .A(N3540), .B(N3542), .Z(N3543) );
  GTECH_OR2 C6178 ( .A(N3538), .B(N3539), .Z(N3540) );
  GTECH_OR2 C6179 ( .A(N3535), .B(N3537), .Z(N3538) );
  GTECH_AND2 C6180 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[76]), .Z(N3535)
         );
  GTECH_AND2 C6181 ( .A(N3536), .B(a2stg_shr[75]), .Z(N3537) );
  GTECH_AND2 C6182 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3536) );
  GTECH_AND2 C6183 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3539) );
  GTECH_AND2 C6185 ( .A(N3541), .B(a3stg_frac2[23]), .Z(N3542) );
  GTECH_NOT I_565 ( .A(a6stg_step), .Z(N3541) );
  GTECH_NOT I_566 ( .A(N3552), .Z(a2stg_shr_frac2_inv[22]) );
  GTECH_OR2 C6188 ( .A(N3549), .B(N3551), .Z(N3552) );
  GTECH_OR2 C6189 ( .A(N3547), .B(N3548), .Z(N3549) );
  GTECH_OR2 C6190 ( .A(N3544), .B(N3546), .Z(N3547) );
  GTECH_AND2 C6191 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[75]), .Z(N3544)
         );
  GTECH_AND2 C6192 ( .A(N3545), .B(a2stg_shr[74]), .Z(N3546) );
  GTECH_AND2 C6193 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3545) );
  GTECH_AND2 C6194 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3548) );
  GTECH_AND2 C6196 ( .A(N3550), .B(a3stg_frac2[22]), .Z(N3551) );
  GTECH_NOT I_567 ( .A(a6stg_step), .Z(N3550) );
  GTECH_NOT I_568 ( .A(N3561), .Z(a2stg_shr_frac2_inv[21]) );
  GTECH_OR2 C6199 ( .A(N3558), .B(N3560), .Z(N3561) );
  GTECH_OR2 C6200 ( .A(N3556), .B(N3557), .Z(N3558) );
  GTECH_OR2 C6201 ( .A(N3553), .B(N3555), .Z(N3556) );
  GTECH_AND2 C6202 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[74]), .Z(N3553)
         );
  GTECH_AND2 C6203 ( .A(N3554), .B(a2stg_shr[73]), .Z(N3555) );
  GTECH_AND2 C6204 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3554) );
  GTECH_AND2 C6205 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3557) );
  GTECH_AND2 C6207 ( .A(N3559), .B(a3stg_frac2[21]), .Z(N3560) );
  GTECH_NOT I_569 ( .A(a6stg_step), .Z(N3559) );
  GTECH_NOT I_570 ( .A(N3570), .Z(a2stg_shr_frac2_inv[20]) );
  GTECH_OR2 C6210 ( .A(N3567), .B(N3569), .Z(N3570) );
  GTECH_OR2 C6211 ( .A(N3565), .B(N3566), .Z(N3567) );
  GTECH_OR2 C6212 ( .A(N3562), .B(N3564), .Z(N3565) );
  GTECH_AND2 C6213 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[73]), .Z(N3562)
         );
  GTECH_AND2 C6214 ( .A(N3563), .B(a2stg_shr[72]), .Z(N3564) );
  GTECH_AND2 C6215 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3563) );
  GTECH_AND2 C6216 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3566) );
  GTECH_AND2 C6218 ( .A(N3568), .B(a3stg_frac2[20]), .Z(N3569) );
  GTECH_NOT I_571 ( .A(a6stg_step), .Z(N3568) );
  GTECH_NOT I_572 ( .A(N3579), .Z(a2stg_shr_frac2_inv[19]) );
  GTECH_OR2 C6221 ( .A(N3576), .B(N3578), .Z(N3579) );
  GTECH_OR2 C6222 ( .A(N3574), .B(N3575), .Z(N3576) );
  GTECH_OR2 C6223 ( .A(N3571), .B(N3573), .Z(N3574) );
  GTECH_AND2 C6224 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[72]), .Z(N3571)
         );
  GTECH_AND2 C6225 ( .A(N3572), .B(a2stg_shr[71]), .Z(N3573) );
  GTECH_AND2 C6226 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3572) );
  GTECH_AND2 C6227 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3575) );
  GTECH_AND2 C6229 ( .A(N3577), .B(a3stg_frac2[19]), .Z(N3578) );
  GTECH_NOT I_573 ( .A(a6stg_step), .Z(N3577) );
  GTECH_NOT I_574 ( .A(N3588), .Z(a2stg_shr_frac2_inv[18]) );
  GTECH_OR2 C6232 ( .A(N3585), .B(N3587), .Z(N3588) );
  GTECH_OR2 C6233 ( .A(N3583), .B(N3584), .Z(N3585) );
  GTECH_OR2 C6234 ( .A(N3580), .B(N3582), .Z(N3583) );
  GTECH_AND2 C6235 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[71]), .Z(N3580)
         );
  GTECH_AND2 C6236 ( .A(N3581), .B(a2stg_shr[70]), .Z(N3582) );
  GTECH_AND2 C6237 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3581) );
  GTECH_AND2 C6238 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3584) );
  GTECH_AND2 C6240 ( .A(N3586), .B(a3stg_frac2[18]), .Z(N3587) );
  GTECH_NOT I_575 ( .A(a6stg_step), .Z(N3586) );
  GTECH_NOT I_576 ( .A(N3597), .Z(a2stg_shr_frac2_inv[17]) );
  GTECH_OR2 C6243 ( .A(N3594), .B(N3596), .Z(N3597) );
  GTECH_OR2 C6244 ( .A(N3592), .B(N3593), .Z(N3594) );
  GTECH_OR2 C6245 ( .A(N3589), .B(N3591), .Z(N3592) );
  GTECH_AND2 C6246 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[70]), .Z(N3589)
         );
  GTECH_AND2 C6247 ( .A(N3590), .B(a2stg_shr[69]), .Z(N3591) );
  GTECH_AND2 C6248 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3590) );
  GTECH_AND2 C6249 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3593) );
  GTECH_AND2 C6251 ( .A(N3595), .B(a3stg_frac2[17]), .Z(N3596) );
  GTECH_NOT I_577 ( .A(a6stg_step), .Z(N3595) );
  GTECH_NOT I_578 ( .A(N3606), .Z(a2stg_shr_frac2_inv[16]) );
  GTECH_OR2 C6254 ( .A(N3603), .B(N3605), .Z(N3606) );
  GTECH_OR2 C6255 ( .A(N3601), .B(N3602), .Z(N3603) );
  GTECH_OR2 C6256 ( .A(N3598), .B(N3600), .Z(N3601) );
  GTECH_AND2 C6257 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[69]), .Z(N3598)
         );
  GTECH_AND2 C6258 ( .A(N3599), .B(a2stg_shr[68]), .Z(N3600) );
  GTECH_AND2 C6259 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3599) );
  GTECH_AND2 C6260 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3602) );
  GTECH_AND2 C6262 ( .A(N3604), .B(a3stg_frac2[16]), .Z(N3605) );
  GTECH_NOT I_579 ( .A(a6stg_step), .Z(N3604) );
  GTECH_NOT I_580 ( .A(N3615), .Z(a2stg_shr_frac2_inv[15]) );
  GTECH_OR2 C6265 ( .A(N3612), .B(N3614), .Z(N3615) );
  GTECH_OR2 C6266 ( .A(N3610), .B(N3611), .Z(N3612) );
  GTECH_OR2 C6267 ( .A(N3607), .B(N3609), .Z(N3610) );
  GTECH_AND2 C6268 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[68]), .Z(N3607)
         );
  GTECH_AND2 C6269 ( .A(N3608), .B(a2stg_shr[67]), .Z(N3609) );
  GTECH_AND2 C6270 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3608) );
  GTECH_AND2 C6271 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3611) );
  GTECH_AND2 C6273 ( .A(N3613), .B(a3stg_frac2[15]), .Z(N3614) );
  GTECH_NOT I_581 ( .A(a6stg_step), .Z(N3613) );
  GTECH_NOT I_582 ( .A(N3624), .Z(a2stg_shr_frac2_inv[14]) );
  GTECH_OR2 C6276 ( .A(N3621), .B(N3623), .Z(N3624) );
  GTECH_OR2 C6277 ( .A(N3619), .B(N3620), .Z(N3621) );
  GTECH_OR2 C6278 ( .A(N3616), .B(N3618), .Z(N3619) );
  GTECH_AND2 C6279 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[67]), .Z(N3616)
         );
  GTECH_AND2 C6280 ( .A(N3617), .B(a2stg_shr[66]), .Z(N3618) );
  GTECH_AND2 C6281 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3617) );
  GTECH_AND2 C6282 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3620) );
  GTECH_AND2 C6284 ( .A(N3622), .B(a3stg_frac2[14]), .Z(N3623) );
  GTECH_NOT I_583 ( .A(a6stg_step), .Z(N3622) );
  GTECH_NOT I_584 ( .A(N3633), .Z(a2stg_shr_frac2_inv[13]) );
  GTECH_OR2 C6287 ( .A(N3630), .B(N3632), .Z(N3633) );
  GTECH_OR2 C6288 ( .A(N3628), .B(N3629), .Z(N3630) );
  GTECH_OR2 C6289 ( .A(N3625), .B(N3627), .Z(N3628) );
  GTECH_AND2 C6290 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[66]), .Z(N3625)
         );
  GTECH_AND2 C6291 ( .A(N3626), .B(a2stg_shr[65]), .Z(N3627) );
  GTECH_AND2 C6292 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3626) );
  GTECH_AND2 C6293 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3629) );
  GTECH_AND2 C6295 ( .A(N3631), .B(a3stg_frac2[13]), .Z(N3632) );
  GTECH_NOT I_585 ( .A(a6stg_step), .Z(N3631) );
  GTECH_NOT I_586 ( .A(N3642), .Z(a2stg_shr_frac2_inv[12]) );
  GTECH_OR2 C6298 ( .A(N3639), .B(N3641), .Z(N3642) );
  GTECH_OR2 C6299 ( .A(N3637), .B(N3638), .Z(N3639) );
  GTECH_OR2 C6300 ( .A(N3634), .B(N3636), .Z(N3637) );
  GTECH_AND2 C6301 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[65]), .Z(N3634)
         );
  GTECH_AND2 C6302 ( .A(N3635), .B(a2stg_shr[64]), .Z(N3636) );
  GTECH_AND2 C6303 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3635) );
  GTECH_AND2 C6304 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3638) );
  GTECH_AND2 C6306 ( .A(N3640), .B(a3stg_frac2[12]), .Z(N3641) );
  GTECH_NOT I_587 ( .A(a6stg_step), .Z(N3640) );
  GTECH_NOT I_588 ( .A(N3651), .Z(a2stg_shr_frac2_inv[11]) );
  GTECH_OR2 C6309 ( .A(N3648), .B(N3650), .Z(N3651) );
  GTECH_OR2 C6310 ( .A(N3646), .B(N3647), .Z(N3648) );
  GTECH_OR2 C6311 ( .A(N3643), .B(N3645), .Z(N3646) );
  GTECH_AND2 C6312 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[64]), .Z(N3643)
         );
  GTECH_AND2 C6313 ( .A(N3644), .B(a2stg_shr[63]), .Z(N3645) );
  GTECH_AND2 C6314 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3644) );
  GTECH_AND2 C6315 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3647) );
  GTECH_AND2 C6317 ( .A(N3649), .B(a3stg_frac2[11]), .Z(N3650) );
  GTECH_NOT I_589 ( .A(a6stg_step), .Z(N3649) );
  GTECH_NOT I_590 ( .A(N3660), .Z(a2stg_shr_frac2_inv[10]) );
  GTECH_OR2 C6320 ( .A(N3657), .B(N3659), .Z(N3660) );
  GTECH_OR2 C6321 ( .A(N3655), .B(N3656), .Z(N3657) );
  GTECH_OR2 C6322 ( .A(N3652), .B(N3654), .Z(N3655) );
  GTECH_AND2 C6323 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[63]), .Z(N3652)
         );
  GTECH_AND2 C6324 ( .A(N3653), .B(a2stg_shr[62]), .Z(N3654) );
  GTECH_AND2 C6325 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3653) );
  GTECH_AND2 C6326 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3656) );
  GTECH_AND2 C6328 ( .A(N3658), .B(a3stg_frac2[10]), .Z(N3659) );
  GTECH_NOT I_591 ( .A(a6stg_step), .Z(N3658) );
  GTECH_NOT I_592 ( .A(N3669), .Z(a2stg_shr_frac2_inv[9]) );
  GTECH_OR2 C6331 ( .A(N3666), .B(N3668), .Z(N3669) );
  GTECH_OR2 C6332 ( .A(N3664), .B(N3665), .Z(N3666) );
  GTECH_OR2 C6333 ( .A(N3661), .B(N3663), .Z(N3664) );
  GTECH_AND2 C6334 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[62]), .Z(N3661)
         );
  GTECH_AND2 C6335 ( .A(N3662), .B(a2stg_shr[61]), .Z(N3663) );
  GTECH_AND2 C6336 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3662) );
  GTECH_AND2 C6337 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3665) );
  GTECH_AND2 C6339 ( .A(N3667), .B(a3stg_frac2[9]), .Z(N3668) );
  GTECH_NOT I_593 ( .A(a6stg_step), .Z(N3667) );
  GTECH_NOT I_594 ( .A(N3678), .Z(a2stg_shr_frac2_inv[8]) );
  GTECH_OR2 C6342 ( .A(N3675), .B(N3677), .Z(N3678) );
  GTECH_OR2 C6343 ( .A(N3673), .B(N3674), .Z(N3675) );
  GTECH_OR2 C6344 ( .A(N3670), .B(N3672), .Z(N3673) );
  GTECH_AND2 C6345 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr[61]), .Z(N3670)
         );
  GTECH_AND2 C6346 ( .A(N3671), .B(a2stg_shr[60]), .Z(N3672) );
  GTECH_AND2 C6347 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3671) );
  GTECH_AND2 C6348 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3674) );
  GTECH_AND2 C6350 ( .A(N3676), .B(a3stg_frac2[8]), .Z(N3677) );
  GTECH_NOT I_595 ( .A(a6stg_step), .Z(N3676) );
  GTECH_NOT I_596 ( .A(N3687), .Z(a2stg_shr_frac2_inv[7]) );
  GTECH_OR2 C6353 ( .A(N3684), .B(N3686), .Z(N3687) );
  GTECH_OR2 C6354 ( .A(N3682), .B(N3683), .Z(N3684) );
  GTECH_OR2 C6355 ( .A(N3679), .B(N3681), .Z(N3682) );
  GTECH_AND2 C6356 ( .A(a2stg_shr_frac2_shr_int), .B(a2stg_shr_60_0_neq_0), 
        .Z(N3679) );
  GTECH_AND2 C6357 ( .A(N3680), .B(a2stg_shr[59]), .Z(N3681) );
  GTECH_AND2 C6358 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3680) );
  GTECH_AND2 C6359 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3683) );
  GTECH_AND2 C6361 ( .A(N3685), .B(a3stg_frac2[7]), .Z(N3686) );
  GTECH_NOT I_597 ( .A(a6stg_step), .Z(N3685) );
  GTECH_NOT I_598 ( .A(N3694), .Z(a2stg_shr_frac2_inv[6]) );
  GTECH_OR2 C6364 ( .A(N3691), .B(N3693), .Z(N3694) );
  GTECH_OR2 C6365 ( .A(N3689), .B(N3690), .Z(N3691) );
  GTECH_AND2 C6366 ( .A(N3688), .B(a2stg_shr[58]), .Z(N3689) );
  GTECH_AND2 C6367 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3688) );
  GTECH_AND2 C6368 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3690) );
  GTECH_AND2 C6370 ( .A(N3692), .B(a3stg_frac2[6]), .Z(N3693) );
  GTECH_NOT I_599 ( .A(a6stg_step), .Z(N3692) );
  GTECH_NOT I_600 ( .A(N3701), .Z(a2stg_shr_frac2_inv[5]) );
  GTECH_OR2 C6373 ( .A(N3698), .B(N3700), .Z(N3701) );
  GTECH_OR2 C6374 ( .A(N3696), .B(N3697), .Z(N3698) );
  GTECH_AND2 C6375 ( .A(N3695), .B(a2stg_shr[57]), .Z(N3696) );
  GTECH_AND2 C6376 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3695) );
  GTECH_AND2 C6377 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3697) );
  GTECH_AND2 C6379 ( .A(N3699), .B(a3stg_frac2[5]), .Z(N3700) );
  GTECH_NOT I_601 ( .A(a6stg_step), .Z(N3699) );
  GTECH_NOT I_602 ( .A(N3708), .Z(a2stg_shr_frac2_inv[4]) );
  GTECH_OR2 C6382 ( .A(N3705), .B(N3707), .Z(N3708) );
  GTECH_OR2 C6383 ( .A(N3703), .B(N3704), .Z(N3705) );
  GTECH_AND2 C6384 ( .A(N3702), .B(a2stg_shr[56]), .Z(N3703) );
  GTECH_AND2 C6385 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3702) );
  GTECH_AND2 C6386 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3704) );
  GTECH_AND2 C6388 ( .A(N3706), .B(a3stg_frac2[4]), .Z(N3707) );
  GTECH_NOT I_603 ( .A(a6stg_step), .Z(N3706) );
  GTECH_NOT I_604 ( .A(N3715), .Z(a2stg_shr_frac2_inv[3]) );
  GTECH_OR2 C6391 ( .A(N3712), .B(N3714), .Z(N3715) );
  GTECH_OR2 C6392 ( .A(N3710), .B(N3711), .Z(N3712) );
  GTECH_AND2 C6393 ( .A(N3709), .B(a2stg_shr[55]), .Z(N3710) );
  GTECH_AND2 C6394 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3709) );
  GTECH_AND2 C6395 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3711) );
  GTECH_AND2 C6397 ( .A(N3713), .B(a3stg_frac2[3]), .Z(N3714) );
  GTECH_NOT I_605 ( .A(a6stg_step), .Z(N3713) );
  GTECH_NOT I_606 ( .A(N3722), .Z(a2stg_shr_frac2_inv[2]) );
  GTECH_OR2 C6400 ( .A(N3719), .B(N3721), .Z(N3722) );
  GTECH_OR2 C6401 ( .A(N3717), .B(N3718), .Z(N3719) );
  GTECH_AND2 C6402 ( .A(N3716), .B(a2stg_shr[54]), .Z(N3717) );
  GTECH_AND2 C6403 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3716) );
  GTECH_AND2 C6404 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3718) );
  GTECH_AND2 C6406 ( .A(N3720), .B(a3stg_frac2[2]), .Z(N3721) );
  GTECH_NOT I_607 ( .A(a6stg_step), .Z(N3720) );
  GTECH_NOT I_608 ( .A(N3729), .Z(a2stg_shr_frac2_inv[1]) );
  GTECH_OR2 C6409 ( .A(N3726), .B(N3728), .Z(N3729) );
  GTECH_OR2 C6410 ( .A(N3724), .B(N3725), .Z(N3726) );
  GTECH_AND2 C6411 ( .A(N3723), .B(a2stg_shr[53]), .Z(N3724) );
  GTECH_AND2 C6412 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3723) );
  GTECH_AND2 C6413 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3725) );
  GTECH_AND2 C6415 ( .A(N3727), .B(a3stg_frac2[1]), .Z(N3728) );
  GTECH_NOT I_609 ( .A(a6stg_step), .Z(N3727) );
  GTECH_NOT I_610 ( .A(N3736), .Z(a2stg_shr_frac2_inv[0]) );
  GTECH_OR2 C6418 ( .A(N3733), .B(N3735), .Z(N3736) );
  GTECH_OR2 C6419 ( .A(N3731), .B(N3732), .Z(N3733) );
  GTECH_AND2 C6420 ( .A(N3730), .B(a2stg_shr[52]), .Z(N3731) );
  GTECH_AND2 C6421 ( .A(a2stg_shr_frac2_shr_dbl), .B(a2stg_expadd_11), .Z(
        N3730) );
  GTECH_AND2 C6422 ( .A(a2stg_shr_frac2_max), .B(N3097), .Z(N3732) );
  GTECH_AND2 C6424 ( .A(N3734), .B(a3stg_frac2[0]), .Z(N3735) );
  GTECH_NOT I_611 ( .A(a6stg_step), .Z(N3734) );
  GTECH_NOT I_612 ( .A(N3737), .Z(a3stg_frac2_in[63]) );
  GTECH_XOR2 C6427 ( .A(a2stg_shr_frac2_inv[63]), .B(a2stg_sub_step), .Z(N3737) );
  GTECH_NOT I_613 ( .A(N3738), .Z(a3stg_frac2_in[62]) );
  GTECH_XOR2 C6429 ( .A(a2stg_shr_frac2_inv[62]), .B(a2stg_sub_step), .Z(N3738) );
  GTECH_NOT I_614 ( .A(N3739), .Z(a3stg_frac2_in[61]) );
  GTECH_XOR2 C6431 ( .A(a2stg_shr_frac2_inv[61]), .B(a2stg_sub_step), .Z(N3739) );
  GTECH_NOT I_615 ( .A(N3740), .Z(a3stg_frac2_in[60]) );
  GTECH_XOR2 C6433 ( .A(a2stg_shr_frac2_inv[60]), .B(a2stg_sub_step), .Z(N3740) );
  GTECH_NOT I_616 ( .A(N3741), .Z(a3stg_frac2_in[59]) );
  GTECH_XOR2 C6435 ( .A(a2stg_shr_frac2_inv[59]), .B(a2stg_sub_step), .Z(N3741) );
  GTECH_NOT I_617 ( .A(N3742), .Z(a3stg_frac2_in[58]) );
  GTECH_XOR2 C6437 ( .A(a2stg_shr_frac2_inv[58]), .B(a2stg_sub_step), .Z(N3742) );
  GTECH_NOT I_618 ( .A(N3743), .Z(a3stg_frac2_in[57]) );
  GTECH_XOR2 C6439 ( .A(a2stg_shr_frac2_inv[57]), .B(a2stg_sub_step), .Z(N3743) );
  GTECH_NOT I_619 ( .A(N3744), .Z(a3stg_frac2_in[56]) );
  GTECH_XOR2 C6441 ( .A(a2stg_shr_frac2_inv[56]), .B(a2stg_sub_step), .Z(N3744) );
  GTECH_NOT I_620 ( .A(N3745), .Z(a3stg_frac2_in[55]) );
  GTECH_XOR2 C6443 ( .A(a2stg_shr_frac2_inv[55]), .B(a2stg_sub_step), .Z(N3745) );
  GTECH_NOT I_621 ( .A(N3746), .Z(a3stg_frac2_in[54]) );
  GTECH_XOR2 C6445 ( .A(a2stg_shr_frac2_inv[54]), .B(a2stg_sub_step), .Z(N3746) );
  GTECH_NOT I_622 ( .A(N3747), .Z(a3stg_frac2_in[53]) );
  GTECH_XOR2 C6447 ( .A(a2stg_shr_frac2_inv[53]), .B(a2stg_sub_step), .Z(N3747) );
  GTECH_NOT I_623 ( .A(N3748), .Z(a3stg_frac2_in[52]) );
  GTECH_XOR2 C6449 ( .A(a2stg_shr_frac2_inv[52]), .B(a2stg_sub_step), .Z(N3748) );
  GTECH_NOT I_624 ( .A(N3749), .Z(a3stg_frac2_in[51]) );
  GTECH_XOR2 C6451 ( .A(a2stg_shr_frac2_inv[51]), .B(a2stg_sub_step), .Z(N3749) );
  GTECH_NOT I_625 ( .A(N3750), .Z(a3stg_frac2_in[50]) );
  GTECH_XOR2 C6453 ( .A(a2stg_shr_frac2_inv[50]), .B(a2stg_sub_step), .Z(N3750) );
  GTECH_NOT I_626 ( .A(N3751), .Z(a3stg_frac2_in[49]) );
  GTECH_XOR2 C6455 ( .A(a2stg_shr_frac2_inv[49]), .B(a2stg_sub_step), .Z(N3751) );
  GTECH_NOT I_627 ( .A(N3752), .Z(a3stg_frac2_in[48]) );
  GTECH_XOR2 C6457 ( .A(a2stg_shr_frac2_inv[48]), .B(a2stg_sub_step), .Z(N3752) );
  GTECH_NOT I_628 ( .A(N3753), .Z(a3stg_frac2_in[47]) );
  GTECH_XOR2 C6459 ( .A(a2stg_shr_frac2_inv[47]), .B(a2stg_sub_step), .Z(N3753) );
  GTECH_NOT I_629 ( .A(N3754), .Z(a3stg_frac2_in[46]) );
  GTECH_XOR2 C6461 ( .A(a2stg_shr_frac2_inv[46]), .B(a2stg_sub_step), .Z(N3754) );
  GTECH_NOT I_630 ( .A(N3755), .Z(a3stg_frac2_in[45]) );
  GTECH_XOR2 C6463 ( .A(a2stg_shr_frac2_inv[45]), .B(a2stg_sub_step), .Z(N3755) );
  GTECH_NOT I_631 ( .A(N3756), .Z(a3stg_frac2_in[44]) );
  GTECH_XOR2 C6465 ( .A(a2stg_shr_frac2_inv[44]), .B(a2stg_sub_step), .Z(N3756) );
  GTECH_NOT I_632 ( .A(N3757), .Z(a3stg_frac2_in[43]) );
  GTECH_XOR2 C6467 ( .A(a2stg_shr_frac2_inv[43]), .B(a2stg_sub_step), .Z(N3757) );
  GTECH_NOT I_633 ( .A(N3758), .Z(a3stg_frac2_in[42]) );
  GTECH_XOR2 C6469 ( .A(a2stg_shr_frac2_inv[42]), .B(a2stg_sub_step), .Z(N3758) );
  GTECH_NOT I_634 ( .A(N3759), .Z(a3stg_frac2_in[41]) );
  GTECH_XOR2 C6471 ( .A(a2stg_shr_frac2_inv[41]), .B(a2stg_sub_step), .Z(N3759) );
  GTECH_NOT I_635 ( .A(N3760), .Z(a3stg_frac2_in[40]) );
  GTECH_XOR2 C6473 ( .A(a2stg_shr_frac2_inv[40]), .B(a2stg_sub_step), .Z(N3760) );
  GTECH_NOT I_636 ( .A(N3761), .Z(a3stg_frac2_in[39]) );
  GTECH_XOR2 C6475 ( .A(a2stg_shr_frac2_inv[39]), .B(a2stg_sub_step), .Z(N3761) );
  GTECH_NOT I_637 ( .A(N3762), .Z(a3stg_frac2_in[38]) );
  GTECH_XOR2 C6477 ( .A(a2stg_shr_frac2_inv[38]), .B(a2stg_sub_step), .Z(N3762) );
  GTECH_NOT I_638 ( .A(N3763), .Z(a3stg_frac2_in[37]) );
  GTECH_XOR2 C6479 ( .A(a2stg_shr_frac2_inv[37]), .B(a2stg_sub_step), .Z(N3763) );
  GTECH_NOT I_639 ( .A(N3764), .Z(a3stg_frac2_in[36]) );
  GTECH_XOR2 C6481 ( .A(a2stg_shr_frac2_inv[36]), .B(a2stg_sub_step), .Z(N3764) );
  GTECH_NOT I_640 ( .A(N3765), .Z(a3stg_frac2_in[35]) );
  GTECH_XOR2 C6483 ( .A(a2stg_shr_frac2_inv[35]), .B(a2stg_sub_step), .Z(N3765) );
  GTECH_NOT I_641 ( .A(N3766), .Z(a3stg_frac2_in[34]) );
  GTECH_XOR2 C6485 ( .A(a2stg_shr_frac2_inv[34]), .B(a2stg_sub_step), .Z(N3766) );
  GTECH_NOT I_642 ( .A(N3767), .Z(a3stg_frac2_in[33]) );
  GTECH_XOR2 C6487 ( .A(a2stg_shr_frac2_inv[33]), .B(a2stg_sub_step), .Z(N3767) );
  GTECH_NOT I_643 ( .A(N3768), .Z(a3stg_frac2_in[32]) );
  GTECH_XOR2 C6489 ( .A(a2stg_shr_frac2_inv[32]), .B(a2stg_sub_step), .Z(N3768) );
  GTECH_NOT I_644 ( .A(N3769), .Z(a3stg_frac2_in[31]) );
  GTECH_XOR2 C6491 ( .A(a2stg_shr_frac2_inv[31]), .B(a2stg_sub_step), .Z(N3769) );
  GTECH_NOT I_645 ( .A(N3770), .Z(a3stg_frac2_in[30]) );
  GTECH_XOR2 C6493 ( .A(a2stg_shr_frac2_inv[30]), .B(a2stg_sub_step), .Z(N3770) );
  GTECH_NOT I_646 ( .A(N3771), .Z(a3stg_frac2_in[29]) );
  GTECH_XOR2 C6495 ( .A(a2stg_shr_frac2_inv[29]), .B(a2stg_sub_step), .Z(N3771) );
  GTECH_NOT I_647 ( .A(N3772), .Z(a3stg_frac2_in[28]) );
  GTECH_XOR2 C6497 ( .A(a2stg_shr_frac2_inv[28]), .B(a2stg_sub_step), .Z(N3772) );
  GTECH_NOT I_648 ( .A(N3773), .Z(a3stg_frac2_in[27]) );
  GTECH_XOR2 C6499 ( .A(a2stg_shr_frac2_inv[27]), .B(a2stg_sub_step), .Z(N3773) );
  GTECH_NOT I_649 ( .A(N3774), .Z(a3stg_frac2_in[26]) );
  GTECH_XOR2 C6501 ( .A(a2stg_shr_frac2_inv[26]), .B(a2stg_sub_step), .Z(N3774) );
  GTECH_NOT I_650 ( .A(N3775), .Z(a3stg_frac2_in[25]) );
  GTECH_XOR2 C6503 ( .A(a2stg_shr_frac2_inv[25]), .B(a2stg_sub_step), .Z(N3775) );
  GTECH_NOT I_651 ( .A(N3776), .Z(a3stg_frac2_in[24]) );
  GTECH_XOR2 C6505 ( .A(a2stg_shr_frac2_inv[24]), .B(a2stg_sub_step), .Z(N3776) );
  GTECH_NOT I_652 ( .A(N3777), .Z(a3stg_frac2_in[23]) );
  GTECH_XOR2 C6507 ( .A(a2stg_shr_frac2_inv[23]), .B(a2stg_sub_step), .Z(N3777) );
  GTECH_NOT I_653 ( .A(N3778), .Z(a3stg_frac2_in[22]) );
  GTECH_XOR2 C6509 ( .A(a2stg_shr_frac2_inv[22]), .B(a2stg_sub_step), .Z(N3778) );
  GTECH_NOT I_654 ( .A(N3779), .Z(a3stg_frac2_in[21]) );
  GTECH_XOR2 C6511 ( .A(a2stg_shr_frac2_inv[21]), .B(a2stg_sub_step), .Z(N3779) );
  GTECH_NOT I_655 ( .A(N3780), .Z(a3stg_frac2_in[20]) );
  GTECH_XOR2 C6513 ( .A(a2stg_shr_frac2_inv[20]), .B(a2stg_sub_step), .Z(N3780) );
  GTECH_NOT I_656 ( .A(N3781), .Z(a3stg_frac2_in[19]) );
  GTECH_XOR2 C6515 ( .A(a2stg_shr_frac2_inv[19]), .B(a2stg_sub_step), .Z(N3781) );
  GTECH_NOT I_657 ( .A(N3782), .Z(a3stg_frac2_in[18]) );
  GTECH_XOR2 C6517 ( .A(a2stg_shr_frac2_inv[18]), .B(a2stg_sub_step), .Z(N3782) );
  GTECH_NOT I_658 ( .A(N3783), .Z(a3stg_frac2_in[17]) );
  GTECH_XOR2 C6519 ( .A(a2stg_shr_frac2_inv[17]), .B(a2stg_sub_step), .Z(N3783) );
  GTECH_NOT I_659 ( .A(N3784), .Z(a3stg_frac2_in[16]) );
  GTECH_XOR2 C6521 ( .A(a2stg_shr_frac2_inv[16]), .B(a2stg_sub_step), .Z(N3784) );
  GTECH_NOT I_660 ( .A(N3785), .Z(a3stg_frac2_in[15]) );
  GTECH_XOR2 C6523 ( .A(a2stg_shr_frac2_inv[15]), .B(a2stg_sub_step), .Z(N3785) );
  GTECH_NOT I_661 ( .A(N3786), .Z(a3stg_frac2_in[14]) );
  GTECH_XOR2 C6525 ( .A(a2stg_shr_frac2_inv[14]), .B(a2stg_sub_step), .Z(N3786) );
  GTECH_NOT I_662 ( .A(N3787), .Z(a3stg_frac2_in[13]) );
  GTECH_XOR2 C6527 ( .A(a2stg_shr_frac2_inv[13]), .B(a2stg_sub_step), .Z(N3787) );
  GTECH_NOT I_663 ( .A(N3788), .Z(a3stg_frac2_in[12]) );
  GTECH_XOR2 C6529 ( .A(a2stg_shr_frac2_inv[12]), .B(a2stg_sub_step), .Z(N3788) );
  GTECH_NOT I_664 ( .A(N3789), .Z(a3stg_frac2_in[11]) );
  GTECH_XOR2 C6531 ( .A(a2stg_shr_frac2_inv[11]), .B(a2stg_sub_step), .Z(N3789) );
  GTECH_NOT I_665 ( .A(N3790), .Z(a3stg_frac2_in[10]) );
  GTECH_XOR2 C6533 ( .A(a2stg_shr_frac2_inv[10]), .B(a2stg_sub_step), .Z(N3790) );
  GTECH_NOT I_666 ( .A(N3791), .Z(a3stg_frac2_in[9]) );
  GTECH_XOR2 C6535 ( .A(a2stg_shr_frac2_inv[9]), .B(a2stg_sub_step), .Z(N3791)
         );
  GTECH_NOT I_667 ( .A(N3792), .Z(a3stg_frac2_in[8]) );
  GTECH_XOR2 C6537 ( .A(a2stg_shr_frac2_inv[8]), .B(a2stg_sub_step), .Z(N3792)
         );
  GTECH_NOT I_668 ( .A(N3793), .Z(a3stg_frac2_in[7]) );
  GTECH_XOR2 C6539 ( .A(a2stg_shr_frac2_inv[7]), .B(a2stg_sub_step), .Z(N3793)
         );
  GTECH_NOT I_669 ( .A(N3794), .Z(a3stg_frac2_in[6]) );
  GTECH_XOR2 C6541 ( .A(a2stg_shr_frac2_inv[6]), .B(a2stg_sub_step), .Z(N3794)
         );
  GTECH_NOT I_670 ( .A(N3795), .Z(a3stg_frac2_in[5]) );
  GTECH_XOR2 C6543 ( .A(a2stg_shr_frac2_inv[5]), .B(a2stg_sub_step), .Z(N3795)
         );
  GTECH_NOT I_671 ( .A(N3796), .Z(a3stg_frac2_in[4]) );
  GTECH_XOR2 C6545 ( .A(a2stg_shr_frac2_inv[4]), .B(a2stg_sub_step), .Z(N3796)
         );
  GTECH_NOT I_672 ( .A(N3797), .Z(a3stg_frac2_in[3]) );
  GTECH_XOR2 C6547 ( .A(a2stg_shr_frac2_inv[3]), .B(a2stg_sub_step), .Z(N3797)
         );
  GTECH_NOT I_673 ( .A(N3798), .Z(a3stg_frac2_in[2]) );
  GTECH_XOR2 C6549 ( .A(a2stg_shr_frac2_inv[2]), .B(a2stg_sub_step), .Z(N3798)
         );
  GTECH_NOT I_674 ( .A(N3799), .Z(a3stg_frac2_in[1]) );
  GTECH_XOR2 C6551 ( .A(a2stg_shr_frac2_inv[1]), .B(a2stg_sub_step), .Z(N3799)
         );
  GTECH_NOT I_675 ( .A(N3800), .Z(a3stg_frac2_in[0]) );
  GTECH_XOR2 C6553 ( .A(a2stg_shr_frac2_inv[0]), .B(a2stg_sub_step), .Z(N3800)
         );
  GTECH_OR2 C6554 ( .A(N3803), .B(N3804), .Z(a2stg_fracadd_in2[63]) );
  GTECH_OR2 C6555 ( .A(N3802), .B(a2stg_fracadd_frac2_inv_shr1), .Z(N3803) );
  GTECH_AND2 C6556 ( .A(a2stg_fracadd_frac2_inv), .B(N3801), .Z(N3802) );
  GTECH_NOT I_676 ( .A(a2stg_frac2_63), .Z(N3801) );
  GTECH_AND2 C6558 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2_63), .Z(N3804) );
  GTECH_OR2 C6559 ( .A(N3808), .B(N3809), .Z(a2stg_fracadd_in2[62]) );
  GTECH_OR2 C6560 ( .A(N3806), .B(N3807), .Z(N3808) );
  GTECH_AND2 C6561 ( .A(a2stg_fracadd_frac2_inv), .B(N3805), .Z(N3806) );
  GTECH_NOT I_677 ( .A(a2stg_frac2[62]), .Z(N3805) );
  GTECH_AND2 C6563 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3801), .Z(N3807) );
  GTECH_AND2 C6565 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[62]), .Z(N3809)
         );
  GTECH_OR2 C6566 ( .A(N3813), .B(N3814), .Z(a2stg_fracadd_in2[61]) );
  GTECH_OR2 C6567 ( .A(N3811), .B(N3812), .Z(N3813) );
  GTECH_AND2 C6568 ( .A(a2stg_fracadd_frac2_inv), .B(N3810), .Z(N3811) );
  GTECH_NOT I_678 ( .A(a2stg_frac2[61]), .Z(N3810) );
  GTECH_AND2 C6570 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3805), .Z(N3812) );
  GTECH_AND2 C6572 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[61]), .Z(N3814)
         );
  GTECH_OR2 C6573 ( .A(N3818), .B(N3819), .Z(a2stg_fracadd_in2[60]) );
  GTECH_OR2 C6574 ( .A(N3816), .B(N3817), .Z(N3818) );
  GTECH_AND2 C6575 ( .A(a2stg_fracadd_frac2_inv), .B(N3815), .Z(N3816) );
  GTECH_NOT I_679 ( .A(a2stg_frac2[60]), .Z(N3815) );
  GTECH_AND2 C6577 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3810), .Z(N3817) );
  GTECH_AND2 C6579 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[60]), .Z(N3819)
         );
  GTECH_OR2 C6580 ( .A(N3823), .B(N3824), .Z(a2stg_fracadd_in2[59]) );
  GTECH_OR2 C6581 ( .A(N3821), .B(N3822), .Z(N3823) );
  GTECH_AND2 C6582 ( .A(a2stg_fracadd_frac2_inv), .B(N3820), .Z(N3821) );
  GTECH_NOT I_680 ( .A(a2stg_frac2[59]), .Z(N3820) );
  GTECH_AND2 C6584 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3815), .Z(N3822) );
  GTECH_AND2 C6586 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[59]), .Z(N3824)
         );
  GTECH_OR2 C6587 ( .A(N3828), .B(N3829), .Z(a2stg_fracadd_in2[58]) );
  GTECH_OR2 C6588 ( .A(N3826), .B(N3827), .Z(N3828) );
  GTECH_AND2 C6589 ( .A(a2stg_fracadd_frac2_inv), .B(N3825), .Z(N3826) );
  GTECH_NOT I_681 ( .A(a2stg_frac2[58]), .Z(N3825) );
  GTECH_AND2 C6591 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3820), .Z(N3827) );
  GTECH_AND2 C6593 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[58]), .Z(N3829)
         );
  GTECH_OR2 C6594 ( .A(N3833), .B(N3834), .Z(a2stg_fracadd_in2[57]) );
  GTECH_OR2 C6595 ( .A(N3831), .B(N3832), .Z(N3833) );
  GTECH_AND2 C6596 ( .A(a2stg_fracadd_frac2_inv), .B(N3830), .Z(N3831) );
  GTECH_NOT I_682 ( .A(a2stg_frac2[57]), .Z(N3830) );
  GTECH_AND2 C6598 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3825), .Z(N3832) );
  GTECH_AND2 C6600 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[57]), .Z(N3834)
         );
  GTECH_OR2 C6601 ( .A(N3838), .B(N3839), .Z(a2stg_fracadd_in2[56]) );
  GTECH_OR2 C6602 ( .A(N3836), .B(N3837), .Z(N3838) );
  GTECH_AND2 C6603 ( .A(a2stg_fracadd_frac2_inv), .B(N3835), .Z(N3836) );
  GTECH_NOT I_683 ( .A(a2stg_frac2[56]), .Z(N3835) );
  GTECH_AND2 C6605 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3830), .Z(N3837) );
  GTECH_AND2 C6607 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[56]), .Z(N3839)
         );
  GTECH_OR2 C6608 ( .A(N3843), .B(N3844), .Z(a2stg_fracadd_in2[55]) );
  GTECH_OR2 C6609 ( .A(N3841), .B(N3842), .Z(N3843) );
  GTECH_AND2 C6610 ( .A(a2stg_fracadd_frac2_inv), .B(N3840), .Z(N3841) );
  GTECH_NOT I_684 ( .A(a2stg_frac2[55]), .Z(N3840) );
  GTECH_AND2 C6612 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3835), .Z(N3842) );
  GTECH_AND2 C6614 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[55]), .Z(N3844)
         );
  GTECH_OR2 C6615 ( .A(N3848), .B(N3849), .Z(a2stg_fracadd_in2[54]) );
  GTECH_OR2 C6616 ( .A(N3846), .B(N3847), .Z(N3848) );
  GTECH_AND2 C6617 ( .A(a2stg_fracadd_frac2_inv), .B(N3845), .Z(N3846) );
  GTECH_NOT I_685 ( .A(a2stg_frac2[54]), .Z(N3845) );
  GTECH_AND2 C6619 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3840), .Z(N3847) );
  GTECH_AND2 C6621 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[54]), .Z(N3849)
         );
  GTECH_OR2 C6622 ( .A(N3853), .B(N3854), .Z(a2stg_fracadd_in2[53]) );
  GTECH_OR2 C6623 ( .A(N3851), .B(N3852), .Z(N3853) );
  GTECH_AND2 C6624 ( .A(a2stg_fracadd_frac2_inv), .B(N3850), .Z(N3851) );
  GTECH_NOT I_686 ( .A(a2stg_frac2[53]), .Z(N3850) );
  GTECH_AND2 C6626 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3845), .Z(N3852) );
  GTECH_AND2 C6628 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[53]), .Z(N3854)
         );
  GTECH_OR2 C6629 ( .A(N3858), .B(N3859), .Z(a2stg_fracadd_in2[52]) );
  GTECH_OR2 C6630 ( .A(N3856), .B(N3857), .Z(N3858) );
  GTECH_AND2 C6631 ( .A(a2stg_fracadd_frac2_inv), .B(N3855), .Z(N3856) );
  GTECH_NOT I_687 ( .A(a2stg_frac2[52]), .Z(N3855) );
  GTECH_AND2 C6633 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3850), .Z(N3857) );
  GTECH_AND2 C6635 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[52]), .Z(N3859)
         );
  GTECH_OR2 C6636 ( .A(N3863), .B(N3864), .Z(a2stg_fracadd_in2[51]) );
  GTECH_OR2 C6637 ( .A(N3861), .B(N3862), .Z(N3863) );
  GTECH_AND2 C6638 ( .A(a2stg_fracadd_frac2_inv), .B(N3860), .Z(N3861) );
  GTECH_NOT I_688 ( .A(a2stg_frac2[51]), .Z(N3860) );
  GTECH_AND2 C6640 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3855), .Z(N3862) );
  GTECH_AND2 C6642 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[51]), .Z(N3864)
         );
  GTECH_OR2 C6643 ( .A(N3868), .B(N3869), .Z(a2stg_fracadd_in2[50]) );
  GTECH_OR2 C6644 ( .A(N3866), .B(N3867), .Z(N3868) );
  GTECH_AND2 C6645 ( .A(a2stg_fracadd_frac2_inv), .B(N3865), .Z(N3866) );
  GTECH_NOT I_689 ( .A(a2stg_frac2[50]), .Z(N3865) );
  GTECH_AND2 C6647 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3860), .Z(N3867) );
  GTECH_AND2 C6649 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[50]), .Z(N3869)
         );
  GTECH_OR2 C6650 ( .A(N3873), .B(N3874), .Z(a2stg_fracadd_in2[49]) );
  GTECH_OR2 C6651 ( .A(N3871), .B(N3872), .Z(N3873) );
  GTECH_AND2 C6652 ( .A(a2stg_fracadd_frac2_inv), .B(N3870), .Z(N3871) );
  GTECH_NOT I_690 ( .A(a2stg_frac2[49]), .Z(N3870) );
  GTECH_AND2 C6654 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3865), .Z(N3872) );
  GTECH_AND2 C6656 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[49]), .Z(N3874)
         );
  GTECH_OR2 C6657 ( .A(N3878), .B(N3879), .Z(a2stg_fracadd_in2[48]) );
  GTECH_OR2 C6658 ( .A(N3876), .B(N3877), .Z(N3878) );
  GTECH_AND2 C6659 ( .A(a2stg_fracadd_frac2_inv), .B(N3875), .Z(N3876) );
  GTECH_NOT I_691 ( .A(a2stg_frac2[48]), .Z(N3875) );
  GTECH_AND2 C6661 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3870), .Z(N3877) );
  GTECH_AND2 C6663 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[48]), .Z(N3879)
         );
  GTECH_OR2 C6664 ( .A(N3883), .B(N3884), .Z(a2stg_fracadd_in2[47]) );
  GTECH_OR2 C6665 ( .A(N3881), .B(N3882), .Z(N3883) );
  GTECH_AND2 C6666 ( .A(a2stg_fracadd_frac2_inv), .B(N3880), .Z(N3881) );
  GTECH_NOT I_692 ( .A(a2stg_frac2[47]), .Z(N3880) );
  GTECH_AND2 C6668 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3875), .Z(N3882) );
  GTECH_AND2 C6670 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[47]), .Z(N3884)
         );
  GTECH_OR2 C6671 ( .A(N3888), .B(N3889), .Z(a2stg_fracadd_in2[46]) );
  GTECH_OR2 C6672 ( .A(N3886), .B(N3887), .Z(N3888) );
  GTECH_AND2 C6673 ( .A(a2stg_fracadd_frac2_inv), .B(N3885), .Z(N3886) );
  GTECH_NOT I_693 ( .A(a2stg_frac2[46]), .Z(N3885) );
  GTECH_AND2 C6675 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3880), .Z(N3887) );
  GTECH_AND2 C6677 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[46]), .Z(N3889)
         );
  GTECH_OR2 C6678 ( .A(N3893), .B(N3894), .Z(a2stg_fracadd_in2[45]) );
  GTECH_OR2 C6679 ( .A(N3891), .B(N3892), .Z(N3893) );
  GTECH_AND2 C6680 ( .A(a2stg_fracadd_frac2_inv), .B(N3890), .Z(N3891) );
  GTECH_NOT I_694 ( .A(a2stg_frac2[45]), .Z(N3890) );
  GTECH_AND2 C6682 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3885), .Z(N3892) );
  GTECH_AND2 C6684 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[45]), .Z(N3894)
         );
  GTECH_OR2 C6685 ( .A(N3898), .B(N3899), .Z(a2stg_fracadd_in2[44]) );
  GTECH_OR2 C6686 ( .A(N3896), .B(N3897), .Z(N3898) );
  GTECH_AND2 C6687 ( .A(a2stg_fracadd_frac2_inv), .B(N3895), .Z(N3896) );
  GTECH_NOT I_695 ( .A(a2stg_frac2[44]), .Z(N3895) );
  GTECH_AND2 C6689 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3890), .Z(N3897) );
  GTECH_AND2 C6691 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[44]), .Z(N3899)
         );
  GTECH_OR2 C6692 ( .A(N3903), .B(N3904), .Z(a2stg_fracadd_in2[43]) );
  GTECH_OR2 C6693 ( .A(N3901), .B(N3902), .Z(N3903) );
  GTECH_AND2 C6694 ( .A(a2stg_fracadd_frac2_inv), .B(N3900), .Z(N3901) );
  GTECH_NOT I_696 ( .A(a2stg_frac2[43]), .Z(N3900) );
  GTECH_AND2 C6696 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3895), .Z(N3902) );
  GTECH_AND2 C6698 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[43]), .Z(N3904)
         );
  GTECH_OR2 C6699 ( .A(N3908), .B(N3909), .Z(a2stg_fracadd_in2[42]) );
  GTECH_OR2 C6700 ( .A(N3906), .B(N3907), .Z(N3908) );
  GTECH_AND2 C6701 ( .A(a2stg_fracadd_frac2_inv), .B(N3905), .Z(N3906) );
  GTECH_NOT I_697 ( .A(a2stg_frac2[42]), .Z(N3905) );
  GTECH_AND2 C6703 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3900), .Z(N3907) );
  GTECH_AND2 C6705 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[42]), .Z(N3909)
         );
  GTECH_OR2 C6706 ( .A(N3913), .B(N3914), .Z(a2stg_fracadd_in2[41]) );
  GTECH_OR2 C6707 ( .A(N3911), .B(N3912), .Z(N3913) );
  GTECH_AND2 C6708 ( .A(a2stg_fracadd_frac2_inv), .B(N3910), .Z(N3911) );
  GTECH_NOT I_698 ( .A(a2stg_frac2[41]), .Z(N3910) );
  GTECH_AND2 C6710 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3905), .Z(N3912) );
  GTECH_AND2 C6712 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[41]), .Z(N3914)
         );
  GTECH_OR2 C6713 ( .A(N3918), .B(N3919), .Z(a2stg_fracadd_in2[40]) );
  GTECH_OR2 C6714 ( .A(N3916), .B(N3917), .Z(N3918) );
  GTECH_AND2 C6715 ( .A(a2stg_fracadd_frac2_inv), .B(N3915), .Z(N3916) );
  GTECH_NOT I_699 ( .A(a2stg_frac2[40]), .Z(N3915) );
  GTECH_AND2 C6717 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3910), .Z(N3917) );
  GTECH_AND2 C6719 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[40]), .Z(N3919)
         );
  GTECH_OR2 C6720 ( .A(N3923), .B(N3924), .Z(a2stg_fracadd_in2[39]) );
  GTECH_OR2 C6721 ( .A(N3921), .B(N3922), .Z(N3923) );
  GTECH_AND2 C6722 ( .A(a2stg_fracadd_frac2_inv), .B(N3920), .Z(N3921) );
  GTECH_NOT I_700 ( .A(a2stg_frac2[39]), .Z(N3920) );
  GTECH_AND2 C6724 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3915), .Z(N3922) );
  GTECH_AND2 C6726 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[39]), .Z(N3924)
         );
  GTECH_OR2 C6727 ( .A(N3928), .B(N3929), .Z(a2stg_fracadd_in2[38]) );
  GTECH_OR2 C6728 ( .A(N3926), .B(N3927), .Z(N3928) );
  GTECH_AND2 C6729 ( .A(a2stg_fracadd_frac2_inv), .B(N3925), .Z(N3926) );
  GTECH_NOT I_701 ( .A(a2stg_frac2[38]), .Z(N3925) );
  GTECH_AND2 C6731 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3920), .Z(N3927) );
  GTECH_AND2 C6733 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[38]), .Z(N3929)
         );
  GTECH_OR2 C6734 ( .A(N3933), .B(N3934), .Z(a2stg_fracadd_in2[37]) );
  GTECH_OR2 C6735 ( .A(N3931), .B(N3932), .Z(N3933) );
  GTECH_AND2 C6736 ( .A(a2stg_fracadd_frac2_inv), .B(N3930), .Z(N3931) );
  GTECH_NOT I_702 ( .A(a2stg_frac2[37]), .Z(N3930) );
  GTECH_AND2 C6738 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3925), .Z(N3932) );
  GTECH_AND2 C6740 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[37]), .Z(N3934)
         );
  GTECH_OR2 C6741 ( .A(N3938), .B(N3939), .Z(a2stg_fracadd_in2[36]) );
  GTECH_OR2 C6742 ( .A(N3936), .B(N3937), .Z(N3938) );
  GTECH_AND2 C6743 ( .A(a2stg_fracadd_frac2_inv), .B(N3935), .Z(N3936) );
  GTECH_NOT I_703 ( .A(a2stg_frac2[36]), .Z(N3935) );
  GTECH_AND2 C6745 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3930), .Z(N3937) );
  GTECH_AND2 C6747 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[36]), .Z(N3939)
         );
  GTECH_OR2 C6748 ( .A(N3943), .B(N3944), .Z(a2stg_fracadd_in2[35]) );
  GTECH_OR2 C6749 ( .A(N3941), .B(N3942), .Z(N3943) );
  GTECH_AND2 C6750 ( .A(a2stg_fracadd_frac2_inv), .B(N3940), .Z(N3941) );
  GTECH_NOT I_704 ( .A(a2stg_frac2[35]), .Z(N3940) );
  GTECH_AND2 C6752 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3935), .Z(N3942) );
  GTECH_AND2 C6754 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[35]), .Z(N3944)
         );
  GTECH_OR2 C6755 ( .A(N3948), .B(N3949), .Z(a2stg_fracadd_in2[34]) );
  GTECH_OR2 C6756 ( .A(N3946), .B(N3947), .Z(N3948) );
  GTECH_AND2 C6757 ( .A(a2stg_fracadd_frac2_inv), .B(N3945), .Z(N3946) );
  GTECH_NOT I_705 ( .A(a2stg_frac2[34]), .Z(N3945) );
  GTECH_AND2 C6759 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3940), .Z(N3947) );
  GTECH_AND2 C6761 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[34]), .Z(N3949)
         );
  GTECH_OR2 C6762 ( .A(N3953), .B(N3954), .Z(a2stg_fracadd_in2[33]) );
  GTECH_OR2 C6763 ( .A(N3951), .B(N3952), .Z(N3953) );
  GTECH_AND2 C6764 ( .A(a2stg_fracadd_frac2_inv), .B(N3950), .Z(N3951) );
  GTECH_NOT I_706 ( .A(a2stg_frac2[33]), .Z(N3950) );
  GTECH_AND2 C6766 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3945), .Z(N3952) );
  GTECH_AND2 C6768 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[33]), .Z(N3954)
         );
  GTECH_OR2 C6769 ( .A(N3958), .B(N3959), .Z(a2stg_fracadd_in2[32]) );
  GTECH_OR2 C6770 ( .A(N3956), .B(N3957), .Z(N3958) );
  GTECH_AND2 C6771 ( .A(a2stg_fracadd_frac2_inv), .B(N3955), .Z(N3956) );
  GTECH_NOT I_707 ( .A(a2stg_frac2[32]), .Z(N3955) );
  GTECH_AND2 C6773 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3950), .Z(N3957) );
  GTECH_AND2 C6775 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[32]), .Z(N3959)
         );
  GTECH_OR2 C6776 ( .A(N3963), .B(N3964), .Z(a2stg_fracadd_in2[31]) );
  GTECH_OR2 C6777 ( .A(N3961), .B(N3962), .Z(N3963) );
  GTECH_AND2 C6778 ( .A(a2stg_fracadd_frac2_inv), .B(N3960), .Z(N3961) );
  GTECH_NOT I_708 ( .A(a2stg_frac2[31]), .Z(N3960) );
  GTECH_AND2 C6780 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3955), .Z(N3962) );
  GTECH_AND2 C6782 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[31]), .Z(N3964)
         );
  GTECH_OR2 C6783 ( .A(N3968), .B(N3969), .Z(a2stg_fracadd_in2[30]) );
  GTECH_OR2 C6784 ( .A(N3966), .B(N3967), .Z(N3968) );
  GTECH_AND2 C6785 ( .A(a2stg_fracadd_frac2_inv), .B(N3965), .Z(N3966) );
  GTECH_NOT I_709 ( .A(a2stg_frac2[30]), .Z(N3965) );
  GTECH_AND2 C6787 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3960), .Z(N3967) );
  GTECH_AND2 C6789 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[30]), .Z(N3969)
         );
  GTECH_OR2 C6790 ( .A(N3973), .B(N3974), .Z(a2stg_fracadd_in2[29]) );
  GTECH_OR2 C6791 ( .A(N3971), .B(N3972), .Z(N3973) );
  GTECH_AND2 C6792 ( .A(a2stg_fracadd_frac2_inv), .B(N3970), .Z(N3971) );
  GTECH_NOT I_710 ( .A(a2stg_frac2[29]), .Z(N3970) );
  GTECH_AND2 C6794 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3965), .Z(N3972) );
  GTECH_AND2 C6796 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[29]), .Z(N3974)
         );
  GTECH_OR2 C6797 ( .A(N3978), .B(N3979), .Z(a2stg_fracadd_in2[28]) );
  GTECH_OR2 C6798 ( .A(N3976), .B(N3977), .Z(N3978) );
  GTECH_AND2 C6799 ( .A(a2stg_fracadd_frac2_inv), .B(N3975), .Z(N3976) );
  GTECH_NOT I_711 ( .A(a2stg_frac2[28]), .Z(N3975) );
  GTECH_AND2 C6801 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3970), .Z(N3977) );
  GTECH_AND2 C6803 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[28]), .Z(N3979)
         );
  GTECH_OR2 C6804 ( .A(N3983), .B(N3984), .Z(a2stg_fracadd_in2[27]) );
  GTECH_OR2 C6805 ( .A(N3981), .B(N3982), .Z(N3983) );
  GTECH_AND2 C6806 ( .A(a2stg_fracadd_frac2_inv), .B(N3980), .Z(N3981) );
  GTECH_NOT I_712 ( .A(a2stg_frac2[27]), .Z(N3980) );
  GTECH_AND2 C6808 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3975), .Z(N3982) );
  GTECH_AND2 C6810 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[27]), .Z(N3984)
         );
  GTECH_OR2 C6811 ( .A(N3988), .B(N3989), .Z(a2stg_fracadd_in2[26]) );
  GTECH_OR2 C6812 ( .A(N3986), .B(N3987), .Z(N3988) );
  GTECH_AND2 C6813 ( .A(a2stg_fracadd_frac2_inv), .B(N3985), .Z(N3986) );
  GTECH_NOT I_713 ( .A(a2stg_frac2[26]), .Z(N3985) );
  GTECH_AND2 C6815 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3980), .Z(N3987) );
  GTECH_AND2 C6817 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[26]), .Z(N3989)
         );
  GTECH_OR2 C6818 ( .A(N3993), .B(N3994), .Z(a2stg_fracadd_in2[25]) );
  GTECH_OR2 C6819 ( .A(N3991), .B(N3992), .Z(N3993) );
  GTECH_AND2 C6820 ( .A(a2stg_fracadd_frac2_inv), .B(N3990), .Z(N3991) );
  GTECH_NOT I_714 ( .A(a2stg_frac2[25]), .Z(N3990) );
  GTECH_AND2 C6822 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3985), .Z(N3992) );
  GTECH_AND2 C6824 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[25]), .Z(N3994)
         );
  GTECH_OR2 C6825 ( .A(N3998), .B(N3999), .Z(a2stg_fracadd_in2[24]) );
  GTECH_OR2 C6826 ( .A(N3996), .B(N3997), .Z(N3998) );
  GTECH_AND2 C6827 ( .A(a2stg_fracadd_frac2_inv), .B(N3995), .Z(N3996) );
  GTECH_NOT I_715 ( .A(a2stg_frac2[24]), .Z(N3995) );
  GTECH_AND2 C6829 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3990), .Z(N3997) );
  GTECH_AND2 C6831 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[24]), .Z(N3999)
         );
  GTECH_OR2 C6832 ( .A(N4003), .B(N4004), .Z(a2stg_fracadd_in2[23]) );
  GTECH_OR2 C6833 ( .A(N4001), .B(N4002), .Z(N4003) );
  GTECH_AND2 C6834 ( .A(a2stg_fracadd_frac2_inv), .B(N4000), .Z(N4001) );
  GTECH_NOT I_716 ( .A(a2stg_frac2[23]), .Z(N4000) );
  GTECH_AND2 C6836 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N3995), .Z(N4002) );
  GTECH_AND2 C6838 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[23]), .Z(N4004)
         );
  GTECH_OR2 C6839 ( .A(N4008), .B(N4009), .Z(a2stg_fracadd_in2[22]) );
  GTECH_OR2 C6840 ( .A(N4006), .B(N4007), .Z(N4008) );
  GTECH_AND2 C6841 ( .A(a2stg_fracadd_frac2_inv), .B(N4005), .Z(N4006) );
  GTECH_NOT I_717 ( .A(a2stg_frac2[22]), .Z(N4005) );
  GTECH_AND2 C6843 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4000), .Z(N4007) );
  GTECH_AND2 C6845 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[22]), .Z(N4009)
         );
  GTECH_OR2 C6846 ( .A(N4013), .B(N4014), .Z(a2stg_fracadd_in2[21]) );
  GTECH_OR2 C6847 ( .A(N4011), .B(N4012), .Z(N4013) );
  GTECH_AND2 C6848 ( .A(a2stg_fracadd_frac2_inv), .B(N4010), .Z(N4011) );
  GTECH_NOT I_718 ( .A(a2stg_frac2[21]), .Z(N4010) );
  GTECH_AND2 C6850 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4005), .Z(N4012) );
  GTECH_AND2 C6852 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[21]), .Z(N4014)
         );
  GTECH_OR2 C6853 ( .A(N4018), .B(N4019), .Z(a2stg_fracadd_in2[20]) );
  GTECH_OR2 C6854 ( .A(N4016), .B(N4017), .Z(N4018) );
  GTECH_AND2 C6855 ( .A(a2stg_fracadd_frac2_inv), .B(N4015), .Z(N4016) );
  GTECH_NOT I_719 ( .A(a2stg_frac2[20]), .Z(N4015) );
  GTECH_AND2 C6857 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4010), .Z(N4017) );
  GTECH_AND2 C6859 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[20]), .Z(N4019)
         );
  GTECH_OR2 C6860 ( .A(N4023), .B(N4024), .Z(a2stg_fracadd_in2[19]) );
  GTECH_OR2 C6861 ( .A(N4021), .B(N4022), .Z(N4023) );
  GTECH_AND2 C6862 ( .A(a2stg_fracadd_frac2_inv), .B(N4020), .Z(N4021) );
  GTECH_NOT I_720 ( .A(a2stg_frac2[19]), .Z(N4020) );
  GTECH_AND2 C6864 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4015), .Z(N4022) );
  GTECH_AND2 C6866 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[19]), .Z(N4024)
         );
  GTECH_OR2 C6867 ( .A(N4028), .B(N4029), .Z(a2stg_fracadd_in2[18]) );
  GTECH_OR2 C6868 ( .A(N4026), .B(N4027), .Z(N4028) );
  GTECH_AND2 C6869 ( .A(a2stg_fracadd_frac2_inv), .B(N4025), .Z(N4026) );
  GTECH_NOT I_721 ( .A(a2stg_frac2[18]), .Z(N4025) );
  GTECH_AND2 C6871 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4020), .Z(N4027) );
  GTECH_AND2 C6873 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[18]), .Z(N4029)
         );
  GTECH_OR2 C6874 ( .A(N4033), .B(N4034), .Z(a2stg_fracadd_in2[17]) );
  GTECH_OR2 C6875 ( .A(N4031), .B(N4032), .Z(N4033) );
  GTECH_AND2 C6876 ( .A(a2stg_fracadd_frac2_inv), .B(N4030), .Z(N4031) );
  GTECH_NOT I_722 ( .A(a2stg_frac2[17]), .Z(N4030) );
  GTECH_AND2 C6878 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4025), .Z(N4032) );
  GTECH_AND2 C6880 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[17]), .Z(N4034)
         );
  GTECH_OR2 C6881 ( .A(N4038), .B(N4039), .Z(a2stg_fracadd_in2[16]) );
  GTECH_OR2 C6882 ( .A(N4036), .B(N4037), .Z(N4038) );
  GTECH_AND2 C6883 ( .A(a2stg_fracadd_frac2_inv), .B(N4035), .Z(N4036) );
  GTECH_NOT I_723 ( .A(a2stg_frac2[16]), .Z(N4035) );
  GTECH_AND2 C6885 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4030), .Z(N4037) );
  GTECH_AND2 C6887 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[16]), .Z(N4039)
         );
  GTECH_OR2 C6888 ( .A(N4043), .B(N4044), .Z(a2stg_fracadd_in2[15]) );
  GTECH_OR2 C6889 ( .A(N4041), .B(N4042), .Z(N4043) );
  GTECH_AND2 C6890 ( .A(a2stg_fracadd_frac2_inv), .B(N4040), .Z(N4041) );
  GTECH_NOT I_724 ( .A(a2stg_frac2[15]), .Z(N4040) );
  GTECH_AND2 C6892 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4035), .Z(N4042) );
  GTECH_AND2 C6894 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[15]), .Z(N4044)
         );
  GTECH_OR2 C6895 ( .A(N4048), .B(N4049), .Z(a2stg_fracadd_in2[14]) );
  GTECH_OR2 C6896 ( .A(N4046), .B(N4047), .Z(N4048) );
  GTECH_AND2 C6897 ( .A(a2stg_fracadd_frac2_inv), .B(N4045), .Z(N4046) );
  GTECH_NOT I_725 ( .A(a2stg_frac2[14]), .Z(N4045) );
  GTECH_AND2 C6899 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4040), .Z(N4047) );
  GTECH_AND2 C6901 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[14]), .Z(N4049)
         );
  GTECH_OR2 C6902 ( .A(N4053), .B(N4054), .Z(a2stg_fracadd_in2[13]) );
  GTECH_OR2 C6903 ( .A(N4051), .B(N4052), .Z(N4053) );
  GTECH_AND2 C6904 ( .A(a2stg_fracadd_frac2_inv), .B(N4050), .Z(N4051) );
  GTECH_NOT I_726 ( .A(a2stg_frac2[13]), .Z(N4050) );
  GTECH_AND2 C6906 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4045), .Z(N4052) );
  GTECH_AND2 C6908 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[13]), .Z(N4054)
         );
  GTECH_OR2 C6909 ( .A(N4058), .B(N4059), .Z(a2stg_fracadd_in2[12]) );
  GTECH_OR2 C6910 ( .A(N4056), .B(N4057), .Z(N4058) );
  GTECH_AND2 C6911 ( .A(a2stg_fracadd_frac2_inv), .B(N4055), .Z(N4056) );
  GTECH_NOT I_727 ( .A(a2stg_frac2[12]), .Z(N4055) );
  GTECH_AND2 C6913 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4050), .Z(N4057) );
  GTECH_AND2 C6915 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[12]), .Z(N4059)
         );
  GTECH_OR2 C6916 ( .A(N4063), .B(N4064), .Z(a2stg_fracadd_in2[11]) );
  GTECH_OR2 C6917 ( .A(N4061), .B(N4062), .Z(N4063) );
  GTECH_AND2 C6918 ( .A(a2stg_fracadd_frac2_inv), .B(N4060), .Z(N4061) );
  GTECH_NOT I_728 ( .A(a2stg_frac2[11]), .Z(N4060) );
  GTECH_AND2 C6920 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4055), .Z(N4062) );
  GTECH_AND2 C6922 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[11]), .Z(N4064)
         );
  GTECH_OR2 C6923 ( .A(N4068), .B(N4069), .Z(a2stg_fracadd_in2[10]) );
  GTECH_OR2 C6924 ( .A(N4066), .B(N4067), .Z(N4068) );
  GTECH_AND2 C6925 ( .A(a2stg_fracadd_frac2_inv), .B(N4065), .Z(N4066) );
  GTECH_NOT I_729 ( .A(a2stg_frac2[10]), .Z(N4065) );
  GTECH_AND2 C6927 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4060), .Z(N4067) );
  GTECH_AND2 C6929 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[10]), .Z(N4069)
         );
  GTECH_OR2 C6930 ( .A(N4073), .B(N4074), .Z(a2stg_fracadd_in2[9]) );
  GTECH_OR2 C6931 ( .A(N4071), .B(N4072), .Z(N4073) );
  GTECH_AND2 C6932 ( .A(a2stg_fracadd_frac2_inv), .B(N4070), .Z(N4071) );
  GTECH_NOT I_730 ( .A(a2stg_frac2[9]), .Z(N4070) );
  GTECH_AND2 C6934 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4065), .Z(N4072) );
  GTECH_AND2 C6936 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[9]), .Z(N4074) );
  GTECH_OR2 C6937 ( .A(N4078), .B(N4079), .Z(a2stg_fracadd_in2[8]) );
  GTECH_OR2 C6938 ( .A(N4076), .B(N4077), .Z(N4078) );
  GTECH_AND2 C6939 ( .A(a2stg_fracadd_frac2_inv), .B(N4075), .Z(N4076) );
  GTECH_NOT I_731 ( .A(a2stg_frac2[8]), .Z(N4075) );
  GTECH_AND2 C6941 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4070), .Z(N4077) );
  GTECH_AND2 C6943 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[8]), .Z(N4079) );
  GTECH_OR2 C6944 ( .A(N4083), .B(N4084), .Z(a2stg_fracadd_in2[7]) );
  GTECH_OR2 C6945 ( .A(N4081), .B(N4082), .Z(N4083) );
  GTECH_AND2 C6946 ( .A(a2stg_fracadd_frac2_inv), .B(N4080), .Z(N4081) );
  GTECH_NOT I_732 ( .A(a2stg_frac2[7]), .Z(N4080) );
  GTECH_AND2 C6948 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4075), .Z(N4082) );
  GTECH_AND2 C6950 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[7]), .Z(N4084) );
  GTECH_OR2 C6951 ( .A(N4088), .B(N4089), .Z(a2stg_fracadd_in2[6]) );
  GTECH_OR2 C6952 ( .A(N4086), .B(N4087), .Z(N4088) );
  GTECH_AND2 C6953 ( .A(a2stg_fracadd_frac2_inv), .B(N4085), .Z(N4086) );
  GTECH_NOT I_733 ( .A(a2stg_frac2[6]), .Z(N4085) );
  GTECH_AND2 C6955 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4080), .Z(N4087) );
  GTECH_AND2 C6957 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[6]), .Z(N4089) );
  GTECH_OR2 C6958 ( .A(N4093), .B(N4094), .Z(a2stg_fracadd_in2[5]) );
  GTECH_OR2 C6959 ( .A(N4091), .B(N4092), .Z(N4093) );
  GTECH_AND2 C6960 ( .A(a2stg_fracadd_frac2_inv), .B(N4090), .Z(N4091) );
  GTECH_NOT I_734 ( .A(a2stg_frac2[5]), .Z(N4090) );
  GTECH_AND2 C6962 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4085), .Z(N4092) );
  GTECH_AND2 C6964 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[5]), .Z(N4094) );
  GTECH_OR2 C6965 ( .A(N4098), .B(N4099), .Z(a2stg_fracadd_in2[4]) );
  GTECH_OR2 C6966 ( .A(N4096), .B(N4097), .Z(N4098) );
  GTECH_AND2 C6967 ( .A(a2stg_fracadd_frac2_inv), .B(N4095), .Z(N4096) );
  GTECH_NOT I_735 ( .A(a2stg_frac2[4]), .Z(N4095) );
  GTECH_AND2 C6969 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4090), .Z(N4097) );
  GTECH_AND2 C6971 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[4]), .Z(N4099) );
  GTECH_OR2 C6972 ( .A(N4103), .B(N4104), .Z(a2stg_fracadd_in2[3]) );
  GTECH_OR2 C6973 ( .A(N4101), .B(N4102), .Z(N4103) );
  GTECH_AND2 C6974 ( .A(a2stg_fracadd_frac2_inv), .B(N4100), .Z(N4101) );
  GTECH_NOT I_736 ( .A(a2stg_frac2[3]), .Z(N4100) );
  GTECH_AND2 C6976 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4095), .Z(N4102) );
  GTECH_AND2 C6978 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[3]), .Z(N4104) );
  GTECH_OR2 C6979 ( .A(N4108), .B(N4109), .Z(a2stg_fracadd_in2[2]) );
  GTECH_OR2 C6980 ( .A(N4106), .B(N4107), .Z(N4108) );
  GTECH_AND2 C6981 ( .A(a2stg_fracadd_frac2_inv), .B(N4105), .Z(N4106) );
  GTECH_NOT I_737 ( .A(a2stg_frac2[2]), .Z(N4105) );
  GTECH_AND2 C6983 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4100), .Z(N4107) );
  GTECH_AND2 C6985 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[2]), .Z(N4109) );
  GTECH_OR2 C6986 ( .A(N4113), .B(N4114), .Z(a2stg_fracadd_in2[1]) );
  GTECH_OR2 C6987 ( .A(N4111), .B(N4112), .Z(N4113) );
  GTECH_AND2 C6988 ( .A(a2stg_fracadd_frac2_inv), .B(N4110), .Z(N4111) );
  GTECH_NOT I_738 ( .A(a2stg_frac2[1]), .Z(N4110) );
  GTECH_AND2 C6990 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4105), .Z(N4112) );
  GTECH_AND2 C6992 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[1]), .Z(N4114) );
  GTECH_OR2 C6993 ( .A(N4118), .B(N4119), .Z(a2stg_fracadd_in2[0]) );
  GTECH_OR2 C6994 ( .A(N4116), .B(N4117), .Z(N4118) );
  GTECH_AND2 C6995 ( .A(a2stg_fracadd_frac2_inv), .B(N4115), .Z(N4116) );
  GTECH_NOT I_739 ( .A(a2stg_frac2[0]), .Z(N4115) );
  GTECH_AND2 C6997 ( .A(a2stg_fracadd_frac2_inv_shr1), .B(N4110), .Z(N4117) );
  GTECH_AND2 C6999 ( .A(a2stg_fracadd_frac2), .B(a2stg_frac2[0]), .Z(N4119) );
  GTECH_AND2 C7000 ( .A(a2stg_expdec_tmp[53]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[53]) );
  GTECH_AND2 C7001 ( .A(a2stg_expdec_tmp[52]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[52]) );
  GTECH_AND2 C7002 ( .A(a2stg_expdec_tmp[51]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[51]) );
  GTECH_AND2 C7003 ( .A(a2stg_expdec_tmp[50]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[50]) );
  GTECH_AND2 C7004 ( .A(a2stg_expdec_tmp[49]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[49]) );
  GTECH_AND2 C7005 ( .A(a2stg_expdec_tmp[48]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[48]) );
  GTECH_AND2 C7006 ( .A(a2stg_expdec_tmp[47]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[47]) );
  GTECH_AND2 C7007 ( .A(a2stg_expdec_tmp[46]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[46]) );
  GTECH_AND2 C7008 ( .A(a2stg_expdec_tmp[45]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[45]) );
  GTECH_AND2 C7009 ( .A(a2stg_expdec_tmp[44]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[44]) );
  GTECH_AND2 C7010 ( .A(a2stg_expdec_tmp[43]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[43]) );
  GTECH_AND2 C7011 ( .A(a2stg_expdec_tmp[42]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[42]) );
  GTECH_AND2 C7012 ( .A(a2stg_expdec_tmp[41]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[41]) );
  GTECH_AND2 C7013 ( .A(a2stg_expdec_tmp[40]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[40]) );
  GTECH_AND2 C7014 ( .A(a2stg_expdec_tmp[39]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[39]) );
  GTECH_AND2 C7015 ( .A(a2stg_expdec_tmp[38]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[38]) );
  GTECH_AND2 C7016 ( .A(a2stg_expdec_tmp[37]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[37]) );
  GTECH_AND2 C7017 ( .A(a2stg_expdec_tmp[36]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[36]) );
  GTECH_AND2 C7018 ( .A(a2stg_expdec_tmp[35]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[35]) );
  GTECH_AND2 C7019 ( .A(a2stg_expdec_tmp[34]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[34]) );
  GTECH_AND2 C7020 ( .A(a2stg_expdec_tmp[33]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[33]) );
  GTECH_AND2 C7021 ( .A(a2stg_expdec_tmp[32]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[32]) );
  GTECH_AND2 C7022 ( .A(a2stg_expdec_tmp[31]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[31]) );
  GTECH_AND2 C7023 ( .A(a2stg_expdec_tmp[30]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[30]) );
  GTECH_AND2 C7024 ( .A(a2stg_expdec_tmp[29]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[29]) );
  GTECH_AND2 C7025 ( .A(a2stg_expdec_tmp[28]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[28]) );
  GTECH_AND2 C7026 ( .A(a2stg_expdec_tmp[27]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[27]) );
  GTECH_AND2 C7027 ( .A(a2stg_expdec_tmp[26]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[26]) );
  GTECH_AND2 C7028 ( .A(a2stg_expdec_tmp[25]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[25]) );
  GTECH_AND2 C7029 ( .A(a2stg_expdec_tmp[24]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[24]) );
  GTECH_AND2 C7030 ( .A(a2stg_expdec_tmp[23]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[23]) );
  GTECH_AND2 C7031 ( .A(a2stg_expdec_tmp[22]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[22]) );
  GTECH_AND2 C7032 ( .A(a2stg_expdec_tmp[21]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[21]) );
  GTECH_AND2 C7033 ( .A(a2stg_expdec_tmp[20]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[20]) );
  GTECH_AND2 C7034 ( .A(a2stg_expdec_tmp[19]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[19]) );
  GTECH_AND2 C7035 ( .A(a2stg_expdec_tmp[18]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[18]) );
  GTECH_AND2 C7036 ( .A(a2stg_expdec_tmp[17]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[17]) );
  GTECH_AND2 C7037 ( .A(a2stg_expdec_tmp[16]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[16]) );
  GTECH_AND2 C7038 ( .A(a2stg_expdec_tmp[15]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[15]) );
  GTECH_AND2 C7039 ( .A(a2stg_expdec_tmp[14]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[14]) );
  GTECH_AND2 C7040 ( .A(a2stg_expdec_tmp[13]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[13]) );
  GTECH_AND2 C7041 ( .A(a2stg_expdec_tmp[12]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[12]) );
  GTECH_AND2 C7042 ( .A(a2stg_expdec_tmp[11]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[11]) );
  GTECH_AND2 C7043 ( .A(a2stg_expdec_tmp[10]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[10]) );
  GTECH_AND2 C7044 ( .A(a2stg_expdec_tmp[9]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[9]) );
  GTECH_AND2 C7045 ( .A(a2stg_expdec_tmp[8]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[8]) );
  GTECH_AND2 C7046 ( .A(a2stg_expdec_tmp[7]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[7]) );
  GTECH_AND2 C7047 ( .A(a2stg_expdec_tmp[6]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[6]) );
  GTECH_AND2 C7048 ( .A(a2stg_expdec_tmp[5]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[5]) );
  GTECH_AND2 C7049 ( .A(a2stg_expdec_tmp[4]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[4]) );
  GTECH_AND2 C7050 ( .A(a2stg_expdec_tmp[3]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[3]) );
  GTECH_AND2 C7051 ( .A(a2stg_expdec_tmp[2]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[2]) );
  GTECH_AND2 C7052 ( .A(a2stg_expdec_tmp[1]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[1]) );
  GTECH_AND2 C7053 ( .A(a2stg_expdec_tmp[0]), .B(a2stg_expdec_neq_0), .Z(
        a2stg_expdec[0]) );
  GTECH_OR2 C7054 ( .A(N4120), .B(N4132), .Z(a3stg_ld0_dnrm_10) );
  GTECH_AND2 C7055 ( .A(a3stg_faddsubopa[0]), .B(a3stg_ld0_frac[10]), .Z(N4120) );
  GTECH_AND2 C7056 ( .A(N4121), .B(N4131), .Z(N4132) );
  GTECH_NOT I_740 ( .A(a3stg_faddsubopa[0]), .Z(N4121) );
  GTECH_OR2 C7058 ( .A(N4130), .B(a3stg_ld0_frac[0]), .Z(N4131) );
  GTECH_OR2 C7059 ( .A(N4129), .B(a3stg_ld0_frac[1]), .Z(N4130) );
  GTECH_OR2 C7060 ( .A(N4128), .B(a3stg_ld0_frac[2]), .Z(N4129) );
  GTECH_OR2 C7061 ( .A(N4127), .B(a3stg_ld0_frac[3]), .Z(N4128) );
  GTECH_OR2 C7062 ( .A(N4126), .B(a3stg_ld0_frac[4]), .Z(N4127) );
  GTECH_OR2 C7063 ( .A(N4125), .B(a3stg_ld0_frac[5]), .Z(N4126) );
  GTECH_OR2 C7064 ( .A(N4124), .B(a3stg_ld0_frac[6]), .Z(N4125) );
  GTECH_OR2 C7065 ( .A(N4123), .B(a3stg_ld0_frac[7]), .Z(N4124) );
  GTECH_OR2 C7066 ( .A(N4122), .B(a3stg_ld0_frac[8]), .Z(N4123) );
  GTECH_OR2 C7067 ( .A(a3stg_ld0_frac[10]), .B(a3stg_ld0_frac[9]), .Z(N4122)
         );
  GTECH_OR2 C7068 ( .A(N4133), .B(a3stg_fracadd[63]), .Z(a4stg_round_in) );
  GTECH_OR2 C7069 ( .A(a3stg_fracadd[61]), .B(a3stg_fracadd[62]), .Z(N4133) );
  GTECH_NOT I_741 ( .A(a3stg_fracadd[63]), .Z(a3stg_inc_exp_inv) );
  GTECH_NOT I_742 ( .A(a3stg_fracadd[63]), .Z(N130) );
  GTECH_NOT I_743 ( .A(N4136), .Z(a3stg_same_exp_inv) );
  GTECH_OR2 C7073 ( .A(N4134), .B(N4135), .Z(N4136) );
  GTECH_AND2 C7074 ( .A(N130), .B(a3stg_fracadd[62]), .Z(N4134) );
  GTECH_AND2 C7075 ( .A(N130), .B(a3stg_exp10_0_eq0), .Z(N4135) );
  GTECH_NOT I_744 ( .A(N4141), .Z(a3stg_dec_exp_inv) );
  GTECH_AND2 C7077 ( .A(N4139), .B(N4140), .Z(N4141) );
  GTECH_AND2 C7078 ( .A(N4138), .B(a3stg_fracadd[61]), .Z(N4139) );
  GTECH_AND2 C7079 ( .A(N130), .B(N4137), .Z(N4138) );
  GTECH_NOT I_745 ( .A(a3stg_fracadd[62]), .Z(N4137) );
  GTECH_NOT I_746 ( .A(a3stg_exp10_0_eq0), .Z(N4140) );
  GTECH_NOT I_747 ( .A(a3stg_fracadd[63]), .Z(a3stg_inc_exp_inva) );
  GTECH_NOT I_748 ( .A(N4148), .Z(a3stg_fsame_exp_inv) );
  GTECH_OR2 C7086 ( .A(N4145), .B(N4147), .Z(N4148) );
  GTECH_AND2 C7087 ( .A(N4144), .B(a3stg_exp_0), .Z(N4145) );
  GTECH_AND2 C7088 ( .A(N4143), .B(a3stg_exp10_1_eq0), .Z(N4144) );
  GTECH_AND2 C7089 ( .A(N4142), .B(a3stg_fracadd[61]), .Z(N4143) );
  GTECH_AND2 C7090 ( .A(N130), .B(N4137), .Z(N4142) );
  GTECH_AND2 C7092 ( .A(N4146), .B(N4140), .Z(N4147) );
  GTECH_AND2 C7093 ( .A(N130), .B(a3stg_fracadd[62]), .Z(N4146) );
  GTECH_NOT I_749 ( .A(N4152), .Z(a3stg_fdec_exp_inv) );
  GTECH_AND2 C7096 ( .A(N4150), .B(N4151), .Z(N4152) );
  GTECH_AND2 C7097 ( .A(N4149), .B(a3stg_fracadd[61]), .Z(N4150) );
  GTECH_AND2 C7098 ( .A(N130), .B(N4137), .Z(N4149) );
  GTECH_NOT I_750 ( .A(a3stg_exp10_1_eq0), .Z(N4151) );
  GTECH_AND2 C7102 ( .A(N4155), .B(a3stg_fracadd[61]), .Z(
        a4stg_rnd_frac_pre1_in[63]) );
  GTECH_AND2 C7103 ( .A(N4153), .B(N4154), .Z(N4155) );
  GTECH_AND2 C7104 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4153) );
  GTECH_NOT I_751 ( .A(a3stg_fdec_exp_inv), .Z(N4154) );
  GTECH_AND2 C7106 ( .A(N4157), .B(a3stg_fracadd[60]), .Z(
        a4stg_rnd_frac_pre1_in[62]) );
  GTECH_AND2 C7107 ( .A(N4156), .B(N4154), .Z(N4157) );
  GTECH_AND2 C7108 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4156) );
  GTECH_AND2 C7110 ( .A(N4159), .B(a3stg_fracadd[59]), .Z(
        a4stg_rnd_frac_pre1_in[61]) );
  GTECH_AND2 C7111 ( .A(N4158), .B(N4154), .Z(N4159) );
  GTECH_AND2 C7112 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4158) );
  GTECH_AND2 C7114 ( .A(N4161), .B(a3stg_fracadd[58]), .Z(
        a4stg_rnd_frac_pre1_in[60]) );
  GTECH_AND2 C7115 ( .A(N4160), .B(N4154), .Z(N4161) );
  GTECH_AND2 C7116 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4160) );
  GTECH_AND2 C7118 ( .A(N4163), .B(a3stg_fracadd[57]), .Z(
        a4stg_rnd_frac_pre1_in[59]) );
  GTECH_AND2 C7119 ( .A(N4162), .B(N4154), .Z(N4163) );
  GTECH_AND2 C7120 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4162) );
  GTECH_AND2 C7122 ( .A(N4165), .B(a3stg_fracadd[56]), .Z(
        a4stg_rnd_frac_pre1_in[58]) );
  GTECH_AND2 C7123 ( .A(N4164), .B(N4154), .Z(N4165) );
  GTECH_AND2 C7124 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4164) );
  GTECH_AND2 C7126 ( .A(N4167), .B(a3stg_fracadd[55]), .Z(
        a4stg_rnd_frac_pre1_in[57]) );
  GTECH_AND2 C7127 ( .A(N4166), .B(N4154), .Z(N4167) );
  GTECH_AND2 C7128 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4166) );
  GTECH_AND2 C7130 ( .A(N4169), .B(a3stg_fracadd[54]), .Z(
        a4stg_rnd_frac_pre1_in[56]) );
  GTECH_AND2 C7131 ( .A(N4168), .B(N4154), .Z(N4169) );
  GTECH_AND2 C7132 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4168) );
  GTECH_AND2 C7134 ( .A(N4171), .B(a3stg_fracadd[53]), .Z(
        a4stg_rnd_frac_pre1_in[55]) );
  GTECH_AND2 C7135 ( .A(N4170), .B(N4154), .Z(N4171) );
  GTECH_AND2 C7136 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4170) );
  GTECH_AND2 C7138 ( .A(N4173), .B(a3stg_fracadd[52]), .Z(
        a4stg_rnd_frac_pre1_in[54]) );
  GTECH_AND2 C7139 ( .A(N4172), .B(N4154), .Z(N4173) );
  GTECH_AND2 C7140 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4172) );
  GTECH_AND2 C7142 ( .A(N4175), .B(a3stg_fracadd[51]), .Z(
        a4stg_rnd_frac_pre1_in[53]) );
  GTECH_AND2 C7143 ( .A(N4174), .B(N4154), .Z(N4175) );
  GTECH_AND2 C7144 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4174) );
  GTECH_AND2 C7146 ( .A(N4177), .B(a3stg_fracadd[50]), .Z(
        a4stg_rnd_frac_pre1_in[52]) );
  GTECH_AND2 C7147 ( .A(N4176), .B(N4154), .Z(N4177) );
  GTECH_AND2 C7148 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4176) );
  GTECH_AND2 C7150 ( .A(N4179), .B(a3stg_fracadd[49]), .Z(
        a4stg_rnd_frac_pre1_in[51]) );
  GTECH_AND2 C7151 ( .A(N4178), .B(N4154), .Z(N4179) );
  GTECH_AND2 C7152 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4178) );
  GTECH_AND2 C7154 ( .A(N4181), .B(a3stg_fracadd[48]), .Z(
        a4stg_rnd_frac_pre1_in[50]) );
  GTECH_AND2 C7155 ( .A(N4180), .B(N4154), .Z(N4181) );
  GTECH_AND2 C7156 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4180) );
  GTECH_AND2 C7158 ( .A(N4183), .B(a3stg_fracadd[47]), .Z(
        a4stg_rnd_frac_pre1_in[49]) );
  GTECH_AND2 C7159 ( .A(N4182), .B(N4154), .Z(N4183) );
  GTECH_AND2 C7160 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4182) );
  GTECH_AND2 C7162 ( .A(N4185), .B(a3stg_fracadd[46]), .Z(
        a4stg_rnd_frac_pre1_in[48]) );
  GTECH_AND2 C7163 ( .A(N4184), .B(N4154), .Z(N4185) );
  GTECH_AND2 C7164 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4184) );
  GTECH_AND2 C7166 ( .A(N4187), .B(a3stg_fracadd[45]), .Z(
        a4stg_rnd_frac_pre1_in[47]) );
  GTECH_AND2 C7167 ( .A(N4186), .B(N4154), .Z(N4187) );
  GTECH_AND2 C7168 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4186) );
  GTECH_AND2 C7170 ( .A(N4189), .B(a3stg_fracadd[44]), .Z(
        a4stg_rnd_frac_pre1_in[46]) );
  GTECH_AND2 C7171 ( .A(N4188), .B(N4154), .Z(N4189) );
  GTECH_AND2 C7172 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4188) );
  GTECH_AND2 C7174 ( .A(N4191), .B(a3stg_fracadd[43]), .Z(
        a4stg_rnd_frac_pre1_in[45]) );
  GTECH_AND2 C7175 ( .A(N4190), .B(N4154), .Z(N4191) );
  GTECH_AND2 C7176 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4190) );
  GTECH_AND2 C7178 ( .A(N4193), .B(a3stg_fracadd[42]), .Z(
        a4stg_rnd_frac_pre1_in[44]) );
  GTECH_AND2 C7179 ( .A(N4192), .B(N4154), .Z(N4193) );
  GTECH_AND2 C7180 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4192) );
  GTECH_AND2 C7182 ( .A(N4195), .B(a3stg_fracadd[41]), .Z(
        a4stg_rnd_frac_pre1_in[43]) );
  GTECH_AND2 C7183 ( .A(N4194), .B(N4154), .Z(N4195) );
  GTECH_AND2 C7184 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4194) );
  GTECH_AND2 C7186 ( .A(N4197), .B(a3stg_fracadd[40]), .Z(
        a4stg_rnd_frac_pre1_in[42]) );
  GTECH_AND2 C7187 ( .A(N4196), .B(N4154), .Z(N4197) );
  GTECH_AND2 C7188 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4196) );
  GTECH_AND2 C7190 ( .A(N4199), .B(a3stg_fracadd[39]), .Z(
        a4stg_rnd_frac_pre1_in[41]) );
  GTECH_AND2 C7191 ( .A(N4198), .B(N4154), .Z(N4199) );
  GTECH_AND2 C7192 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4198) );
  GTECH_AND2 C7194 ( .A(N4201), .B(a3stg_fracadd[38]), .Z(
        a4stg_rnd_frac_pre1_in[40]) );
  GTECH_AND2 C7195 ( .A(N4200), .B(N4154), .Z(N4201) );
  GTECH_AND2 C7196 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4200) );
  GTECH_AND2 C7198 ( .A(N4203), .B(a3stg_fracadd[37]), .Z(
        a4stg_rnd_frac_pre1_in[39]) );
  GTECH_AND2 C7199 ( .A(N4202), .B(N4154), .Z(N4203) );
  GTECH_AND2 C7200 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4202) );
  GTECH_AND2 C7202 ( .A(N4205), .B(a3stg_fracadd[36]), .Z(
        a4stg_rnd_frac_pre1_in[38]) );
  GTECH_AND2 C7203 ( .A(N4204), .B(N4154), .Z(N4205) );
  GTECH_AND2 C7204 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4204) );
  GTECH_AND2 C7206 ( .A(N4207), .B(a3stg_fracadd[35]), .Z(
        a4stg_rnd_frac_pre1_in[37]) );
  GTECH_AND2 C7207 ( .A(N4206), .B(N4154), .Z(N4207) );
  GTECH_AND2 C7208 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4206) );
  GTECH_AND2 C7210 ( .A(N4209), .B(a3stg_fracadd[34]), .Z(
        a4stg_rnd_frac_pre1_in[36]) );
  GTECH_AND2 C7211 ( .A(N4208), .B(N4154), .Z(N4209) );
  GTECH_AND2 C7212 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4208) );
  GTECH_AND2 C7214 ( .A(N4211), .B(a3stg_fracadd[33]), .Z(
        a4stg_rnd_frac_pre1_in[35]) );
  GTECH_AND2 C7215 ( .A(N4210), .B(N4154), .Z(N4211) );
  GTECH_AND2 C7216 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4210) );
  GTECH_AND2 C7218 ( .A(N4213), .B(a3stg_fracadd[32]), .Z(
        a4stg_rnd_frac_pre1_in[34]) );
  GTECH_AND2 C7219 ( .A(N4212), .B(N4154), .Z(N4213) );
  GTECH_AND2 C7220 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4212) );
  GTECH_AND2 C7222 ( .A(N4215), .B(a3stg_fracadd[31]), .Z(
        a4stg_rnd_frac_pre1_in[33]) );
  GTECH_AND2 C7223 ( .A(N4214), .B(N4154), .Z(N4215) );
  GTECH_AND2 C7224 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4214) );
  GTECH_AND2 C7226 ( .A(N4217), .B(a3stg_fracadd[30]), .Z(
        a4stg_rnd_frac_pre1_in[32]) );
  GTECH_AND2 C7227 ( .A(N4216), .B(N4154), .Z(N4217) );
  GTECH_AND2 C7228 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4216) );
  GTECH_AND2 C7230 ( .A(N4219), .B(a3stg_fracadd[29]), .Z(
        a4stg_rnd_frac_pre1_in[31]) );
  GTECH_AND2 C7231 ( .A(N4218), .B(N4154), .Z(N4219) );
  GTECH_AND2 C7232 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4218) );
  GTECH_AND2 C7234 ( .A(N4221), .B(a3stg_fracadd[28]), .Z(
        a4stg_rnd_frac_pre1_in[30]) );
  GTECH_AND2 C7235 ( .A(N4220), .B(N4154), .Z(N4221) );
  GTECH_AND2 C7236 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4220) );
  GTECH_AND2 C7238 ( .A(N4223), .B(a3stg_fracadd[27]), .Z(
        a4stg_rnd_frac_pre1_in[29]) );
  GTECH_AND2 C7239 ( .A(N4222), .B(N4154), .Z(N4223) );
  GTECH_AND2 C7240 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4222) );
  GTECH_AND2 C7242 ( .A(N4225), .B(a3stg_fracadd[26]), .Z(
        a4stg_rnd_frac_pre1_in[28]) );
  GTECH_AND2 C7243 ( .A(N4224), .B(N4154), .Z(N4225) );
  GTECH_AND2 C7244 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4224) );
  GTECH_AND2 C7246 ( .A(N4227), .B(a3stg_fracadd[25]), .Z(
        a4stg_rnd_frac_pre1_in[27]) );
  GTECH_AND2 C7247 ( .A(N4226), .B(N4154), .Z(N4227) );
  GTECH_AND2 C7248 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4226) );
  GTECH_AND2 C7250 ( .A(N4229), .B(a3stg_fracadd[24]), .Z(
        a4stg_rnd_frac_pre1_in[26]) );
  GTECH_AND2 C7251 ( .A(N4228), .B(N4154), .Z(N4229) );
  GTECH_AND2 C7252 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4228) );
  GTECH_AND2 C7254 ( .A(N4231), .B(a3stg_fracadd[23]), .Z(
        a4stg_rnd_frac_pre1_in[25]) );
  GTECH_AND2 C7255 ( .A(N4230), .B(N4154), .Z(N4231) );
  GTECH_AND2 C7256 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4230) );
  GTECH_AND2 C7258 ( .A(N4233), .B(a3stg_fracadd[22]), .Z(
        a4stg_rnd_frac_pre1_in[24]) );
  GTECH_AND2 C7259 ( .A(N4232), .B(N4154), .Z(N4233) );
  GTECH_AND2 C7260 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4232) );
  GTECH_AND2 C7262 ( .A(N4235), .B(a3stg_fracadd[21]), .Z(
        a4stg_rnd_frac_pre1_in[23]) );
  GTECH_AND2 C7263 ( .A(N4234), .B(N4154), .Z(N4235) );
  GTECH_AND2 C7264 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4234) );
  GTECH_AND2 C7266 ( .A(N4237), .B(a3stg_fracadd[20]), .Z(
        a4stg_rnd_frac_pre1_in[22]) );
  GTECH_AND2 C7267 ( .A(N4236), .B(N4154), .Z(N4237) );
  GTECH_AND2 C7268 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4236) );
  GTECH_AND2 C7270 ( .A(N4239), .B(a3stg_fracadd[19]), .Z(
        a4stg_rnd_frac_pre1_in[21]) );
  GTECH_AND2 C7271 ( .A(N4238), .B(N4154), .Z(N4239) );
  GTECH_AND2 C7272 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4238) );
  GTECH_AND2 C7274 ( .A(N4241), .B(a3stg_fracadd[18]), .Z(
        a4stg_rnd_frac_pre1_in[20]) );
  GTECH_AND2 C7275 ( .A(N4240), .B(N4154), .Z(N4241) );
  GTECH_AND2 C7276 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4240) );
  GTECH_AND2 C7278 ( .A(N4243), .B(a3stg_fracadd[17]), .Z(
        a4stg_rnd_frac_pre1_in[19]) );
  GTECH_AND2 C7279 ( .A(N4242), .B(N4154), .Z(N4243) );
  GTECH_AND2 C7280 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4242) );
  GTECH_AND2 C7282 ( .A(N4245), .B(a3stg_fracadd[16]), .Z(
        a4stg_rnd_frac_pre1_in[18]) );
  GTECH_AND2 C7283 ( .A(N4244), .B(N4154), .Z(N4245) );
  GTECH_AND2 C7284 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4244) );
  GTECH_AND2 C7286 ( .A(N4247), .B(a3stg_fracadd[15]), .Z(
        a4stg_rnd_frac_pre1_in[17]) );
  GTECH_AND2 C7287 ( .A(N4246), .B(N4154), .Z(N4247) );
  GTECH_AND2 C7288 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4246) );
  GTECH_AND2 C7290 ( .A(N4249), .B(a3stg_fracadd[14]), .Z(
        a4stg_rnd_frac_pre1_in[16]) );
  GTECH_AND2 C7291 ( .A(N4248), .B(N4154), .Z(N4249) );
  GTECH_AND2 C7292 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4248) );
  GTECH_AND2 C7294 ( .A(N4251), .B(a3stg_fracadd[13]), .Z(
        a4stg_rnd_frac_pre1_in[15]) );
  GTECH_AND2 C7295 ( .A(N4250), .B(N4154), .Z(N4251) );
  GTECH_AND2 C7296 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4250) );
  GTECH_AND2 C7298 ( .A(N4253), .B(a3stg_fracadd[12]), .Z(
        a4stg_rnd_frac_pre1_in[14]) );
  GTECH_AND2 C7299 ( .A(N4252), .B(N4154), .Z(N4253) );
  GTECH_AND2 C7300 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4252) );
  GTECH_AND2 C7302 ( .A(N4255), .B(a3stg_fracadd[11]), .Z(
        a4stg_rnd_frac_pre1_in[13]) );
  GTECH_AND2 C7303 ( .A(N4254), .B(N4154), .Z(N4255) );
  GTECH_AND2 C7304 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4254) );
  GTECH_AND2 C7306 ( .A(N4257), .B(a3stg_fracadd[10]), .Z(
        a4stg_rnd_frac_pre1_in[12]) );
  GTECH_AND2 C7307 ( .A(N4256), .B(N4154), .Z(N4257) );
  GTECH_AND2 C7308 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4256) );
  GTECH_AND2 C7310 ( .A(N4259), .B(a3stg_fracadd[9]), .Z(
        a4stg_rnd_frac_pre1_in[11]) );
  GTECH_AND2 C7311 ( .A(N4258), .B(N4154), .Z(N4259) );
  GTECH_AND2 C7312 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4258) );
  GTECH_AND2 C7314 ( .A(N4261), .B(a3stg_fracadd[8]), .Z(
        a4stg_rnd_frac_pre1_in[10]) );
  GTECH_AND2 C7315 ( .A(N4260), .B(N4154), .Z(N4261) );
  GTECH_AND2 C7316 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4260) );
  GTECH_AND2 C7318 ( .A(N4263), .B(a3stg_fracadd[7]), .Z(
        a4stg_rnd_frac_pre1_in[9]) );
  GTECH_AND2 C7319 ( .A(N4262), .B(N4154), .Z(N4263) );
  GTECH_AND2 C7320 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4262) );
  GTECH_AND2 C7322 ( .A(N4265), .B(a3stg_fracadd[6]), .Z(
        a4stg_rnd_frac_pre1_in[8]) );
  GTECH_AND2 C7323 ( .A(N4264), .B(N4154), .Z(N4265) );
  GTECH_AND2 C7324 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4264) );
  GTECH_AND2 C7326 ( .A(N4267), .B(a3stg_fracadd[5]), .Z(
        a4stg_rnd_frac_pre1_in[7]) );
  GTECH_AND2 C7327 ( .A(N4266), .B(N4154), .Z(N4267) );
  GTECH_AND2 C7328 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4266) );
  GTECH_AND2 C7330 ( .A(N4269), .B(a3stg_fracadd[4]), .Z(
        a4stg_rnd_frac_pre1_in[6]) );
  GTECH_AND2 C7331 ( .A(N4268), .B(N4154), .Z(N4269) );
  GTECH_AND2 C7332 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4268) );
  GTECH_AND2 C7334 ( .A(N4271), .B(a3stg_fracadd[3]), .Z(
        a4stg_rnd_frac_pre1_in[5]) );
  GTECH_AND2 C7335 ( .A(N4270), .B(N4154), .Z(N4271) );
  GTECH_AND2 C7336 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4270) );
  GTECH_AND2 C7338 ( .A(N4273), .B(a3stg_fracadd[2]), .Z(
        a4stg_rnd_frac_pre1_in[4]) );
  GTECH_AND2 C7339 ( .A(N4272), .B(N4154), .Z(N4273) );
  GTECH_AND2 C7340 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4272) );
  GTECH_AND2 C7342 ( .A(N4275), .B(a3stg_fracadd[1]), .Z(
        a4stg_rnd_frac_pre1_in[3]) );
  GTECH_AND2 C7343 ( .A(N4274), .B(N4154), .Z(N4275) );
  GTECH_AND2 C7344 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4274) );
  GTECH_AND2 C7346 ( .A(N4277), .B(a3stg_fracadd[0]), .Z(
        a4stg_rnd_frac_pre1_in[2]) );
  GTECH_AND2 C7347 ( .A(N4276), .B(N4154), .Z(N4277) );
  GTECH_AND2 C7348 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4276) );
  GTECH_AND2 C7350 ( .A(N4280), .B(a3stg_fracadd[62]), .Z(
        a4stg_rnd_frac_pre3_in[63]) );
  GTECH_AND2 C7351 ( .A(N4278), .B(N4279), .Z(N4280) );
  GTECH_AND2 C7352 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4278) );
  GTECH_NOT I_752 ( .A(a3stg_fsame_exp_inv), .Z(N4279) );
  GTECH_AND2 C7354 ( .A(N4282), .B(a3stg_fracadd[61]), .Z(
        a4stg_rnd_frac_pre3_in[62]) );
  GTECH_AND2 C7355 ( .A(N4281), .B(N4279), .Z(N4282) );
  GTECH_AND2 C7356 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4281) );
  GTECH_AND2 C7358 ( .A(N4284), .B(a3stg_fracadd[60]), .Z(
        a4stg_rnd_frac_pre3_in[61]) );
  GTECH_AND2 C7359 ( .A(N4283), .B(N4279), .Z(N4284) );
  GTECH_AND2 C7360 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4283) );
  GTECH_AND2 C7362 ( .A(N4286), .B(a3stg_fracadd[59]), .Z(
        a4stg_rnd_frac_pre3_in[60]) );
  GTECH_AND2 C7363 ( .A(N4285), .B(N4279), .Z(N4286) );
  GTECH_AND2 C7364 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4285) );
  GTECH_AND2 C7366 ( .A(N4288), .B(a3stg_fracadd[58]), .Z(
        a4stg_rnd_frac_pre3_in[59]) );
  GTECH_AND2 C7367 ( .A(N4287), .B(N4279), .Z(N4288) );
  GTECH_AND2 C7368 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4287) );
  GTECH_AND2 C7370 ( .A(N4290), .B(a3stg_fracadd[57]), .Z(
        a4stg_rnd_frac_pre3_in[58]) );
  GTECH_AND2 C7371 ( .A(N4289), .B(N4279), .Z(N4290) );
  GTECH_AND2 C7372 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4289) );
  GTECH_AND2 C7374 ( .A(N4292), .B(a3stg_fracadd[56]), .Z(
        a4stg_rnd_frac_pre3_in[57]) );
  GTECH_AND2 C7375 ( .A(N4291), .B(N4279), .Z(N4292) );
  GTECH_AND2 C7376 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4291) );
  GTECH_AND2 C7378 ( .A(N4294), .B(a3stg_fracadd[55]), .Z(
        a4stg_rnd_frac_pre3_in[56]) );
  GTECH_AND2 C7379 ( .A(N4293), .B(N4279), .Z(N4294) );
  GTECH_AND2 C7380 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4293) );
  GTECH_AND2 C7382 ( .A(N4296), .B(a3stg_fracadd[54]), .Z(
        a4stg_rnd_frac_pre3_in[55]) );
  GTECH_AND2 C7383 ( .A(N4295), .B(N4279), .Z(N4296) );
  GTECH_AND2 C7384 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4295) );
  GTECH_AND2 C7386 ( .A(N4298), .B(a3stg_fracadd[53]), .Z(
        a4stg_rnd_frac_pre3_in[54]) );
  GTECH_AND2 C7387 ( .A(N4297), .B(N4279), .Z(N4298) );
  GTECH_AND2 C7388 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4297) );
  GTECH_AND2 C7390 ( .A(N4300), .B(a3stg_fracadd[52]), .Z(
        a4stg_rnd_frac_pre3_in[53]) );
  GTECH_AND2 C7391 ( .A(N4299), .B(N4279), .Z(N4300) );
  GTECH_AND2 C7392 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4299) );
  GTECH_AND2 C7394 ( .A(N4302), .B(a3stg_fracadd[51]), .Z(
        a4stg_rnd_frac_pre3_in[52]) );
  GTECH_AND2 C7395 ( .A(N4301), .B(N4279), .Z(N4302) );
  GTECH_AND2 C7396 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4301) );
  GTECH_AND2 C7398 ( .A(N4304), .B(a3stg_fracadd[50]), .Z(
        a4stg_rnd_frac_pre3_in[51]) );
  GTECH_AND2 C7399 ( .A(N4303), .B(N4279), .Z(N4304) );
  GTECH_AND2 C7400 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4303) );
  GTECH_AND2 C7402 ( .A(N4306), .B(a3stg_fracadd[49]), .Z(
        a4stg_rnd_frac_pre3_in[50]) );
  GTECH_AND2 C7403 ( .A(N4305), .B(N4279), .Z(N4306) );
  GTECH_AND2 C7404 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4305) );
  GTECH_AND2 C7406 ( .A(N4308), .B(a3stg_fracadd[48]), .Z(
        a4stg_rnd_frac_pre3_in[49]) );
  GTECH_AND2 C7407 ( .A(N4307), .B(N4279), .Z(N4308) );
  GTECH_AND2 C7408 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4307) );
  GTECH_AND2 C7410 ( .A(N4310), .B(a3stg_fracadd[47]), .Z(
        a4stg_rnd_frac_pre3_in[48]) );
  GTECH_AND2 C7411 ( .A(N4309), .B(N4279), .Z(N4310) );
  GTECH_AND2 C7412 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4309) );
  GTECH_AND2 C7414 ( .A(N4312), .B(a3stg_fracadd[46]), .Z(
        a4stg_rnd_frac_pre3_in[47]) );
  GTECH_AND2 C7415 ( .A(N4311), .B(N4279), .Z(N4312) );
  GTECH_AND2 C7416 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4311) );
  GTECH_AND2 C7418 ( .A(N4314), .B(a3stg_fracadd[45]), .Z(
        a4stg_rnd_frac_pre3_in[46]) );
  GTECH_AND2 C7419 ( .A(N4313), .B(N4279), .Z(N4314) );
  GTECH_AND2 C7420 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4313) );
  GTECH_AND2 C7422 ( .A(N4316), .B(a3stg_fracadd[44]), .Z(
        a4stg_rnd_frac_pre3_in[45]) );
  GTECH_AND2 C7423 ( .A(N4315), .B(N4279), .Z(N4316) );
  GTECH_AND2 C7424 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4315) );
  GTECH_AND2 C7426 ( .A(N4318), .B(a3stg_fracadd[43]), .Z(
        a4stg_rnd_frac_pre3_in[44]) );
  GTECH_AND2 C7427 ( .A(N4317), .B(N4279), .Z(N4318) );
  GTECH_AND2 C7428 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4317) );
  GTECH_AND2 C7430 ( .A(N4320), .B(a3stg_fracadd[42]), .Z(
        a4stg_rnd_frac_pre3_in[43]) );
  GTECH_AND2 C7431 ( .A(N4319), .B(N4279), .Z(N4320) );
  GTECH_AND2 C7432 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4319) );
  GTECH_AND2 C7434 ( .A(N4322), .B(a3stg_fracadd[41]), .Z(
        a4stg_rnd_frac_pre3_in[42]) );
  GTECH_AND2 C7435 ( .A(N4321), .B(N4279), .Z(N4322) );
  GTECH_AND2 C7436 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4321) );
  GTECH_AND2 C7438 ( .A(N4324), .B(a3stg_fracadd[40]), .Z(
        a4stg_rnd_frac_pre3_in[41]) );
  GTECH_AND2 C7439 ( .A(N4323), .B(N4279), .Z(N4324) );
  GTECH_AND2 C7440 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4323) );
  GTECH_AND2 C7442 ( .A(N4326), .B(a3stg_fracadd[39]), .Z(
        a4stg_rnd_frac_pre3_in[40]) );
  GTECH_AND2 C7443 ( .A(N4325), .B(N4279), .Z(N4326) );
  GTECH_AND2 C7444 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4325) );
  GTECH_AND2 C7446 ( .A(N4328), .B(a3stg_fracadd[38]), .Z(
        a4stg_rnd_frac_pre3_in[39]) );
  GTECH_AND2 C7447 ( .A(N4327), .B(N4279), .Z(N4328) );
  GTECH_AND2 C7448 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4327) );
  GTECH_AND2 C7450 ( .A(N4330), .B(a3stg_fracadd[37]), .Z(
        a4stg_rnd_frac_pre3_in[38]) );
  GTECH_AND2 C7451 ( .A(N4329), .B(N4279), .Z(N4330) );
  GTECH_AND2 C7452 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4329) );
  GTECH_AND2 C7454 ( .A(N4332), .B(a3stg_fracadd[36]), .Z(
        a4stg_rnd_frac_pre3_in[37]) );
  GTECH_AND2 C7455 ( .A(N4331), .B(N4279), .Z(N4332) );
  GTECH_AND2 C7456 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4331) );
  GTECH_AND2 C7458 ( .A(N4334), .B(a3stg_fracadd[35]), .Z(
        a4stg_rnd_frac_pre3_in[36]) );
  GTECH_AND2 C7459 ( .A(N4333), .B(N4279), .Z(N4334) );
  GTECH_AND2 C7460 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4333) );
  GTECH_AND2 C7462 ( .A(N4336), .B(a3stg_fracadd[34]), .Z(
        a4stg_rnd_frac_pre3_in[35]) );
  GTECH_AND2 C7463 ( .A(N4335), .B(N4279), .Z(N4336) );
  GTECH_AND2 C7464 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4335) );
  GTECH_AND2 C7466 ( .A(N4338), .B(a3stg_fracadd[33]), .Z(
        a4stg_rnd_frac_pre3_in[34]) );
  GTECH_AND2 C7467 ( .A(N4337), .B(N4279), .Z(N4338) );
  GTECH_AND2 C7468 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4337) );
  GTECH_AND2 C7470 ( .A(N4340), .B(a3stg_fracadd[32]), .Z(
        a4stg_rnd_frac_pre3_in[33]) );
  GTECH_AND2 C7471 ( .A(N4339), .B(N4279), .Z(N4340) );
  GTECH_AND2 C7472 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4339) );
  GTECH_AND2 C7474 ( .A(N4342), .B(a3stg_fracadd[31]), .Z(
        a4stg_rnd_frac_pre3_in[32]) );
  GTECH_AND2 C7475 ( .A(N4341), .B(N4279), .Z(N4342) );
  GTECH_AND2 C7476 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4341) );
  GTECH_AND2 C7478 ( .A(N4344), .B(a3stg_fracadd[30]), .Z(
        a4stg_rnd_frac_pre3_in[31]) );
  GTECH_AND2 C7479 ( .A(N4343), .B(N4279), .Z(N4344) );
  GTECH_AND2 C7480 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4343) );
  GTECH_AND2 C7482 ( .A(N4346), .B(a3stg_fracadd[29]), .Z(
        a4stg_rnd_frac_pre3_in[30]) );
  GTECH_AND2 C7483 ( .A(N4345), .B(N4279), .Z(N4346) );
  GTECH_AND2 C7484 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4345) );
  GTECH_AND2 C7486 ( .A(N4348), .B(a3stg_fracadd[28]), .Z(
        a4stg_rnd_frac_pre3_in[29]) );
  GTECH_AND2 C7487 ( .A(N4347), .B(N4279), .Z(N4348) );
  GTECH_AND2 C7488 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4347) );
  GTECH_AND2 C7490 ( .A(N4350), .B(a3stg_fracadd[27]), .Z(
        a4stg_rnd_frac_pre3_in[28]) );
  GTECH_AND2 C7491 ( .A(N4349), .B(N4279), .Z(N4350) );
  GTECH_AND2 C7492 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4349) );
  GTECH_AND2 C7494 ( .A(N4352), .B(a3stg_fracadd[26]), .Z(
        a4stg_rnd_frac_pre3_in[27]) );
  GTECH_AND2 C7495 ( .A(N4351), .B(N4279), .Z(N4352) );
  GTECH_AND2 C7496 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4351) );
  GTECH_AND2 C7498 ( .A(N4354), .B(a3stg_fracadd[25]), .Z(
        a4stg_rnd_frac_pre3_in[26]) );
  GTECH_AND2 C7499 ( .A(N4353), .B(N4279), .Z(N4354) );
  GTECH_AND2 C7500 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4353) );
  GTECH_AND2 C7502 ( .A(N4356), .B(a3stg_fracadd[24]), .Z(
        a4stg_rnd_frac_pre3_in[25]) );
  GTECH_AND2 C7503 ( .A(N4355), .B(N4279), .Z(N4356) );
  GTECH_AND2 C7504 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4355) );
  GTECH_AND2 C7506 ( .A(N4358), .B(a3stg_fracadd[23]), .Z(
        a4stg_rnd_frac_pre3_in[24]) );
  GTECH_AND2 C7507 ( .A(N4357), .B(N4279), .Z(N4358) );
  GTECH_AND2 C7508 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4357) );
  GTECH_AND2 C7510 ( .A(N4360), .B(a3stg_fracadd[22]), .Z(
        a4stg_rnd_frac_pre3_in[23]) );
  GTECH_AND2 C7511 ( .A(N4359), .B(N4279), .Z(N4360) );
  GTECH_AND2 C7512 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4359) );
  GTECH_AND2 C7514 ( .A(N4362), .B(a3stg_fracadd[21]), .Z(
        a4stg_rnd_frac_pre3_in[22]) );
  GTECH_AND2 C7515 ( .A(N4361), .B(N4279), .Z(N4362) );
  GTECH_AND2 C7516 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4361) );
  GTECH_AND2 C7518 ( .A(N4364), .B(a3stg_fracadd[20]), .Z(
        a4stg_rnd_frac_pre3_in[21]) );
  GTECH_AND2 C7519 ( .A(N4363), .B(N4279), .Z(N4364) );
  GTECH_AND2 C7520 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4363) );
  GTECH_AND2 C7522 ( .A(N4366), .B(a3stg_fracadd[19]), .Z(
        a4stg_rnd_frac_pre3_in[20]) );
  GTECH_AND2 C7523 ( .A(N4365), .B(N4279), .Z(N4366) );
  GTECH_AND2 C7524 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4365) );
  GTECH_AND2 C7526 ( .A(N4368), .B(a3stg_fracadd[18]), .Z(
        a4stg_rnd_frac_pre3_in[19]) );
  GTECH_AND2 C7527 ( .A(N4367), .B(N4279), .Z(N4368) );
  GTECH_AND2 C7528 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4367) );
  GTECH_AND2 C7530 ( .A(N4370), .B(a3stg_fracadd[17]), .Z(
        a4stg_rnd_frac_pre3_in[18]) );
  GTECH_AND2 C7531 ( .A(N4369), .B(N4279), .Z(N4370) );
  GTECH_AND2 C7532 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4369) );
  GTECH_AND2 C7534 ( .A(N4372), .B(a3stg_fracadd[16]), .Z(
        a4stg_rnd_frac_pre3_in[17]) );
  GTECH_AND2 C7535 ( .A(N4371), .B(N4279), .Z(N4372) );
  GTECH_AND2 C7536 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4371) );
  GTECH_AND2 C7538 ( .A(N4374), .B(a3stg_fracadd[15]), .Z(
        a4stg_rnd_frac_pre3_in[16]) );
  GTECH_AND2 C7539 ( .A(N4373), .B(N4279), .Z(N4374) );
  GTECH_AND2 C7540 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4373) );
  GTECH_AND2 C7542 ( .A(N4376), .B(a3stg_fracadd[14]), .Z(
        a4stg_rnd_frac_pre3_in[15]) );
  GTECH_AND2 C7543 ( .A(N4375), .B(N4279), .Z(N4376) );
  GTECH_AND2 C7544 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4375) );
  GTECH_AND2 C7546 ( .A(N4378), .B(a3stg_fracadd[13]), .Z(
        a4stg_rnd_frac_pre3_in[14]) );
  GTECH_AND2 C7547 ( .A(N4377), .B(N4279), .Z(N4378) );
  GTECH_AND2 C7548 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4377) );
  GTECH_AND2 C7550 ( .A(N4380), .B(a3stg_fracadd[12]), .Z(
        a4stg_rnd_frac_pre3_in[13]) );
  GTECH_AND2 C7551 ( .A(N4379), .B(N4279), .Z(N4380) );
  GTECH_AND2 C7552 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4379) );
  GTECH_AND2 C7554 ( .A(N4382), .B(a3stg_fracadd[11]), .Z(
        a4stg_rnd_frac_pre3_in[12]) );
  GTECH_AND2 C7555 ( .A(N4381), .B(N4279), .Z(N4382) );
  GTECH_AND2 C7556 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4381) );
  GTECH_AND2 C7558 ( .A(N4384), .B(a3stg_fracadd[10]), .Z(
        a4stg_rnd_frac_pre3_in[11]) );
  GTECH_AND2 C7559 ( .A(N4383), .B(N4279), .Z(N4384) );
  GTECH_AND2 C7560 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4383) );
  GTECH_AND2 C7562 ( .A(N4386), .B(a3stg_fracadd[9]), .Z(
        a4stg_rnd_frac_pre3_in[10]) );
  GTECH_AND2 C7563 ( .A(N4385), .B(N4279), .Z(N4386) );
  GTECH_AND2 C7564 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4385) );
  GTECH_AND2 C7566 ( .A(N4388), .B(a3stg_fracadd[8]), .Z(
        a4stg_rnd_frac_pre3_in[9]) );
  GTECH_AND2 C7567 ( .A(N4387), .B(N4279), .Z(N4388) );
  GTECH_AND2 C7568 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4387) );
  GTECH_AND2 C7570 ( .A(N4390), .B(a3stg_fracadd[7]), .Z(
        a4stg_rnd_frac_pre3_in[8]) );
  GTECH_AND2 C7571 ( .A(N4389), .B(N4279), .Z(N4390) );
  GTECH_AND2 C7572 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4389) );
  GTECH_AND2 C7574 ( .A(N4392), .B(a3stg_fracadd[6]), .Z(
        a4stg_rnd_frac_pre3_in[7]) );
  GTECH_AND2 C7575 ( .A(N4391), .B(N4279), .Z(N4392) );
  GTECH_AND2 C7576 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4391) );
  GTECH_AND2 C7578 ( .A(N4394), .B(a3stg_fracadd[5]), .Z(
        a4stg_rnd_frac_pre3_in[6]) );
  GTECH_AND2 C7579 ( .A(N4393), .B(N4279), .Z(N4394) );
  GTECH_AND2 C7580 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4393) );
  GTECH_AND2 C7582 ( .A(N4396), .B(a3stg_fracadd[4]), .Z(
        a4stg_rnd_frac_pre3_in[5]) );
  GTECH_AND2 C7583 ( .A(N4395), .B(N4279), .Z(N4396) );
  GTECH_AND2 C7584 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4395) );
  GTECH_AND2 C7586 ( .A(N4398), .B(a3stg_fracadd[3]), .Z(
        a4stg_rnd_frac_pre3_in[4]) );
  GTECH_AND2 C7587 ( .A(N4397), .B(N4279), .Z(N4398) );
  GTECH_AND2 C7588 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4397) );
  GTECH_AND2 C7590 ( .A(N4400), .B(a3stg_fracadd[2]), .Z(
        a4stg_rnd_frac_pre3_in[3]) );
  GTECH_AND2 C7591 ( .A(N4399), .B(N4279), .Z(N4400) );
  GTECH_AND2 C7592 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4399) );
  GTECH_AND2 C7594 ( .A(N4402), .B(a3stg_fracadd[1]), .Z(
        a4stg_rnd_frac_pre3_in[2]) );
  GTECH_AND2 C7595 ( .A(N4401), .B(N4279), .Z(N4402) );
  GTECH_AND2 C7596 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4401) );
  GTECH_AND2 C7598 ( .A(N4404), .B(a3stg_fracadd[0]), .Z(
        a4stg_rnd_frac_pre3_in[1]) );
  GTECH_AND2 C7599 ( .A(N4403), .B(N4279), .Z(N4404) );
  GTECH_AND2 C7600 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4403) );
  GTECH_OR2 C7602 ( .A(N4420), .B(N4422), .Z(a4stg_rnd_frac_pre2_in[63]) );
  GTECH_OR2 C7603 ( .A(N4416), .B(N4419), .Z(N4420) );
  GTECH_OR2 C7604 ( .A(N4412), .B(N4415), .Z(N4416) );
  GTECH_OR2 C7605 ( .A(N4408), .B(N4411), .Z(N4412) );
  GTECH_AND2 C7606 ( .A(N4407), .B(a3stg_fracadd[63]), .Z(N4408) );
  GTECH_AND2 C7607 ( .A(N4405), .B(N4406), .Z(N4407) );
  GTECH_AND2 C7608 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4405) );
  GTECH_NOT I_753 ( .A(a3stg_inc_exp_inva), .Z(N4406) );
  GTECH_AND2 C7610 ( .A(N4410), .B(a3stg_fracadd[63]), .Z(N4411) );
  GTECH_AND2 C7611 ( .A(N4409), .B(a6stg_step), .Z(N4410) );
  GTECH_NOT I_754 ( .A(a4stg_rnd_frac_add_inv), .Z(N4409) );
  GTECH_AND2 C7613 ( .A(N4414), .B(a3stg_fracadd[62]), .Z(N4415) );
  GTECH_AND2 C7614 ( .A(N4413), .B(a6stg_step), .Z(N4414) );
  GTECH_NOT I_755 ( .A(a3stg_fdtos_inv), .Z(N4413) );
  GTECH_AND2 C7616 ( .A(N4418), .B(a4stg_shl[63]), .Z(N4419) );
  GTECH_AND2 C7617 ( .A(N4417), .B(a6stg_step), .Z(N4418) );
  GTECH_NOT I_756 ( .A(a4stg_fixtos_fxtod_inv), .Z(N4417) );
  GTECH_AND2 C7619 ( .A(N4421), .B(a4stg_rnd_frac_63), .Z(N4422) );
  GTECH_NOT I_757 ( .A(a6stg_step), .Z(N4421) );
  GTECH_OR2 C7621 ( .A(N4434), .B(N4436), .Z(a4stg_rnd_frac_pre2_in[62]) );
  GTECH_OR2 C7622 ( .A(N4431), .B(N4433), .Z(N4434) );
  GTECH_OR2 C7623 ( .A(N4428), .B(N4430), .Z(N4431) );
  GTECH_OR2 C7624 ( .A(N4425), .B(N4427), .Z(N4428) );
  GTECH_AND2 C7625 ( .A(N4424), .B(a3stg_fracadd[62]), .Z(N4425) );
  GTECH_AND2 C7626 ( .A(N4423), .B(N4406), .Z(N4424) );
  GTECH_AND2 C7627 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4423) );
  GTECH_AND2 C7629 ( .A(N4426), .B(a3stg_fracadd[62]), .Z(N4427) );
  GTECH_AND2 C7630 ( .A(N4409), .B(a6stg_step), .Z(N4426) );
  GTECH_AND2 C7632 ( .A(N4429), .B(a3stg_fracadd[61]), .Z(N4430) );
  GTECH_AND2 C7633 ( .A(N4413), .B(a6stg_step), .Z(N4429) );
  GTECH_AND2 C7635 ( .A(N4432), .B(a4stg_shl[62]), .Z(N4433) );
  GTECH_AND2 C7636 ( .A(N4417), .B(a6stg_step), .Z(N4432) );
  GTECH_AND2 C7638 ( .A(N4435), .B(a4stg_rnd_frac_62), .Z(N4436) );
  GTECH_NOT I_758 ( .A(a6stg_step), .Z(N4435) );
  GTECH_OR2 C7640 ( .A(N4448), .B(N4450), .Z(a4stg_rnd_frac_pre2_in[61]) );
  GTECH_OR2 C7641 ( .A(N4445), .B(N4447), .Z(N4448) );
  GTECH_OR2 C7642 ( .A(N4442), .B(N4444), .Z(N4445) );
  GTECH_OR2 C7643 ( .A(N4439), .B(N4441), .Z(N4442) );
  GTECH_AND2 C7644 ( .A(N4438), .B(a3stg_fracadd[61]), .Z(N4439) );
  GTECH_AND2 C7645 ( .A(N4437), .B(N4406), .Z(N4438) );
  GTECH_AND2 C7646 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4437) );
  GTECH_AND2 C7648 ( .A(N4440), .B(a3stg_fracadd[61]), .Z(N4441) );
  GTECH_AND2 C7649 ( .A(N4409), .B(a6stg_step), .Z(N4440) );
  GTECH_AND2 C7651 ( .A(N4443), .B(a3stg_fracadd[60]), .Z(N4444) );
  GTECH_AND2 C7652 ( .A(N4413), .B(a6stg_step), .Z(N4443) );
  GTECH_AND2 C7654 ( .A(N4446), .B(a4stg_shl[61]), .Z(N4447) );
  GTECH_AND2 C7655 ( .A(N4417), .B(a6stg_step), .Z(N4446) );
  GTECH_AND2 C7657 ( .A(N4449), .B(a4stg_rnd_frac_61), .Z(N4450) );
  GTECH_NOT I_759 ( .A(a6stg_step), .Z(N4449) );
  GTECH_OR2 C7659 ( .A(N4462), .B(N4464), .Z(a4stg_rnd_frac_pre2_in[60]) );
  GTECH_OR2 C7660 ( .A(N4459), .B(N4461), .Z(N4462) );
  GTECH_OR2 C7661 ( .A(N4456), .B(N4458), .Z(N4459) );
  GTECH_OR2 C7662 ( .A(N4453), .B(N4455), .Z(N4456) );
  GTECH_AND2 C7663 ( .A(N4452), .B(a3stg_fracadd[60]), .Z(N4453) );
  GTECH_AND2 C7664 ( .A(N4451), .B(N4406), .Z(N4452) );
  GTECH_AND2 C7665 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4451) );
  GTECH_AND2 C7667 ( .A(N4454), .B(a3stg_fracadd[60]), .Z(N4455) );
  GTECH_AND2 C7668 ( .A(N4409), .B(a6stg_step), .Z(N4454) );
  GTECH_AND2 C7670 ( .A(N4457), .B(a3stg_fracadd[59]), .Z(N4458) );
  GTECH_AND2 C7671 ( .A(N4413), .B(a6stg_step), .Z(N4457) );
  GTECH_AND2 C7673 ( .A(N4460), .B(a4stg_shl[60]), .Z(N4461) );
  GTECH_AND2 C7674 ( .A(N4417), .B(a6stg_step), .Z(N4460) );
  GTECH_AND2 C7676 ( .A(N4463), .B(a4stg_rnd_frac_60), .Z(N4464) );
  GTECH_NOT I_760 ( .A(a6stg_step), .Z(N4463) );
  GTECH_OR2 C7678 ( .A(N4476), .B(N4478), .Z(a4stg_rnd_frac_pre2_in[59]) );
  GTECH_OR2 C7679 ( .A(N4473), .B(N4475), .Z(N4476) );
  GTECH_OR2 C7680 ( .A(N4470), .B(N4472), .Z(N4473) );
  GTECH_OR2 C7681 ( .A(N4467), .B(N4469), .Z(N4470) );
  GTECH_AND2 C7682 ( .A(N4466), .B(a3stg_fracadd[59]), .Z(N4467) );
  GTECH_AND2 C7683 ( .A(N4465), .B(N4406), .Z(N4466) );
  GTECH_AND2 C7684 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4465) );
  GTECH_AND2 C7686 ( .A(N4468), .B(a3stg_fracadd[59]), .Z(N4469) );
  GTECH_AND2 C7687 ( .A(N4409), .B(a6stg_step), .Z(N4468) );
  GTECH_AND2 C7689 ( .A(N4471), .B(a3stg_fracadd[58]), .Z(N4472) );
  GTECH_AND2 C7690 ( .A(N4413), .B(a6stg_step), .Z(N4471) );
  GTECH_AND2 C7692 ( .A(N4474), .B(a4stg_shl[59]), .Z(N4475) );
  GTECH_AND2 C7693 ( .A(N4417), .B(a6stg_step), .Z(N4474) );
  GTECH_AND2 C7695 ( .A(N4477), .B(a4stg_rnd_frac_59), .Z(N4478) );
  GTECH_NOT I_761 ( .A(a6stg_step), .Z(N4477) );
  GTECH_OR2 C7697 ( .A(N4490), .B(N4492), .Z(a4stg_rnd_frac_pre2_in[58]) );
  GTECH_OR2 C7698 ( .A(N4487), .B(N4489), .Z(N4490) );
  GTECH_OR2 C7699 ( .A(N4484), .B(N4486), .Z(N4487) );
  GTECH_OR2 C7700 ( .A(N4481), .B(N4483), .Z(N4484) );
  GTECH_AND2 C7701 ( .A(N4480), .B(a3stg_fracadd[58]), .Z(N4481) );
  GTECH_AND2 C7702 ( .A(N4479), .B(N4406), .Z(N4480) );
  GTECH_AND2 C7703 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4479) );
  GTECH_AND2 C7705 ( .A(N4482), .B(a3stg_fracadd[58]), .Z(N4483) );
  GTECH_AND2 C7706 ( .A(N4409), .B(a6stg_step), .Z(N4482) );
  GTECH_AND2 C7708 ( .A(N4485), .B(a3stg_fracadd[57]), .Z(N4486) );
  GTECH_AND2 C7709 ( .A(N4413), .B(a6stg_step), .Z(N4485) );
  GTECH_AND2 C7711 ( .A(N4488), .B(a4stg_shl[58]), .Z(N4489) );
  GTECH_AND2 C7712 ( .A(N4417), .B(a6stg_step), .Z(N4488) );
  GTECH_AND2 C7714 ( .A(N4491), .B(a4stg_rnd_frac_58), .Z(N4492) );
  GTECH_NOT I_762 ( .A(a6stg_step), .Z(N4491) );
  GTECH_OR2 C7716 ( .A(N4504), .B(N4506), .Z(a4stg_rnd_frac_pre2_in[57]) );
  GTECH_OR2 C7717 ( .A(N4501), .B(N4503), .Z(N4504) );
  GTECH_OR2 C7718 ( .A(N4498), .B(N4500), .Z(N4501) );
  GTECH_OR2 C7719 ( .A(N4495), .B(N4497), .Z(N4498) );
  GTECH_AND2 C7720 ( .A(N4494), .B(a3stg_fracadd[57]), .Z(N4495) );
  GTECH_AND2 C7721 ( .A(N4493), .B(N4406), .Z(N4494) );
  GTECH_AND2 C7722 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4493) );
  GTECH_AND2 C7724 ( .A(N4496), .B(a3stg_fracadd[57]), .Z(N4497) );
  GTECH_AND2 C7725 ( .A(N4409), .B(a6stg_step), .Z(N4496) );
  GTECH_AND2 C7727 ( .A(N4499), .B(a3stg_fracadd[56]), .Z(N4500) );
  GTECH_AND2 C7728 ( .A(N4413), .B(a6stg_step), .Z(N4499) );
  GTECH_AND2 C7730 ( .A(N4502), .B(a4stg_shl[57]), .Z(N4503) );
  GTECH_AND2 C7731 ( .A(N4417), .B(a6stg_step), .Z(N4502) );
  GTECH_AND2 C7733 ( .A(N4505), .B(a4stg_rnd_frac_57), .Z(N4506) );
  GTECH_NOT I_763 ( .A(a6stg_step), .Z(N4505) );
  GTECH_OR2 C7735 ( .A(N4518), .B(N4520), .Z(a4stg_rnd_frac_pre2_in[56]) );
  GTECH_OR2 C7736 ( .A(N4515), .B(N4517), .Z(N4518) );
  GTECH_OR2 C7737 ( .A(N4512), .B(N4514), .Z(N4515) );
  GTECH_OR2 C7738 ( .A(N4509), .B(N4511), .Z(N4512) );
  GTECH_AND2 C7739 ( .A(N4508), .B(a3stg_fracadd[56]), .Z(N4509) );
  GTECH_AND2 C7740 ( .A(N4507), .B(N4406), .Z(N4508) );
  GTECH_AND2 C7741 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4507) );
  GTECH_AND2 C7743 ( .A(N4510), .B(a3stg_fracadd[56]), .Z(N4511) );
  GTECH_AND2 C7744 ( .A(N4409), .B(a6stg_step), .Z(N4510) );
  GTECH_AND2 C7746 ( .A(N4513), .B(a3stg_fracadd[55]), .Z(N4514) );
  GTECH_AND2 C7747 ( .A(N4413), .B(a6stg_step), .Z(N4513) );
  GTECH_AND2 C7749 ( .A(N4516), .B(a4stg_shl[56]), .Z(N4517) );
  GTECH_AND2 C7750 ( .A(N4417), .B(a6stg_step), .Z(N4516) );
  GTECH_AND2 C7752 ( .A(N4519), .B(a4stg_rnd_frac_56), .Z(N4520) );
  GTECH_NOT I_764 ( .A(a6stg_step), .Z(N4519) );
  GTECH_OR2 C7754 ( .A(N4532), .B(N4534), .Z(a4stg_rnd_frac_pre2_in[55]) );
  GTECH_OR2 C7755 ( .A(N4529), .B(N4531), .Z(N4532) );
  GTECH_OR2 C7756 ( .A(N4526), .B(N4528), .Z(N4529) );
  GTECH_OR2 C7757 ( .A(N4523), .B(N4525), .Z(N4526) );
  GTECH_AND2 C7758 ( .A(N4522), .B(a3stg_fracadd[55]), .Z(N4523) );
  GTECH_AND2 C7759 ( .A(N4521), .B(N4406), .Z(N4522) );
  GTECH_AND2 C7760 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4521) );
  GTECH_AND2 C7762 ( .A(N4524), .B(a3stg_fracadd[55]), .Z(N4525) );
  GTECH_AND2 C7763 ( .A(N4409), .B(a6stg_step), .Z(N4524) );
  GTECH_AND2 C7765 ( .A(N4527), .B(a3stg_fracadd[54]), .Z(N4528) );
  GTECH_AND2 C7766 ( .A(N4413), .B(a6stg_step), .Z(N4527) );
  GTECH_AND2 C7768 ( .A(N4530), .B(a4stg_shl[55]), .Z(N4531) );
  GTECH_AND2 C7769 ( .A(N4417), .B(a6stg_step), .Z(N4530) );
  GTECH_AND2 C7771 ( .A(N4533), .B(a4stg_rnd_frac_55), .Z(N4534) );
  GTECH_NOT I_765 ( .A(a6stg_step), .Z(N4533) );
  GTECH_OR2 C7773 ( .A(N4546), .B(N4548), .Z(a4stg_rnd_frac_pre2_in[54]) );
  GTECH_OR2 C7774 ( .A(N4543), .B(N4545), .Z(N4546) );
  GTECH_OR2 C7775 ( .A(N4540), .B(N4542), .Z(N4543) );
  GTECH_OR2 C7776 ( .A(N4537), .B(N4539), .Z(N4540) );
  GTECH_AND2 C7777 ( .A(N4536), .B(a3stg_fracadd[54]), .Z(N4537) );
  GTECH_AND2 C7778 ( .A(N4535), .B(N4406), .Z(N4536) );
  GTECH_AND2 C7779 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4535) );
  GTECH_AND2 C7781 ( .A(N4538), .B(a3stg_fracadd[54]), .Z(N4539) );
  GTECH_AND2 C7782 ( .A(N4409), .B(a6stg_step), .Z(N4538) );
  GTECH_AND2 C7784 ( .A(N4541), .B(a3stg_fracadd[53]), .Z(N4542) );
  GTECH_AND2 C7785 ( .A(N4413), .B(a6stg_step), .Z(N4541) );
  GTECH_AND2 C7787 ( .A(N4544), .B(a4stg_shl[54]), .Z(N4545) );
  GTECH_AND2 C7788 ( .A(N4417), .B(a6stg_step), .Z(N4544) );
  GTECH_AND2 C7790 ( .A(N4547), .B(a4stg_rnd_frac_54), .Z(N4548) );
  GTECH_NOT I_766 ( .A(a6stg_step), .Z(N4547) );
  GTECH_OR2 C7792 ( .A(N4560), .B(N4562), .Z(a4stg_rnd_frac_pre2_in[53]) );
  GTECH_OR2 C7793 ( .A(N4557), .B(N4559), .Z(N4560) );
  GTECH_OR2 C7794 ( .A(N4554), .B(N4556), .Z(N4557) );
  GTECH_OR2 C7795 ( .A(N4551), .B(N4553), .Z(N4554) );
  GTECH_AND2 C7796 ( .A(N4550), .B(a3stg_fracadd[53]), .Z(N4551) );
  GTECH_AND2 C7797 ( .A(N4549), .B(N4406), .Z(N4550) );
  GTECH_AND2 C7798 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4549) );
  GTECH_AND2 C7800 ( .A(N4552), .B(a3stg_fracadd[53]), .Z(N4553) );
  GTECH_AND2 C7801 ( .A(N4409), .B(a6stg_step), .Z(N4552) );
  GTECH_AND2 C7803 ( .A(N4555), .B(a3stg_fracadd[52]), .Z(N4556) );
  GTECH_AND2 C7804 ( .A(N4413), .B(a6stg_step), .Z(N4555) );
  GTECH_AND2 C7806 ( .A(N4558), .B(a4stg_shl[53]), .Z(N4559) );
  GTECH_AND2 C7807 ( .A(N4417), .B(a6stg_step), .Z(N4558) );
  GTECH_AND2 C7809 ( .A(N4561), .B(a4stg_rnd_frac_53), .Z(N4562) );
  GTECH_NOT I_767 ( .A(a6stg_step), .Z(N4561) );
  GTECH_OR2 C7811 ( .A(N4574), .B(N4576), .Z(a4stg_rnd_frac_pre2_in[52]) );
  GTECH_OR2 C7812 ( .A(N4571), .B(N4573), .Z(N4574) );
  GTECH_OR2 C7813 ( .A(N4568), .B(N4570), .Z(N4571) );
  GTECH_OR2 C7814 ( .A(N4565), .B(N4567), .Z(N4568) );
  GTECH_AND2 C7815 ( .A(N4564), .B(a3stg_fracadd[52]), .Z(N4565) );
  GTECH_AND2 C7816 ( .A(N4563), .B(N4406), .Z(N4564) );
  GTECH_AND2 C7817 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4563) );
  GTECH_AND2 C7819 ( .A(N4566), .B(a3stg_fracadd[52]), .Z(N4567) );
  GTECH_AND2 C7820 ( .A(N4409), .B(a6stg_step), .Z(N4566) );
  GTECH_AND2 C7822 ( .A(N4569), .B(a3stg_fracadd[51]), .Z(N4570) );
  GTECH_AND2 C7823 ( .A(N4413), .B(a6stg_step), .Z(N4569) );
  GTECH_AND2 C7825 ( .A(N4572), .B(a4stg_shl[52]), .Z(N4573) );
  GTECH_AND2 C7826 ( .A(N4417), .B(a6stg_step), .Z(N4572) );
  GTECH_AND2 C7828 ( .A(N4575), .B(a4stg_rnd_frac_52), .Z(N4576) );
  GTECH_NOT I_768 ( .A(a6stg_step), .Z(N4575) );
  GTECH_OR2 C7830 ( .A(N4588), .B(N4590), .Z(a4stg_rnd_frac_pre2_in[51]) );
  GTECH_OR2 C7831 ( .A(N4585), .B(N4587), .Z(N4588) );
  GTECH_OR2 C7832 ( .A(N4582), .B(N4584), .Z(N4585) );
  GTECH_OR2 C7833 ( .A(N4579), .B(N4581), .Z(N4582) );
  GTECH_AND2 C7834 ( .A(N4578), .B(a3stg_fracadd[51]), .Z(N4579) );
  GTECH_AND2 C7835 ( .A(N4577), .B(N4406), .Z(N4578) );
  GTECH_AND2 C7836 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4577) );
  GTECH_AND2 C7838 ( .A(N4580), .B(a3stg_fracadd[51]), .Z(N4581) );
  GTECH_AND2 C7839 ( .A(N4409), .B(a6stg_step), .Z(N4580) );
  GTECH_AND2 C7841 ( .A(N4583), .B(a3stg_fracadd[50]), .Z(N4584) );
  GTECH_AND2 C7842 ( .A(N4413), .B(a6stg_step), .Z(N4583) );
  GTECH_AND2 C7844 ( .A(N4586), .B(a4stg_shl[51]), .Z(N4587) );
  GTECH_AND2 C7845 ( .A(N4417), .B(a6stg_step), .Z(N4586) );
  GTECH_AND2 C7847 ( .A(N4589), .B(a4stg_rnd_frac_51), .Z(N4590) );
  GTECH_NOT I_769 ( .A(a6stg_step), .Z(N4589) );
  GTECH_OR2 C7849 ( .A(N4602), .B(N4604), .Z(a4stg_rnd_frac_pre2_in[50]) );
  GTECH_OR2 C7850 ( .A(N4599), .B(N4601), .Z(N4602) );
  GTECH_OR2 C7851 ( .A(N4596), .B(N4598), .Z(N4599) );
  GTECH_OR2 C7852 ( .A(N4593), .B(N4595), .Z(N4596) );
  GTECH_AND2 C7853 ( .A(N4592), .B(a3stg_fracadd[50]), .Z(N4593) );
  GTECH_AND2 C7854 ( .A(N4591), .B(N4406), .Z(N4592) );
  GTECH_AND2 C7855 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4591) );
  GTECH_AND2 C7857 ( .A(N4594), .B(a3stg_fracadd[50]), .Z(N4595) );
  GTECH_AND2 C7858 ( .A(N4409), .B(a6stg_step), .Z(N4594) );
  GTECH_AND2 C7860 ( .A(N4597), .B(a3stg_fracadd[49]), .Z(N4598) );
  GTECH_AND2 C7861 ( .A(N4413), .B(a6stg_step), .Z(N4597) );
  GTECH_AND2 C7863 ( .A(N4600), .B(a4stg_shl[50]), .Z(N4601) );
  GTECH_AND2 C7864 ( .A(N4417), .B(a6stg_step), .Z(N4600) );
  GTECH_AND2 C7866 ( .A(N4603), .B(a4stg_rnd_frac_50), .Z(N4604) );
  GTECH_NOT I_770 ( .A(a6stg_step), .Z(N4603) );
  GTECH_OR2 C7868 ( .A(N4616), .B(N4618), .Z(a4stg_rnd_frac_pre2_in[49]) );
  GTECH_OR2 C7869 ( .A(N4613), .B(N4615), .Z(N4616) );
  GTECH_OR2 C7870 ( .A(N4610), .B(N4612), .Z(N4613) );
  GTECH_OR2 C7871 ( .A(N4607), .B(N4609), .Z(N4610) );
  GTECH_AND2 C7872 ( .A(N4606), .B(a3stg_fracadd[49]), .Z(N4607) );
  GTECH_AND2 C7873 ( .A(N4605), .B(N4406), .Z(N4606) );
  GTECH_AND2 C7874 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4605) );
  GTECH_AND2 C7876 ( .A(N4608), .B(a3stg_fracadd[49]), .Z(N4609) );
  GTECH_AND2 C7877 ( .A(N4409), .B(a6stg_step), .Z(N4608) );
  GTECH_AND2 C7879 ( .A(N4611), .B(a3stg_fracadd[48]), .Z(N4612) );
  GTECH_AND2 C7880 ( .A(N4413), .B(a6stg_step), .Z(N4611) );
  GTECH_AND2 C7882 ( .A(N4614), .B(a4stg_shl[49]), .Z(N4615) );
  GTECH_AND2 C7883 ( .A(N4417), .B(a6stg_step), .Z(N4614) );
  GTECH_AND2 C7885 ( .A(N4617), .B(a4stg_rnd_frac_49), .Z(N4618) );
  GTECH_NOT I_771 ( .A(a6stg_step), .Z(N4617) );
  GTECH_OR2 C7887 ( .A(N4630), .B(N4632), .Z(a4stg_rnd_frac_pre2_in[48]) );
  GTECH_OR2 C7888 ( .A(N4627), .B(N4629), .Z(N4630) );
  GTECH_OR2 C7889 ( .A(N4624), .B(N4626), .Z(N4627) );
  GTECH_OR2 C7890 ( .A(N4621), .B(N4623), .Z(N4624) );
  GTECH_AND2 C7891 ( .A(N4620), .B(a3stg_fracadd[48]), .Z(N4621) );
  GTECH_AND2 C7892 ( .A(N4619), .B(N4406), .Z(N4620) );
  GTECH_AND2 C7893 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4619) );
  GTECH_AND2 C7895 ( .A(N4622), .B(a3stg_fracadd[48]), .Z(N4623) );
  GTECH_AND2 C7896 ( .A(N4409), .B(a6stg_step), .Z(N4622) );
  GTECH_AND2 C7898 ( .A(N4625), .B(a3stg_fracadd[47]), .Z(N4626) );
  GTECH_AND2 C7899 ( .A(N4413), .B(a6stg_step), .Z(N4625) );
  GTECH_AND2 C7901 ( .A(N4628), .B(a4stg_shl[48]), .Z(N4629) );
  GTECH_AND2 C7902 ( .A(N4417), .B(a6stg_step), .Z(N4628) );
  GTECH_AND2 C7904 ( .A(N4631), .B(a4stg_rnd_frac_48), .Z(N4632) );
  GTECH_NOT I_772 ( .A(a6stg_step), .Z(N4631) );
  GTECH_OR2 C7906 ( .A(N4644), .B(N4646), .Z(a4stg_rnd_frac_pre2_in[47]) );
  GTECH_OR2 C7907 ( .A(N4641), .B(N4643), .Z(N4644) );
  GTECH_OR2 C7908 ( .A(N4638), .B(N4640), .Z(N4641) );
  GTECH_OR2 C7909 ( .A(N4635), .B(N4637), .Z(N4638) );
  GTECH_AND2 C7910 ( .A(N4634), .B(a3stg_fracadd[47]), .Z(N4635) );
  GTECH_AND2 C7911 ( .A(N4633), .B(N4406), .Z(N4634) );
  GTECH_AND2 C7912 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4633) );
  GTECH_AND2 C7914 ( .A(N4636), .B(a3stg_fracadd[47]), .Z(N4637) );
  GTECH_AND2 C7915 ( .A(N4409), .B(a6stg_step), .Z(N4636) );
  GTECH_AND2 C7917 ( .A(N4639), .B(a3stg_fracadd[46]), .Z(N4640) );
  GTECH_AND2 C7918 ( .A(N4413), .B(a6stg_step), .Z(N4639) );
  GTECH_AND2 C7920 ( .A(N4642), .B(a4stg_shl[47]), .Z(N4643) );
  GTECH_AND2 C7921 ( .A(N4417), .B(a6stg_step), .Z(N4642) );
  GTECH_AND2 C7923 ( .A(N4645), .B(a4stg_rnd_frac_47), .Z(N4646) );
  GTECH_NOT I_773 ( .A(a6stg_step), .Z(N4645) );
  GTECH_OR2 C7925 ( .A(N4658), .B(N4660), .Z(a4stg_rnd_frac_pre2_in[46]) );
  GTECH_OR2 C7926 ( .A(N4655), .B(N4657), .Z(N4658) );
  GTECH_OR2 C7927 ( .A(N4652), .B(N4654), .Z(N4655) );
  GTECH_OR2 C7928 ( .A(N4649), .B(N4651), .Z(N4652) );
  GTECH_AND2 C7929 ( .A(N4648), .B(a3stg_fracadd[46]), .Z(N4649) );
  GTECH_AND2 C7930 ( .A(N4647), .B(N4406), .Z(N4648) );
  GTECH_AND2 C7931 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4647) );
  GTECH_AND2 C7933 ( .A(N4650), .B(a3stg_fracadd[46]), .Z(N4651) );
  GTECH_AND2 C7934 ( .A(N4409), .B(a6stg_step), .Z(N4650) );
  GTECH_AND2 C7936 ( .A(N4653), .B(a3stg_fracadd[45]), .Z(N4654) );
  GTECH_AND2 C7937 ( .A(N4413), .B(a6stg_step), .Z(N4653) );
  GTECH_AND2 C7939 ( .A(N4656), .B(a4stg_shl[46]), .Z(N4657) );
  GTECH_AND2 C7940 ( .A(N4417), .B(a6stg_step), .Z(N4656) );
  GTECH_AND2 C7942 ( .A(N4659), .B(a4stg_rnd_frac_46), .Z(N4660) );
  GTECH_NOT I_774 ( .A(a6stg_step), .Z(N4659) );
  GTECH_OR2 C7944 ( .A(N4672), .B(N4674), .Z(a4stg_rnd_frac_pre2_in[45]) );
  GTECH_OR2 C7945 ( .A(N4669), .B(N4671), .Z(N4672) );
  GTECH_OR2 C7946 ( .A(N4666), .B(N4668), .Z(N4669) );
  GTECH_OR2 C7947 ( .A(N4663), .B(N4665), .Z(N4666) );
  GTECH_AND2 C7948 ( .A(N4662), .B(a3stg_fracadd[45]), .Z(N4663) );
  GTECH_AND2 C7949 ( .A(N4661), .B(N4406), .Z(N4662) );
  GTECH_AND2 C7950 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4661) );
  GTECH_AND2 C7952 ( .A(N4664), .B(a3stg_fracadd[45]), .Z(N4665) );
  GTECH_AND2 C7953 ( .A(N4409), .B(a6stg_step), .Z(N4664) );
  GTECH_AND2 C7955 ( .A(N4667), .B(a3stg_fracadd[44]), .Z(N4668) );
  GTECH_AND2 C7956 ( .A(N4413), .B(a6stg_step), .Z(N4667) );
  GTECH_AND2 C7958 ( .A(N4670), .B(a4stg_shl[45]), .Z(N4671) );
  GTECH_AND2 C7959 ( .A(N4417), .B(a6stg_step), .Z(N4670) );
  GTECH_AND2 C7961 ( .A(N4673), .B(a4stg_rnd_frac_45), .Z(N4674) );
  GTECH_NOT I_775 ( .A(a6stg_step), .Z(N4673) );
  GTECH_OR2 C7963 ( .A(N4686), .B(N4688), .Z(a4stg_rnd_frac_pre2_in[44]) );
  GTECH_OR2 C7964 ( .A(N4683), .B(N4685), .Z(N4686) );
  GTECH_OR2 C7965 ( .A(N4680), .B(N4682), .Z(N4683) );
  GTECH_OR2 C7966 ( .A(N4677), .B(N4679), .Z(N4680) );
  GTECH_AND2 C7967 ( .A(N4676), .B(a3stg_fracadd[44]), .Z(N4677) );
  GTECH_AND2 C7968 ( .A(N4675), .B(N4406), .Z(N4676) );
  GTECH_AND2 C7969 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4675) );
  GTECH_AND2 C7971 ( .A(N4678), .B(a3stg_fracadd[44]), .Z(N4679) );
  GTECH_AND2 C7972 ( .A(N4409), .B(a6stg_step), .Z(N4678) );
  GTECH_AND2 C7974 ( .A(N4681), .B(a3stg_fracadd[43]), .Z(N4682) );
  GTECH_AND2 C7975 ( .A(N4413), .B(a6stg_step), .Z(N4681) );
  GTECH_AND2 C7977 ( .A(N4684), .B(a4stg_shl[44]), .Z(N4685) );
  GTECH_AND2 C7978 ( .A(N4417), .B(a6stg_step), .Z(N4684) );
  GTECH_AND2 C7980 ( .A(N4687), .B(a4stg_rnd_frac_44), .Z(N4688) );
  GTECH_NOT I_776 ( .A(a6stg_step), .Z(N4687) );
  GTECH_OR2 C7982 ( .A(N4700), .B(N4702), .Z(a4stg_rnd_frac_pre2_in[43]) );
  GTECH_OR2 C7983 ( .A(N4697), .B(N4699), .Z(N4700) );
  GTECH_OR2 C7984 ( .A(N4694), .B(N4696), .Z(N4697) );
  GTECH_OR2 C7985 ( .A(N4691), .B(N4693), .Z(N4694) );
  GTECH_AND2 C7986 ( .A(N4690), .B(a3stg_fracadd[43]), .Z(N4691) );
  GTECH_AND2 C7987 ( .A(N4689), .B(N4406), .Z(N4690) );
  GTECH_AND2 C7988 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4689) );
  GTECH_AND2 C7990 ( .A(N4692), .B(a3stg_fracadd[43]), .Z(N4693) );
  GTECH_AND2 C7991 ( .A(N4409), .B(a6stg_step), .Z(N4692) );
  GTECH_AND2 C7993 ( .A(N4695), .B(a3stg_fracadd[42]), .Z(N4696) );
  GTECH_AND2 C7994 ( .A(N4413), .B(a6stg_step), .Z(N4695) );
  GTECH_AND2 C7996 ( .A(N4698), .B(a4stg_shl[43]), .Z(N4699) );
  GTECH_AND2 C7997 ( .A(N4417), .B(a6stg_step), .Z(N4698) );
  GTECH_AND2 C7999 ( .A(N4701), .B(a4stg_rnd_frac_43), .Z(N4702) );
  GTECH_NOT I_777 ( .A(a6stg_step), .Z(N4701) );
  GTECH_OR2 C8001 ( .A(N4714), .B(N4716), .Z(a4stg_rnd_frac_pre2_in[42]) );
  GTECH_OR2 C8002 ( .A(N4711), .B(N4713), .Z(N4714) );
  GTECH_OR2 C8003 ( .A(N4708), .B(N4710), .Z(N4711) );
  GTECH_OR2 C8004 ( .A(N4705), .B(N4707), .Z(N4708) );
  GTECH_AND2 C8005 ( .A(N4704), .B(a3stg_fracadd[42]), .Z(N4705) );
  GTECH_AND2 C8006 ( .A(N4703), .B(N4406), .Z(N4704) );
  GTECH_AND2 C8007 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4703) );
  GTECH_AND2 C8009 ( .A(N4706), .B(a3stg_fracadd[42]), .Z(N4707) );
  GTECH_AND2 C8010 ( .A(N4409), .B(a6stg_step), .Z(N4706) );
  GTECH_AND2 C8012 ( .A(N4709), .B(a3stg_fracadd[41]), .Z(N4710) );
  GTECH_AND2 C8013 ( .A(N4413), .B(a6stg_step), .Z(N4709) );
  GTECH_AND2 C8015 ( .A(N4712), .B(a4stg_shl[42]), .Z(N4713) );
  GTECH_AND2 C8016 ( .A(N4417), .B(a6stg_step), .Z(N4712) );
  GTECH_AND2 C8018 ( .A(N4715), .B(a4stg_rnd_frac_42), .Z(N4716) );
  GTECH_NOT I_778 ( .A(a6stg_step), .Z(N4715) );
  GTECH_OR2 C8020 ( .A(N4728), .B(N4730), .Z(a4stg_rnd_frac_pre2_in[41]) );
  GTECH_OR2 C8021 ( .A(N4725), .B(N4727), .Z(N4728) );
  GTECH_OR2 C8022 ( .A(N4722), .B(N4724), .Z(N4725) );
  GTECH_OR2 C8023 ( .A(N4719), .B(N4721), .Z(N4722) );
  GTECH_AND2 C8024 ( .A(N4718), .B(a3stg_fracadd[41]), .Z(N4719) );
  GTECH_AND2 C8025 ( .A(N4717), .B(N4406), .Z(N4718) );
  GTECH_AND2 C8026 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4717) );
  GTECH_AND2 C8028 ( .A(N4720), .B(a3stg_fracadd[41]), .Z(N4721) );
  GTECH_AND2 C8029 ( .A(N4409), .B(a6stg_step), .Z(N4720) );
  GTECH_AND2 C8031 ( .A(N4723), .B(a3stg_fracadd[40]), .Z(N4724) );
  GTECH_AND2 C8032 ( .A(N4413), .B(a6stg_step), .Z(N4723) );
  GTECH_AND2 C8034 ( .A(N4726), .B(a4stg_shl[41]), .Z(N4727) );
  GTECH_AND2 C8035 ( .A(N4417), .B(a6stg_step), .Z(N4726) );
  GTECH_AND2 C8037 ( .A(N4729), .B(a4stg_rnd_frac_41), .Z(N4730) );
  GTECH_NOT I_779 ( .A(a6stg_step), .Z(N4729) );
  GTECH_OR2 C8039 ( .A(N4742), .B(N4744), .Z(a4stg_rnd_frac_pre2_in[40]) );
  GTECH_OR2 C8040 ( .A(N4739), .B(N4741), .Z(N4742) );
  GTECH_OR2 C8041 ( .A(N4736), .B(N4738), .Z(N4739) );
  GTECH_OR2 C8042 ( .A(N4733), .B(N4735), .Z(N4736) );
  GTECH_AND2 C8043 ( .A(N4732), .B(a3stg_fracadd[40]), .Z(N4733) );
  GTECH_AND2 C8044 ( .A(N4731), .B(N4406), .Z(N4732) );
  GTECH_AND2 C8045 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4731) );
  GTECH_AND2 C8047 ( .A(N4734), .B(a3stg_fracadd[40]), .Z(N4735) );
  GTECH_AND2 C8048 ( .A(N4409), .B(a6stg_step), .Z(N4734) );
  GTECH_AND2 C8050 ( .A(N4737), .B(a3stg_fracadd[39]), .Z(N4738) );
  GTECH_AND2 C8051 ( .A(N4413), .B(a6stg_step), .Z(N4737) );
  GTECH_AND2 C8053 ( .A(N4740), .B(a4stg_shl[40]), .Z(N4741) );
  GTECH_AND2 C8054 ( .A(N4417), .B(a6stg_step), .Z(N4740) );
  GTECH_AND2 C8056 ( .A(N4743), .B(a4stg_rnd_frac_40), .Z(N4744) );
  GTECH_NOT I_780 ( .A(a6stg_step), .Z(N4743) );
  GTECH_OR2 C8058 ( .A(N4756), .B(N4758), .Z(a4stg_rnd_frac_pre2_in[39]) );
  GTECH_OR2 C8059 ( .A(N4753), .B(N4755), .Z(N4756) );
  GTECH_OR2 C8060 ( .A(N4750), .B(N4752), .Z(N4753) );
  GTECH_OR2 C8061 ( .A(N4747), .B(N4749), .Z(N4750) );
  GTECH_AND2 C8062 ( .A(N4746), .B(a3stg_fracadd[39]), .Z(N4747) );
  GTECH_AND2 C8063 ( .A(N4745), .B(N4406), .Z(N4746) );
  GTECH_AND2 C8064 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4745) );
  GTECH_AND2 C8066 ( .A(N4748), .B(a3stg_fracadd[39]), .Z(N4749) );
  GTECH_AND2 C8067 ( .A(N4409), .B(a6stg_step), .Z(N4748) );
  GTECH_AND2 C8069 ( .A(N4751), .B(a3stg_fracadd[38]), .Z(N4752) );
  GTECH_AND2 C8070 ( .A(N4413), .B(a6stg_step), .Z(N4751) );
  GTECH_AND2 C8072 ( .A(N4754), .B(a4stg_shl[39]), .Z(N4755) );
  GTECH_AND2 C8073 ( .A(N4417), .B(a6stg_step), .Z(N4754) );
  GTECH_AND2 C8075 ( .A(N4757), .B(a4stg_rnd_frac_39), .Z(N4758) );
  GTECH_NOT I_781 ( .A(a6stg_step), .Z(N4757) );
  GTECH_OR2 C8077 ( .A(N4770), .B(N4772), .Z(a4stg_rnd_frac_pre2_in[38]) );
  GTECH_OR2 C8078 ( .A(N4767), .B(N4769), .Z(N4770) );
  GTECH_OR2 C8079 ( .A(N4764), .B(N4766), .Z(N4767) );
  GTECH_OR2 C8080 ( .A(N4761), .B(N4763), .Z(N4764) );
  GTECH_AND2 C8081 ( .A(N4760), .B(a3stg_fracadd[38]), .Z(N4761) );
  GTECH_AND2 C8082 ( .A(N4759), .B(N4406), .Z(N4760) );
  GTECH_AND2 C8083 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4759) );
  GTECH_AND2 C8085 ( .A(N4762), .B(a3stg_fracadd[38]), .Z(N4763) );
  GTECH_AND2 C8086 ( .A(N4409), .B(a6stg_step), .Z(N4762) );
  GTECH_AND2 C8088 ( .A(N4765), .B(a3stg_fracadd[37]), .Z(N4766) );
  GTECH_AND2 C8089 ( .A(N4413), .B(a6stg_step), .Z(N4765) );
  GTECH_AND2 C8091 ( .A(N4768), .B(a4stg_shl[38]), .Z(N4769) );
  GTECH_AND2 C8092 ( .A(N4417), .B(a6stg_step), .Z(N4768) );
  GTECH_AND2 C8094 ( .A(N4771), .B(a4stg_rnd_frac[38]), .Z(N4772) );
  GTECH_NOT I_782 ( .A(a6stg_step), .Z(N4771) );
  GTECH_OR2 C8096 ( .A(N4784), .B(N4786), .Z(a4stg_rnd_frac_pre2_in[37]) );
  GTECH_OR2 C8097 ( .A(N4781), .B(N4783), .Z(N4784) );
  GTECH_OR2 C8098 ( .A(N4778), .B(N4780), .Z(N4781) );
  GTECH_OR2 C8099 ( .A(N4775), .B(N4777), .Z(N4778) );
  GTECH_AND2 C8100 ( .A(N4774), .B(a3stg_fracadd[37]), .Z(N4775) );
  GTECH_AND2 C8101 ( .A(N4773), .B(N4406), .Z(N4774) );
  GTECH_AND2 C8102 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4773) );
  GTECH_AND2 C8104 ( .A(N4776), .B(a3stg_fracadd[37]), .Z(N4777) );
  GTECH_AND2 C8105 ( .A(N4409), .B(a6stg_step), .Z(N4776) );
  GTECH_AND2 C8107 ( .A(N4779), .B(a3stg_fracadd[36]), .Z(N4780) );
  GTECH_AND2 C8108 ( .A(N4413), .B(a6stg_step), .Z(N4779) );
  GTECH_AND2 C8110 ( .A(N4782), .B(a4stg_shl[37]), .Z(N4783) );
  GTECH_AND2 C8111 ( .A(N4417), .B(a6stg_step), .Z(N4782) );
  GTECH_AND2 C8113 ( .A(N4785), .B(a4stg_rnd_frac[37]), .Z(N4786) );
  GTECH_NOT I_783 ( .A(a6stg_step), .Z(N4785) );
  GTECH_OR2 C8115 ( .A(N4798), .B(N4800), .Z(a4stg_rnd_frac_pre2_in[36]) );
  GTECH_OR2 C8116 ( .A(N4795), .B(N4797), .Z(N4798) );
  GTECH_OR2 C8117 ( .A(N4792), .B(N4794), .Z(N4795) );
  GTECH_OR2 C8118 ( .A(N4789), .B(N4791), .Z(N4792) );
  GTECH_AND2 C8119 ( .A(N4788), .B(a3stg_fracadd[36]), .Z(N4789) );
  GTECH_AND2 C8120 ( .A(N4787), .B(N4406), .Z(N4788) );
  GTECH_AND2 C8121 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4787) );
  GTECH_AND2 C8123 ( .A(N4790), .B(a3stg_fracadd[36]), .Z(N4791) );
  GTECH_AND2 C8124 ( .A(N4409), .B(a6stg_step), .Z(N4790) );
  GTECH_AND2 C8126 ( .A(N4793), .B(a3stg_fracadd[35]), .Z(N4794) );
  GTECH_AND2 C8127 ( .A(N4413), .B(a6stg_step), .Z(N4793) );
  GTECH_AND2 C8129 ( .A(N4796), .B(a4stg_shl[36]), .Z(N4797) );
  GTECH_AND2 C8130 ( .A(N4417), .B(a6stg_step), .Z(N4796) );
  GTECH_AND2 C8132 ( .A(N4799), .B(a4stg_rnd_frac[36]), .Z(N4800) );
  GTECH_NOT I_784 ( .A(a6stg_step), .Z(N4799) );
  GTECH_OR2 C8134 ( .A(N4812), .B(N4814), .Z(a4stg_rnd_frac_pre2_in[35]) );
  GTECH_OR2 C8135 ( .A(N4809), .B(N4811), .Z(N4812) );
  GTECH_OR2 C8136 ( .A(N4806), .B(N4808), .Z(N4809) );
  GTECH_OR2 C8137 ( .A(N4803), .B(N4805), .Z(N4806) );
  GTECH_AND2 C8138 ( .A(N4802), .B(a3stg_fracadd[35]), .Z(N4803) );
  GTECH_AND2 C8139 ( .A(N4801), .B(N4406), .Z(N4802) );
  GTECH_AND2 C8140 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4801) );
  GTECH_AND2 C8142 ( .A(N4804), .B(a3stg_fracadd[35]), .Z(N4805) );
  GTECH_AND2 C8143 ( .A(N4409), .B(a6stg_step), .Z(N4804) );
  GTECH_AND2 C8145 ( .A(N4807), .B(a3stg_fracadd[34]), .Z(N4808) );
  GTECH_AND2 C8146 ( .A(N4413), .B(a6stg_step), .Z(N4807) );
  GTECH_AND2 C8148 ( .A(N4810), .B(a4stg_shl[35]), .Z(N4811) );
  GTECH_AND2 C8149 ( .A(N4417), .B(a6stg_step), .Z(N4810) );
  GTECH_AND2 C8151 ( .A(N4813), .B(a4stg_rnd_frac[35]), .Z(N4814) );
  GTECH_NOT I_785 ( .A(a6stg_step), .Z(N4813) );
  GTECH_OR2 C8153 ( .A(N4826), .B(N4828), .Z(a4stg_rnd_frac_pre2_in[34]) );
  GTECH_OR2 C8154 ( .A(N4823), .B(N4825), .Z(N4826) );
  GTECH_OR2 C8155 ( .A(N4820), .B(N4822), .Z(N4823) );
  GTECH_OR2 C8156 ( .A(N4817), .B(N4819), .Z(N4820) );
  GTECH_AND2 C8157 ( .A(N4816), .B(a3stg_fracadd[34]), .Z(N4817) );
  GTECH_AND2 C8158 ( .A(N4815), .B(N4406), .Z(N4816) );
  GTECH_AND2 C8159 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4815) );
  GTECH_AND2 C8161 ( .A(N4818), .B(a3stg_fracadd[34]), .Z(N4819) );
  GTECH_AND2 C8162 ( .A(N4409), .B(a6stg_step), .Z(N4818) );
  GTECH_AND2 C8164 ( .A(N4821), .B(a3stg_fracadd[33]), .Z(N4822) );
  GTECH_AND2 C8165 ( .A(N4413), .B(a6stg_step), .Z(N4821) );
  GTECH_AND2 C8167 ( .A(N4824), .B(a4stg_shl[34]), .Z(N4825) );
  GTECH_AND2 C8168 ( .A(N4417), .B(a6stg_step), .Z(N4824) );
  GTECH_AND2 C8170 ( .A(N4827), .B(a4stg_rnd_frac[34]), .Z(N4828) );
  GTECH_NOT I_786 ( .A(a6stg_step), .Z(N4827) );
  GTECH_OR2 C8172 ( .A(N4840), .B(N4842), .Z(a4stg_rnd_frac_pre2_in[33]) );
  GTECH_OR2 C8173 ( .A(N4837), .B(N4839), .Z(N4840) );
  GTECH_OR2 C8174 ( .A(N4834), .B(N4836), .Z(N4837) );
  GTECH_OR2 C8175 ( .A(N4831), .B(N4833), .Z(N4834) );
  GTECH_AND2 C8176 ( .A(N4830), .B(a3stg_fracadd[33]), .Z(N4831) );
  GTECH_AND2 C8177 ( .A(N4829), .B(N4406), .Z(N4830) );
  GTECH_AND2 C8178 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4829) );
  GTECH_AND2 C8180 ( .A(N4832), .B(a3stg_fracadd[33]), .Z(N4833) );
  GTECH_AND2 C8181 ( .A(N4409), .B(a6stg_step), .Z(N4832) );
  GTECH_AND2 C8183 ( .A(N4835), .B(a3stg_fracadd[32]), .Z(N4836) );
  GTECH_AND2 C8184 ( .A(N4413), .B(a6stg_step), .Z(N4835) );
  GTECH_AND2 C8186 ( .A(N4838), .B(a4stg_shl[33]), .Z(N4839) );
  GTECH_AND2 C8187 ( .A(N4417), .B(a6stg_step), .Z(N4838) );
  GTECH_AND2 C8189 ( .A(N4841), .B(a4stg_rnd_frac[33]), .Z(N4842) );
  GTECH_NOT I_787 ( .A(a6stg_step), .Z(N4841) );
  GTECH_OR2 C8191 ( .A(N4854), .B(N4856), .Z(a4stg_rnd_frac_pre2_in[32]) );
  GTECH_OR2 C8192 ( .A(N4851), .B(N4853), .Z(N4854) );
  GTECH_OR2 C8193 ( .A(N4848), .B(N4850), .Z(N4851) );
  GTECH_OR2 C8194 ( .A(N4845), .B(N4847), .Z(N4848) );
  GTECH_AND2 C8195 ( .A(N4844), .B(a3stg_fracadd[32]), .Z(N4845) );
  GTECH_AND2 C8196 ( .A(N4843), .B(N4406), .Z(N4844) );
  GTECH_AND2 C8197 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4843) );
  GTECH_AND2 C8199 ( .A(N4846), .B(a3stg_fracadd[32]), .Z(N4847) );
  GTECH_AND2 C8200 ( .A(N4409), .B(a6stg_step), .Z(N4846) );
  GTECH_AND2 C8202 ( .A(N4849), .B(a3stg_fracadd[31]), .Z(N4850) );
  GTECH_AND2 C8203 ( .A(N4413), .B(a6stg_step), .Z(N4849) );
  GTECH_AND2 C8205 ( .A(N4852), .B(a4stg_shl[32]), .Z(N4853) );
  GTECH_AND2 C8206 ( .A(N4417), .B(a6stg_step), .Z(N4852) );
  GTECH_AND2 C8208 ( .A(N4855), .B(a4stg_rnd_frac[32]), .Z(N4856) );
  GTECH_NOT I_788 ( .A(a6stg_step), .Z(N4855) );
  GTECH_OR2 C8210 ( .A(N4868), .B(N4870), .Z(a4stg_rnd_frac_pre2_in[31]) );
  GTECH_OR2 C8211 ( .A(N4865), .B(N4867), .Z(N4868) );
  GTECH_OR2 C8212 ( .A(N4862), .B(N4864), .Z(N4865) );
  GTECH_OR2 C8213 ( .A(N4859), .B(N4861), .Z(N4862) );
  GTECH_AND2 C8214 ( .A(N4858), .B(a3stg_fracadd[31]), .Z(N4859) );
  GTECH_AND2 C8215 ( .A(N4857), .B(N4406), .Z(N4858) );
  GTECH_AND2 C8216 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4857) );
  GTECH_AND2 C8218 ( .A(N4860), .B(a3stg_fracadd[31]), .Z(N4861) );
  GTECH_AND2 C8219 ( .A(N4409), .B(a6stg_step), .Z(N4860) );
  GTECH_AND2 C8221 ( .A(N4863), .B(a3stg_fracadd[30]), .Z(N4864) );
  GTECH_AND2 C8222 ( .A(N4413), .B(a6stg_step), .Z(N4863) );
  GTECH_AND2 C8224 ( .A(N4866), .B(a4stg_shl[31]), .Z(N4867) );
  GTECH_AND2 C8225 ( .A(N4417), .B(a6stg_step), .Z(N4866) );
  GTECH_AND2 C8227 ( .A(N4869), .B(a4stg_rnd_frac[31]), .Z(N4870) );
  GTECH_NOT I_789 ( .A(a6stg_step), .Z(N4869) );
  GTECH_OR2 C8229 ( .A(N4882), .B(N4884), .Z(a4stg_rnd_frac_pre2_in[30]) );
  GTECH_OR2 C8230 ( .A(N4879), .B(N4881), .Z(N4882) );
  GTECH_OR2 C8231 ( .A(N4876), .B(N4878), .Z(N4879) );
  GTECH_OR2 C8232 ( .A(N4873), .B(N4875), .Z(N4876) );
  GTECH_AND2 C8233 ( .A(N4872), .B(a3stg_fracadd[30]), .Z(N4873) );
  GTECH_AND2 C8234 ( .A(N4871), .B(N4406), .Z(N4872) );
  GTECH_AND2 C8235 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4871) );
  GTECH_AND2 C8237 ( .A(N4874), .B(a3stg_fracadd[30]), .Z(N4875) );
  GTECH_AND2 C8238 ( .A(N4409), .B(a6stg_step), .Z(N4874) );
  GTECH_AND2 C8240 ( .A(N4877), .B(a3stg_fracadd[29]), .Z(N4878) );
  GTECH_AND2 C8241 ( .A(N4413), .B(a6stg_step), .Z(N4877) );
  GTECH_AND2 C8243 ( .A(N4880), .B(a4stg_shl[30]), .Z(N4881) );
  GTECH_AND2 C8244 ( .A(N4417), .B(a6stg_step), .Z(N4880) );
  GTECH_AND2 C8246 ( .A(N4883), .B(a4stg_rnd_frac[30]), .Z(N4884) );
  GTECH_NOT I_790 ( .A(a6stg_step), .Z(N4883) );
  GTECH_OR2 C8248 ( .A(N4896), .B(N4898), .Z(a4stg_rnd_frac_pre2_in[29]) );
  GTECH_OR2 C8249 ( .A(N4893), .B(N4895), .Z(N4896) );
  GTECH_OR2 C8250 ( .A(N4890), .B(N4892), .Z(N4893) );
  GTECH_OR2 C8251 ( .A(N4887), .B(N4889), .Z(N4890) );
  GTECH_AND2 C8252 ( .A(N4886), .B(a3stg_fracadd[29]), .Z(N4887) );
  GTECH_AND2 C8253 ( .A(N4885), .B(N4406), .Z(N4886) );
  GTECH_AND2 C8254 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4885) );
  GTECH_AND2 C8256 ( .A(N4888), .B(a3stg_fracadd[29]), .Z(N4889) );
  GTECH_AND2 C8257 ( .A(N4409), .B(a6stg_step), .Z(N4888) );
  GTECH_AND2 C8259 ( .A(N4891), .B(a3stg_fracadd[28]), .Z(N4892) );
  GTECH_AND2 C8260 ( .A(N4413), .B(a6stg_step), .Z(N4891) );
  GTECH_AND2 C8262 ( .A(N4894), .B(a4stg_shl[29]), .Z(N4895) );
  GTECH_AND2 C8263 ( .A(N4417), .B(a6stg_step), .Z(N4894) );
  GTECH_AND2 C8265 ( .A(N4897), .B(a4stg_rnd_frac[29]), .Z(N4898) );
  GTECH_NOT I_791 ( .A(a6stg_step), .Z(N4897) );
  GTECH_OR2 C8267 ( .A(N4910), .B(N4912), .Z(a4stg_rnd_frac_pre2_in[28]) );
  GTECH_OR2 C8268 ( .A(N4907), .B(N4909), .Z(N4910) );
  GTECH_OR2 C8269 ( .A(N4904), .B(N4906), .Z(N4907) );
  GTECH_OR2 C8270 ( .A(N4901), .B(N4903), .Z(N4904) );
  GTECH_AND2 C8271 ( .A(N4900), .B(a3stg_fracadd[28]), .Z(N4901) );
  GTECH_AND2 C8272 ( .A(N4899), .B(N4406), .Z(N4900) );
  GTECH_AND2 C8273 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4899) );
  GTECH_AND2 C8275 ( .A(N4902), .B(a3stg_fracadd[28]), .Z(N4903) );
  GTECH_AND2 C8276 ( .A(N4409), .B(a6stg_step), .Z(N4902) );
  GTECH_AND2 C8278 ( .A(N4905), .B(a3stg_fracadd[27]), .Z(N4906) );
  GTECH_AND2 C8279 ( .A(N4413), .B(a6stg_step), .Z(N4905) );
  GTECH_AND2 C8281 ( .A(N4908), .B(a4stg_shl[28]), .Z(N4909) );
  GTECH_AND2 C8282 ( .A(N4417), .B(a6stg_step), .Z(N4908) );
  GTECH_AND2 C8284 ( .A(N4911), .B(a4stg_rnd_frac[28]), .Z(N4912) );
  GTECH_NOT I_792 ( .A(a6stg_step), .Z(N4911) );
  GTECH_OR2 C8286 ( .A(N4924), .B(N4926), .Z(a4stg_rnd_frac_pre2_in[27]) );
  GTECH_OR2 C8287 ( .A(N4921), .B(N4923), .Z(N4924) );
  GTECH_OR2 C8288 ( .A(N4918), .B(N4920), .Z(N4921) );
  GTECH_OR2 C8289 ( .A(N4915), .B(N4917), .Z(N4918) );
  GTECH_AND2 C8290 ( .A(N4914), .B(a3stg_fracadd[27]), .Z(N4915) );
  GTECH_AND2 C8291 ( .A(N4913), .B(N4406), .Z(N4914) );
  GTECH_AND2 C8292 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4913) );
  GTECH_AND2 C8294 ( .A(N4916), .B(a3stg_fracadd[27]), .Z(N4917) );
  GTECH_AND2 C8295 ( .A(N4409), .B(a6stg_step), .Z(N4916) );
  GTECH_AND2 C8297 ( .A(N4919), .B(a3stg_fracadd[26]), .Z(N4920) );
  GTECH_AND2 C8298 ( .A(N4413), .B(a6stg_step), .Z(N4919) );
  GTECH_AND2 C8300 ( .A(N4922), .B(a4stg_shl[27]), .Z(N4923) );
  GTECH_AND2 C8301 ( .A(N4417), .B(a6stg_step), .Z(N4922) );
  GTECH_AND2 C8303 ( .A(N4925), .B(a4stg_rnd_frac[27]), .Z(N4926) );
  GTECH_NOT I_793 ( .A(a6stg_step), .Z(N4925) );
  GTECH_OR2 C8305 ( .A(N4938), .B(N4940), .Z(a4stg_rnd_frac_pre2_in[26]) );
  GTECH_OR2 C8306 ( .A(N4935), .B(N4937), .Z(N4938) );
  GTECH_OR2 C8307 ( .A(N4932), .B(N4934), .Z(N4935) );
  GTECH_OR2 C8308 ( .A(N4929), .B(N4931), .Z(N4932) );
  GTECH_AND2 C8309 ( .A(N4928), .B(a3stg_fracadd[26]), .Z(N4929) );
  GTECH_AND2 C8310 ( .A(N4927), .B(N4406), .Z(N4928) );
  GTECH_AND2 C8311 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4927) );
  GTECH_AND2 C8313 ( .A(N4930), .B(a3stg_fracadd[26]), .Z(N4931) );
  GTECH_AND2 C8314 ( .A(N4409), .B(a6stg_step), .Z(N4930) );
  GTECH_AND2 C8316 ( .A(N4933), .B(a3stg_fracadd[25]), .Z(N4934) );
  GTECH_AND2 C8317 ( .A(N4413), .B(a6stg_step), .Z(N4933) );
  GTECH_AND2 C8319 ( .A(N4936), .B(a4stg_shl[26]), .Z(N4937) );
  GTECH_AND2 C8320 ( .A(N4417), .B(a6stg_step), .Z(N4936) );
  GTECH_AND2 C8322 ( .A(N4939), .B(a4stg_rnd_frac[26]), .Z(N4940) );
  GTECH_NOT I_794 ( .A(a6stg_step), .Z(N4939) );
  GTECH_OR2 C8324 ( .A(N4952), .B(N4954), .Z(a4stg_rnd_frac_pre2_in[25]) );
  GTECH_OR2 C8325 ( .A(N4949), .B(N4951), .Z(N4952) );
  GTECH_OR2 C8326 ( .A(N4946), .B(N4948), .Z(N4949) );
  GTECH_OR2 C8327 ( .A(N4943), .B(N4945), .Z(N4946) );
  GTECH_AND2 C8328 ( .A(N4942), .B(a3stg_fracadd[25]), .Z(N4943) );
  GTECH_AND2 C8329 ( .A(N4941), .B(N4406), .Z(N4942) );
  GTECH_AND2 C8330 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4941) );
  GTECH_AND2 C8332 ( .A(N4944), .B(a3stg_fracadd[25]), .Z(N4945) );
  GTECH_AND2 C8333 ( .A(N4409), .B(a6stg_step), .Z(N4944) );
  GTECH_AND2 C8335 ( .A(N4947), .B(a3stg_fracadd[24]), .Z(N4948) );
  GTECH_AND2 C8336 ( .A(N4413), .B(a6stg_step), .Z(N4947) );
  GTECH_AND2 C8338 ( .A(N4950), .B(a4stg_shl[25]), .Z(N4951) );
  GTECH_AND2 C8339 ( .A(N4417), .B(a6stg_step), .Z(N4950) );
  GTECH_AND2 C8341 ( .A(N4953), .B(a4stg_rnd_frac[25]), .Z(N4954) );
  GTECH_NOT I_795 ( .A(a6stg_step), .Z(N4953) );
  GTECH_OR2 C8343 ( .A(N4966), .B(N4968), .Z(a4stg_rnd_frac_pre2_in[24]) );
  GTECH_OR2 C8344 ( .A(N4963), .B(N4965), .Z(N4966) );
  GTECH_OR2 C8345 ( .A(N4960), .B(N4962), .Z(N4963) );
  GTECH_OR2 C8346 ( .A(N4957), .B(N4959), .Z(N4960) );
  GTECH_AND2 C8347 ( .A(N4956), .B(a3stg_fracadd[24]), .Z(N4957) );
  GTECH_AND2 C8348 ( .A(N4955), .B(N4406), .Z(N4956) );
  GTECH_AND2 C8349 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4955) );
  GTECH_AND2 C8351 ( .A(N4958), .B(a3stg_fracadd[24]), .Z(N4959) );
  GTECH_AND2 C8352 ( .A(N4409), .B(a6stg_step), .Z(N4958) );
  GTECH_AND2 C8354 ( .A(N4961), .B(a3stg_fracadd[23]), .Z(N4962) );
  GTECH_AND2 C8355 ( .A(N4413), .B(a6stg_step), .Z(N4961) );
  GTECH_AND2 C8357 ( .A(N4964), .B(a4stg_shl[24]), .Z(N4965) );
  GTECH_AND2 C8358 ( .A(N4417), .B(a6stg_step), .Z(N4964) );
  GTECH_AND2 C8360 ( .A(N4967), .B(a4stg_rnd_frac[24]), .Z(N4968) );
  GTECH_NOT I_796 ( .A(a6stg_step), .Z(N4967) );
  GTECH_OR2 C8362 ( .A(N4980), .B(N4982), .Z(a4stg_rnd_frac_pre2_in[23]) );
  GTECH_OR2 C8363 ( .A(N4977), .B(N4979), .Z(N4980) );
  GTECH_OR2 C8364 ( .A(N4974), .B(N4976), .Z(N4977) );
  GTECH_OR2 C8365 ( .A(N4971), .B(N4973), .Z(N4974) );
  GTECH_AND2 C8366 ( .A(N4970), .B(a3stg_fracadd[23]), .Z(N4971) );
  GTECH_AND2 C8367 ( .A(N4969), .B(N4406), .Z(N4970) );
  GTECH_AND2 C8368 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4969) );
  GTECH_AND2 C8370 ( .A(N4972), .B(a3stg_fracadd[23]), .Z(N4973) );
  GTECH_AND2 C8371 ( .A(N4409), .B(a6stg_step), .Z(N4972) );
  GTECH_AND2 C8373 ( .A(N4975), .B(a3stg_fracadd[22]), .Z(N4976) );
  GTECH_AND2 C8374 ( .A(N4413), .B(a6stg_step), .Z(N4975) );
  GTECH_AND2 C8376 ( .A(N4978), .B(a4stg_shl[23]), .Z(N4979) );
  GTECH_AND2 C8377 ( .A(N4417), .B(a6stg_step), .Z(N4978) );
  GTECH_AND2 C8379 ( .A(N4981), .B(a4stg_rnd_frac[23]), .Z(N4982) );
  GTECH_NOT I_797 ( .A(a6stg_step), .Z(N4981) );
  GTECH_OR2 C8381 ( .A(N4994), .B(N4996), .Z(a4stg_rnd_frac_pre2_in[22]) );
  GTECH_OR2 C8382 ( .A(N4991), .B(N4993), .Z(N4994) );
  GTECH_OR2 C8383 ( .A(N4988), .B(N4990), .Z(N4991) );
  GTECH_OR2 C8384 ( .A(N4985), .B(N4987), .Z(N4988) );
  GTECH_AND2 C8385 ( .A(N4984), .B(a3stg_fracadd[22]), .Z(N4985) );
  GTECH_AND2 C8386 ( .A(N4983), .B(N4406), .Z(N4984) );
  GTECH_AND2 C8387 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4983) );
  GTECH_AND2 C8389 ( .A(N4986), .B(a3stg_fracadd[22]), .Z(N4987) );
  GTECH_AND2 C8390 ( .A(N4409), .B(a6stg_step), .Z(N4986) );
  GTECH_AND2 C8392 ( .A(N4989), .B(a3stg_fracadd[21]), .Z(N4990) );
  GTECH_AND2 C8393 ( .A(N4413), .B(a6stg_step), .Z(N4989) );
  GTECH_AND2 C8395 ( .A(N4992), .B(a4stg_shl[22]), .Z(N4993) );
  GTECH_AND2 C8396 ( .A(N4417), .B(a6stg_step), .Z(N4992) );
  GTECH_AND2 C8398 ( .A(N4995), .B(a4stg_rnd_frac[22]), .Z(N4996) );
  GTECH_NOT I_798 ( .A(a6stg_step), .Z(N4995) );
  GTECH_OR2 C8400 ( .A(N5008), .B(N5010), .Z(a4stg_rnd_frac_pre2_in[21]) );
  GTECH_OR2 C8401 ( .A(N5005), .B(N5007), .Z(N5008) );
  GTECH_OR2 C8402 ( .A(N5002), .B(N5004), .Z(N5005) );
  GTECH_OR2 C8403 ( .A(N4999), .B(N5001), .Z(N5002) );
  GTECH_AND2 C8404 ( .A(N4998), .B(a3stg_fracadd[21]), .Z(N4999) );
  GTECH_AND2 C8405 ( .A(N4997), .B(N4406), .Z(N4998) );
  GTECH_AND2 C8406 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N4997) );
  GTECH_AND2 C8408 ( .A(N5000), .B(a3stg_fracadd[21]), .Z(N5001) );
  GTECH_AND2 C8409 ( .A(N4409), .B(a6stg_step), .Z(N5000) );
  GTECH_AND2 C8411 ( .A(N5003), .B(a3stg_fracadd[20]), .Z(N5004) );
  GTECH_AND2 C8412 ( .A(N4413), .B(a6stg_step), .Z(N5003) );
  GTECH_AND2 C8414 ( .A(N5006), .B(a4stg_shl[21]), .Z(N5007) );
  GTECH_AND2 C8415 ( .A(N4417), .B(a6stg_step), .Z(N5006) );
  GTECH_AND2 C8417 ( .A(N5009), .B(a4stg_rnd_frac[21]), .Z(N5010) );
  GTECH_NOT I_799 ( .A(a6stg_step), .Z(N5009) );
  GTECH_OR2 C8419 ( .A(N5022), .B(N5024), .Z(a4stg_rnd_frac_pre2_in[20]) );
  GTECH_OR2 C8420 ( .A(N5019), .B(N5021), .Z(N5022) );
  GTECH_OR2 C8421 ( .A(N5016), .B(N5018), .Z(N5019) );
  GTECH_OR2 C8422 ( .A(N5013), .B(N5015), .Z(N5016) );
  GTECH_AND2 C8423 ( .A(N5012), .B(a3stg_fracadd[20]), .Z(N5013) );
  GTECH_AND2 C8424 ( .A(N5011), .B(N4406), .Z(N5012) );
  GTECH_AND2 C8425 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5011) );
  GTECH_AND2 C8427 ( .A(N5014), .B(a3stg_fracadd[20]), .Z(N5015) );
  GTECH_AND2 C8428 ( .A(N4409), .B(a6stg_step), .Z(N5014) );
  GTECH_AND2 C8430 ( .A(N5017), .B(a3stg_fracadd[19]), .Z(N5018) );
  GTECH_AND2 C8431 ( .A(N4413), .B(a6stg_step), .Z(N5017) );
  GTECH_AND2 C8433 ( .A(N5020), .B(a4stg_shl[20]), .Z(N5021) );
  GTECH_AND2 C8434 ( .A(N4417), .B(a6stg_step), .Z(N5020) );
  GTECH_AND2 C8436 ( .A(N5023), .B(a4stg_rnd_frac[20]), .Z(N5024) );
  GTECH_NOT I_800 ( .A(a6stg_step), .Z(N5023) );
  GTECH_OR2 C8438 ( .A(N5036), .B(N5038), .Z(a4stg_rnd_frac_pre2_in[19]) );
  GTECH_OR2 C8439 ( .A(N5033), .B(N5035), .Z(N5036) );
  GTECH_OR2 C8440 ( .A(N5030), .B(N5032), .Z(N5033) );
  GTECH_OR2 C8441 ( .A(N5027), .B(N5029), .Z(N5030) );
  GTECH_AND2 C8442 ( .A(N5026), .B(a3stg_fracadd[19]), .Z(N5027) );
  GTECH_AND2 C8443 ( .A(N5025), .B(N4406), .Z(N5026) );
  GTECH_AND2 C8444 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5025) );
  GTECH_AND2 C8446 ( .A(N5028), .B(a3stg_fracadd[19]), .Z(N5029) );
  GTECH_AND2 C8447 ( .A(N4409), .B(a6stg_step), .Z(N5028) );
  GTECH_AND2 C8449 ( .A(N5031), .B(a3stg_fracadd[18]), .Z(N5032) );
  GTECH_AND2 C8450 ( .A(N4413), .B(a6stg_step), .Z(N5031) );
  GTECH_AND2 C8452 ( .A(N5034), .B(a4stg_shl[19]), .Z(N5035) );
  GTECH_AND2 C8453 ( .A(N4417), .B(a6stg_step), .Z(N5034) );
  GTECH_AND2 C8455 ( .A(N5037), .B(a4stg_rnd_frac[19]), .Z(N5038) );
  GTECH_NOT I_801 ( .A(a6stg_step), .Z(N5037) );
  GTECH_OR2 C8457 ( .A(N5050), .B(N5052), .Z(a4stg_rnd_frac_pre2_in[18]) );
  GTECH_OR2 C8458 ( .A(N5047), .B(N5049), .Z(N5050) );
  GTECH_OR2 C8459 ( .A(N5044), .B(N5046), .Z(N5047) );
  GTECH_OR2 C8460 ( .A(N5041), .B(N5043), .Z(N5044) );
  GTECH_AND2 C8461 ( .A(N5040), .B(a3stg_fracadd[18]), .Z(N5041) );
  GTECH_AND2 C8462 ( .A(N5039), .B(N4406), .Z(N5040) );
  GTECH_AND2 C8463 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5039) );
  GTECH_AND2 C8465 ( .A(N5042), .B(a3stg_fracadd[18]), .Z(N5043) );
  GTECH_AND2 C8466 ( .A(N4409), .B(a6stg_step), .Z(N5042) );
  GTECH_AND2 C8468 ( .A(N5045), .B(a3stg_fracadd[17]), .Z(N5046) );
  GTECH_AND2 C8469 ( .A(N4413), .B(a6stg_step), .Z(N5045) );
  GTECH_AND2 C8471 ( .A(N5048), .B(a4stg_shl[18]), .Z(N5049) );
  GTECH_AND2 C8472 ( .A(N4417), .B(a6stg_step), .Z(N5048) );
  GTECH_AND2 C8474 ( .A(N5051), .B(a4stg_rnd_frac[18]), .Z(N5052) );
  GTECH_NOT I_802 ( .A(a6stg_step), .Z(N5051) );
  GTECH_OR2 C8476 ( .A(N5064), .B(N5066), .Z(a4stg_rnd_frac_pre2_in[17]) );
  GTECH_OR2 C8477 ( .A(N5061), .B(N5063), .Z(N5064) );
  GTECH_OR2 C8478 ( .A(N5058), .B(N5060), .Z(N5061) );
  GTECH_OR2 C8479 ( .A(N5055), .B(N5057), .Z(N5058) );
  GTECH_AND2 C8480 ( .A(N5054), .B(a3stg_fracadd[17]), .Z(N5055) );
  GTECH_AND2 C8481 ( .A(N5053), .B(N4406), .Z(N5054) );
  GTECH_AND2 C8482 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5053) );
  GTECH_AND2 C8484 ( .A(N5056), .B(a3stg_fracadd[17]), .Z(N5057) );
  GTECH_AND2 C8485 ( .A(N4409), .B(a6stg_step), .Z(N5056) );
  GTECH_AND2 C8487 ( .A(N5059), .B(a3stg_fracadd[16]), .Z(N5060) );
  GTECH_AND2 C8488 ( .A(N4413), .B(a6stg_step), .Z(N5059) );
  GTECH_AND2 C8490 ( .A(N5062), .B(a4stg_shl[17]), .Z(N5063) );
  GTECH_AND2 C8491 ( .A(N4417), .B(a6stg_step), .Z(N5062) );
  GTECH_AND2 C8493 ( .A(N5065), .B(a4stg_rnd_frac[17]), .Z(N5066) );
  GTECH_NOT I_803 ( .A(a6stg_step), .Z(N5065) );
  GTECH_OR2 C8495 ( .A(N5078), .B(N5080), .Z(a4stg_rnd_frac_pre2_in[16]) );
  GTECH_OR2 C8496 ( .A(N5075), .B(N5077), .Z(N5078) );
  GTECH_OR2 C8497 ( .A(N5072), .B(N5074), .Z(N5075) );
  GTECH_OR2 C8498 ( .A(N5069), .B(N5071), .Z(N5072) );
  GTECH_AND2 C8499 ( .A(N5068), .B(a3stg_fracadd[16]), .Z(N5069) );
  GTECH_AND2 C8500 ( .A(N5067), .B(N4406), .Z(N5068) );
  GTECH_AND2 C8501 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5067) );
  GTECH_AND2 C8503 ( .A(N5070), .B(a3stg_fracadd[16]), .Z(N5071) );
  GTECH_AND2 C8504 ( .A(N4409), .B(a6stg_step), .Z(N5070) );
  GTECH_AND2 C8506 ( .A(N5073), .B(a3stg_fracadd[15]), .Z(N5074) );
  GTECH_AND2 C8507 ( .A(N4413), .B(a6stg_step), .Z(N5073) );
  GTECH_AND2 C8509 ( .A(N5076), .B(a4stg_shl[16]), .Z(N5077) );
  GTECH_AND2 C8510 ( .A(N4417), .B(a6stg_step), .Z(N5076) );
  GTECH_AND2 C8512 ( .A(N5079), .B(a4stg_rnd_frac[16]), .Z(N5080) );
  GTECH_NOT I_804 ( .A(a6stg_step), .Z(N5079) );
  GTECH_OR2 C8514 ( .A(N5092), .B(N5094), .Z(a4stg_rnd_frac_pre2_in[15]) );
  GTECH_OR2 C8515 ( .A(N5089), .B(N5091), .Z(N5092) );
  GTECH_OR2 C8516 ( .A(N5086), .B(N5088), .Z(N5089) );
  GTECH_OR2 C8517 ( .A(N5083), .B(N5085), .Z(N5086) );
  GTECH_AND2 C8518 ( .A(N5082), .B(a3stg_fracadd[15]), .Z(N5083) );
  GTECH_AND2 C8519 ( .A(N5081), .B(N4406), .Z(N5082) );
  GTECH_AND2 C8520 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5081) );
  GTECH_AND2 C8522 ( .A(N5084), .B(a3stg_fracadd[15]), .Z(N5085) );
  GTECH_AND2 C8523 ( .A(N4409), .B(a6stg_step), .Z(N5084) );
  GTECH_AND2 C8525 ( .A(N5087), .B(a3stg_fracadd[14]), .Z(N5088) );
  GTECH_AND2 C8526 ( .A(N4413), .B(a6stg_step), .Z(N5087) );
  GTECH_AND2 C8528 ( .A(N5090), .B(a4stg_shl[15]), .Z(N5091) );
  GTECH_AND2 C8529 ( .A(N4417), .B(a6stg_step), .Z(N5090) );
  GTECH_AND2 C8531 ( .A(N5093), .B(a4stg_rnd_frac[15]), .Z(N5094) );
  GTECH_NOT I_805 ( .A(a6stg_step), .Z(N5093) );
  GTECH_OR2 C8533 ( .A(N5106), .B(N5108), .Z(a4stg_rnd_frac_pre2_in[14]) );
  GTECH_OR2 C8534 ( .A(N5103), .B(N5105), .Z(N5106) );
  GTECH_OR2 C8535 ( .A(N5100), .B(N5102), .Z(N5103) );
  GTECH_OR2 C8536 ( .A(N5097), .B(N5099), .Z(N5100) );
  GTECH_AND2 C8537 ( .A(N5096), .B(a3stg_fracadd[14]), .Z(N5097) );
  GTECH_AND2 C8538 ( .A(N5095), .B(N4406), .Z(N5096) );
  GTECH_AND2 C8539 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5095) );
  GTECH_AND2 C8541 ( .A(N5098), .B(a3stg_fracadd[14]), .Z(N5099) );
  GTECH_AND2 C8542 ( .A(N4409), .B(a6stg_step), .Z(N5098) );
  GTECH_AND2 C8544 ( .A(N5101), .B(a3stg_fracadd[13]), .Z(N5102) );
  GTECH_AND2 C8545 ( .A(N4413), .B(a6stg_step), .Z(N5101) );
  GTECH_AND2 C8547 ( .A(N5104), .B(a4stg_shl[14]), .Z(N5105) );
  GTECH_AND2 C8548 ( .A(N4417), .B(a6stg_step), .Z(N5104) );
  GTECH_AND2 C8550 ( .A(N5107), .B(a4stg_rnd_frac[14]), .Z(N5108) );
  GTECH_NOT I_806 ( .A(a6stg_step), .Z(N5107) );
  GTECH_OR2 C8552 ( .A(N5120), .B(N5122), .Z(a4stg_rnd_frac_pre2_in[13]) );
  GTECH_OR2 C8553 ( .A(N5117), .B(N5119), .Z(N5120) );
  GTECH_OR2 C8554 ( .A(N5114), .B(N5116), .Z(N5117) );
  GTECH_OR2 C8555 ( .A(N5111), .B(N5113), .Z(N5114) );
  GTECH_AND2 C8556 ( .A(N5110), .B(a3stg_fracadd[13]), .Z(N5111) );
  GTECH_AND2 C8557 ( .A(N5109), .B(N4406), .Z(N5110) );
  GTECH_AND2 C8558 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5109) );
  GTECH_AND2 C8560 ( .A(N5112), .B(a3stg_fracadd[13]), .Z(N5113) );
  GTECH_AND2 C8561 ( .A(N4409), .B(a6stg_step), .Z(N5112) );
  GTECH_AND2 C8563 ( .A(N5115), .B(a3stg_fracadd[12]), .Z(N5116) );
  GTECH_AND2 C8564 ( .A(N4413), .B(a6stg_step), .Z(N5115) );
  GTECH_AND2 C8566 ( .A(N5118), .B(a4stg_shl[13]), .Z(N5119) );
  GTECH_AND2 C8567 ( .A(N4417), .B(a6stg_step), .Z(N5118) );
  GTECH_AND2 C8569 ( .A(N5121), .B(a4stg_rnd_frac[13]), .Z(N5122) );
  GTECH_NOT I_807 ( .A(a6stg_step), .Z(N5121) );
  GTECH_OR2 C8571 ( .A(N5134), .B(N5136), .Z(a4stg_rnd_frac_pre2_in[12]) );
  GTECH_OR2 C8572 ( .A(N5131), .B(N5133), .Z(N5134) );
  GTECH_OR2 C8573 ( .A(N5128), .B(N5130), .Z(N5131) );
  GTECH_OR2 C8574 ( .A(N5125), .B(N5127), .Z(N5128) );
  GTECH_AND2 C8575 ( .A(N5124), .B(a3stg_fracadd[12]), .Z(N5125) );
  GTECH_AND2 C8576 ( .A(N5123), .B(N4406), .Z(N5124) );
  GTECH_AND2 C8577 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5123) );
  GTECH_AND2 C8579 ( .A(N5126), .B(a3stg_fracadd[12]), .Z(N5127) );
  GTECH_AND2 C8580 ( .A(N4409), .B(a6stg_step), .Z(N5126) );
  GTECH_AND2 C8582 ( .A(N5129), .B(a3stg_fracadd[11]), .Z(N5130) );
  GTECH_AND2 C8583 ( .A(N4413), .B(a6stg_step), .Z(N5129) );
  GTECH_AND2 C8585 ( .A(N5132), .B(a4stg_shl[12]), .Z(N5133) );
  GTECH_AND2 C8586 ( .A(N4417), .B(a6stg_step), .Z(N5132) );
  GTECH_AND2 C8588 ( .A(N5135), .B(a4stg_rnd_frac[12]), .Z(N5136) );
  GTECH_NOT I_808 ( .A(a6stg_step), .Z(N5135) );
  GTECH_OR2 C8590 ( .A(N5148), .B(N5150), .Z(a4stg_rnd_frac_pre2_in[11]) );
  GTECH_OR2 C8591 ( .A(N5145), .B(N5147), .Z(N5148) );
  GTECH_OR2 C8592 ( .A(N5142), .B(N5144), .Z(N5145) );
  GTECH_OR2 C8593 ( .A(N5139), .B(N5141), .Z(N5142) );
  GTECH_AND2 C8594 ( .A(N5138), .B(a3stg_fracadd[11]), .Z(N5139) );
  GTECH_AND2 C8595 ( .A(N5137), .B(N4406), .Z(N5138) );
  GTECH_AND2 C8596 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5137) );
  GTECH_AND2 C8598 ( .A(N5140), .B(a3stg_fracadd[11]), .Z(N5141) );
  GTECH_AND2 C8599 ( .A(N4409), .B(a6stg_step), .Z(N5140) );
  GTECH_AND2 C8601 ( .A(N5143), .B(a3stg_fracadd[10]), .Z(N5144) );
  GTECH_AND2 C8602 ( .A(N4413), .B(a6stg_step), .Z(N5143) );
  GTECH_AND2 C8604 ( .A(N5146), .B(a4stg_shl[11]), .Z(N5147) );
  GTECH_AND2 C8605 ( .A(N4417), .B(a6stg_step), .Z(N5146) );
  GTECH_AND2 C8607 ( .A(N5149), .B(a4stg_rnd_frac_11), .Z(N5150) );
  GTECH_NOT I_809 ( .A(a6stg_step), .Z(N5149) );
  GTECH_OR2 C8609 ( .A(N5162), .B(N5164), .Z(a4stg_rnd_frac_pre2_in[10]) );
  GTECH_OR2 C8610 ( .A(N5159), .B(N5161), .Z(N5162) );
  GTECH_OR2 C8611 ( .A(N5156), .B(N5158), .Z(N5159) );
  GTECH_OR2 C8612 ( .A(N5153), .B(N5155), .Z(N5156) );
  GTECH_AND2 C8613 ( .A(N5152), .B(a3stg_fracadd[10]), .Z(N5153) );
  GTECH_AND2 C8614 ( .A(N5151), .B(N4406), .Z(N5152) );
  GTECH_AND2 C8615 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5151) );
  GTECH_AND2 C8617 ( .A(N5154), .B(a3stg_fracadd[10]), .Z(N5155) );
  GTECH_AND2 C8618 ( .A(N4409), .B(a6stg_step), .Z(N5154) );
  GTECH_AND2 C8620 ( .A(N5157), .B(a3stg_fracadd[9]), .Z(N5158) );
  GTECH_AND2 C8621 ( .A(N4413), .B(a6stg_step), .Z(N5157) );
  GTECH_AND2 C8623 ( .A(N5160), .B(a4stg_shl[10]), .Z(N5161) );
  GTECH_AND2 C8624 ( .A(N4417), .B(a6stg_step), .Z(N5160) );
  GTECH_AND2 C8626 ( .A(N5163), .B(a4stg_rnd_frac_10), .Z(N5164) );
  GTECH_NOT I_810 ( .A(a6stg_step), .Z(N5163) );
  GTECH_OR2 C8628 ( .A(N5176), .B(N5178), .Z(a4stg_rnd_frac_pre2_in[9]) );
  GTECH_OR2 C8629 ( .A(N5173), .B(N5175), .Z(N5176) );
  GTECH_OR2 C8630 ( .A(N5170), .B(N5172), .Z(N5173) );
  GTECH_OR2 C8631 ( .A(N5167), .B(N5169), .Z(N5170) );
  GTECH_AND2 C8632 ( .A(N5166), .B(a3stg_fracadd[9]), .Z(N5167) );
  GTECH_AND2 C8633 ( .A(N5165), .B(N4406), .Z(N5166) );
  GTECH_AND2 C8634 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5165) );
  GTECH_AND2 C8636 ( .A(N5168), .B(a3stg_fracadd[9]), .Z(N5169) );
  GTECH_AND2 C8637 ( .A(N4409), .B(a6stg_step), .Z(N5168) );
  GTECH_AND2 C8639 ( .A(N5171), .B(a3stg_fracadd[8]), .Z(N5172) );
  GTECH_AND2 C8640 ( .A(N4413), .B(a6stg_step), .Z(N5171) );
  GTECH_AND2 C8642 ( .A(N5174), .B(a4stg_shl[9]), .Z(N5175) );
  GTECH_AND2 C8643 ( .A(N4417), .B(a6stg_step), .Z(N5174) );
  GTECH_AND2 C8645 ( .A(N5177), .B(a4stg_rnd_frac_9), .Z(N5178) );
  GTECH_NOT I_811 ( .A(a6stg_step), .Z(N5177) );
  GTECH_OR2 C8647 ( .A(N5190), .B(N5192), .Z(a4stg_rnd_frac_pre2_in[8]) );
  GTECH_OR2 C8648 ( .A(N5187), .B(N5189), .Z(N5190) );
  GTECH_OR2 C8649 ( .A(N5184), .B(N5186), .Z(N5187) );
  GTECH_OR2 C8650 ( .A(N5181), .B(N5183), .Z(N5184) );
  GTECH_AND2 C8651 ( .A(N5180), .B(a3stg_fracadd[8]), .Z(N5181) );
  GTECH_AND2 C8652 ( .A(N5179), .B(N4406), .Z(N5180) );
  GTECH_AND2 C8653 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5179) );
  GTECH_AND2 C8655 ( .A(N5182), .B(a3stg_fracadd[8]), .Z(N5183) );
  GTECH_AND2 C8656 ( .A(N4409), .B(a6stg_step), .Z(N5182) );
  GTECH_AND2 C8658 ( .A(N5185), .B(a3stg_fracadd[7]), .Z(N5186) );
  GTECH_AND2 C8659 ( .A(N4413), .B(a6stg_step), .Z(N5185) );
  GTECH_AND2 C8661 ( .A(N5188), .B(a4stg_shl[8]), .Z(N5189) );
  GTECH_AND2 C8662 ( .A(N4417), .B(a6stg_step), .Z(N5188) );
  GTECH_AND2 C8664 ( .A(N5191), .B(a4stg_rnd_frac_8), .Z(N5192) );
  GTECH_NOT I_812 ( .A(a6stg_step), .Z(N5191) );
  GTECH_OR2 C8666 ( .A(N5204), .B(N5206), .Z(a4stg_rnd_frac_pre2_in[7]) );
  GTECH_OR2 C8667 ( .A(N5201), .B(N5203), .Z(N5204) );
  GTECH_OR2 C8668 ( .A(N5198), .B(N5200), .Z(N5201) );
  GTECH_OR2 C8669 ( .A(N5195), .B(N5197), .Z(N5198) );
  GTECH_AND2 C8670 ( .A(N5194), .B(a3stg_fracadd[7]), .Z(N5195) );
  GTECH_AND2 C8671 ( .A(N5193), .B(N4406), .Z(N5194) );
  GTECH_AND2 C8672 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5193) );
  GTECH_AND2 C8674 ( .A(N5196), .B(a3stg_fracadd[7]), .Z(N5197) );
  GTECH_AND2 C8675 ( .A(N4409), .B(a6stg_step), .Z(N5196) );
  GTECH_AND2 C8677 ( .A(N5199), .B(a3stg_fracadd[6]), .Z(N5200) );
  GTECH_AND2 C8678 ( .A(N4413), .B(a6stg_step), .Z(N5199) );
  GTECH_AND2 C8680 ( .A(N5202), .B(a4stg_shl[7]), .Z(N5203) );
  GTECH_AND2 C8681 ( .A(N4417), .B(a6stg_step), .Z(N5202) );
  GTECH_AND2 C8683 ( .A(N5205), .B(a4stg_rnd_frac_7), .Z(N5206) );
  GTECH_NOT I_813 ( .A(a6stg_step), .Z(N5205) );
  GTECH_OR2 C8685 ( .A(N5218), .B(N5220), .Z(a4stg_rnd_frac_pre2_in[6]) );
  GTECH_OR2 C8686 ( .A(N5215), .B(N5217), .Z(N5218) );
  GTECH_OR2 C8687 ( .A(N5212), .B(N5214), .Z(N5215) );
  GTECH_OR2 C8688 ( .A(N5209), .B(N5211), .Z(N5212) );
  GTECH_AND2 C8689 ( .A(N5208), .B(a3stg_fracadd[6]), .Z(N5209) );
  GTECH_AND2 C8690 ( .A(N5207), .B(N4406), .Z(N5208) );
  GTECH_AND2 C8691 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5207) );
  GTECH_AND2 C8693 ( .A(N5210), .B(a3stg_fracadd[6]), .Z(N5211) );
  GTECH_AND2 C8694 ( .A(N4409), .B(a6stg_step), .Z(N5210) );
  GTECH_AND2 C8696 ( .A(N5213), .B(a3stg_fracadd[5]), .Z(N5214) );
  GTECH_AND2 C8697 ( .A(N4413), .B(a6stg_step), .Z(N5213) );
  GTECH_AND2 C8699 ( .A(N5216), .B(a4stg_shl[6]), .Z(N5217) );
  GTECH_AND2 C8700 ( .A(N4417), .B(a6stg_step), .Z(N5216) );
  GTECH_AND2 C8702 ( .A(N5219), .B(a4stg_rnd_frac_6), .Z(N5220) );
  GTECH_NOT I_814 ( .A(a6stg_step), .Z(N5219) );
  GTECH_OR2 C8704 ( .A(N5232), .B(N5234), .Z(a4stg_rnd_frac_pre2_in[5]) );
  GTECH_OR2 C8705 ( .A(N5229), .B(N5231), .Z(N5232) );
  GTECH_OR2 C8706 ( .A(N5226), .B(N5228), .Z(N5229) );
  GTECH_OR2 C8707 ( .A(N5223), .B(N5225), .Z(N5226) );
  GTECH_AND2 C8708 ( .A(N5222), .B(a3stg_fracadd[5]), .Z(N5223) );
  GTECH_AND2 C8709 ( .A(N5221), .B(N4406), .Z(N5222) );
  GTECH_AND2 C8710 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5221) );
  GTECH_AND2 C8712 ( .A(N5224), .B(a3stg_fracadd[5]), .Z(N5225) );
  GTECH_AND2 C8713 ( .A(N4409), .B(a6stg_step), .Z(N5224) );
  GTECH_AND2 C8715 ( .A(N5227), .B(a3stg_fracadd[4]), .Z(N5228) );
  GTECH_AND2 C8716 ( .A(N4413), .B(a6stg_step), .Z(N5227) );
  GTECH_AND2 C8718 ( .A(N5230), .B(a4stg_shl[5]), .Z(N5231) );
  GTECH_AND2 C8719 ( .A(N4417), .B(a6stg_step), .Z(N5230) );
  GTECH_AND2 C8721 ( .A(N5233), .B(a4stg_rnd_frac_5), .Z(N5234) );
  GTECH_NOT I_815 ( .A(a6stg_step), .Z(N5233) );
  GTECH_OR2 C8723 ( .A(N5246), .B(N5248), .Z(a4stg_rnd_frac_pre2_in[4]) );
  GTECH_OR2 C8724 ( .A(N5243), .B(N5245), .Z(N5246) );
  GTECH_OR2 C8725 ( .A(N5240), .B(N5242), .Z(N5243) );
  GTECH_OR2 C8726 ( .A(N5237), .B(N5239), .Z(N5240) );
  GTECH_AND2 C8727 ( .A(N5236), .B(a3stg_fracadd[4]), .Z(N5237) );
  GTECH_AND2 C8728 ( .A(N5235), .B(N4406), .Z(N5236) );
  GTECH_AND2 C8729 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5235) );
  GTECH_AND2 C8731 ( .A(N5238), .B(a3stg_fracadd[4]), .Z(N5239) );
  GTECH_AND2 C8732 ( .A(N4409), .B(a6stg_step), .Z(N5238) );
  GTECH_AND2 C8734 ( .A(N5241), .B(a3stg_fracadd[3]), .Z(N5242) );
  GTECH_AND2 C8735 ( .A(N4413), .B(a6stg_step), .Z(N5241) );
  GTECH_AND2 C8737 ( .A(N5244), .B(a4stg_shl[4]), .Z(N5245) );
  GTECH_AND2 C8738 ( .A(N4417), .B(a6stg_step), .Z(N5244) );
  GTECH_AND2 C8740 ( .A(N5247), .B(a4stg_rnd_frac_4), .Z(N5248) );
  GTECH_NOT I_816 ( .A(a6stg_step), .Z(N5247) );
  GTECH_OR2 C8742 ( .A(N5260), .B(N5262), .Z(a4stg_rnd_frac_pre2_in[3]) );
  GTECH_OR2 C8743 ( .A(N5257), .B(N5259), .Z(N5260) );
  GTECH_OR2 C8744 ( .A(N5254), .B(N5256), .Z(N5257) );
  GTECH_OR2 C8745 ( .A(N5251), .B(N5253), .Z(N5254) );
  GTECH_AND2 C8746 ( .A(N5250), .B(a3stg_fracadd[3]), .Z(N5251) );
  GTECH_AND2 C8747 ( .A(N5249), .B(N4406), .Z(N5250) );
  GTECH_AND2 C8748 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5249) );
  GTECH_AND2 C8750 ( .A(N5252), .B(a3stg_fracadd[3]), .Z(N5253) );
  GTECH_AND2 C8751 ( .A(N4409), .B(a6stg_step), .Z(N5252) );
  GTECH_AND2 C8753 ( .A(N5255), .B(a3stg_fracadd[2]), .Z(N5256) );
  GTECH_AND2 C8754 ( .A(N4413), .B(a6stg_step), .Z(N5255) );
  GTECH_AND2 C8756 ( .A(N5258), .B(a4stg_shl[3]), .Z(N5259) );
  GTECH_AND2 C8757 ( .A(N4417), .B(a6stg_step), .Z(N5258) );
  GTECH_AND2 C8759 ( .A(N5261), .B(a4stg_rnd_frac_3), .Z(N5262) );
  GTECH_NOT I_817 ( .A(a6stg_step), .Z(N5261) );
  GTECH_OR2 C8761 ( .A(N5274), .B(N5276), .Z(a4stg_rnd_frac_pre2_in[2]) );
  GTECH_OR2 C8762 ( .A(N5271), .B(N5273), .Z(N5274) );
  GTECH_OR2 C8763 ( .A(N5268), .B(N5270), .Z(N5271) );
  GTECH_OR2 C8764 ( .A(N5265), .B(N5267), .Z(N5268) );
  GTECH_AND2 C8765 ( .A(N5264), .B(a3stg_fracadd[2]), .Z(N5265) );
  GTECH_AND2 C8766 ( .A(N5263), .B(N4406), .Z(N5264) );
  GTECH_AND2 C8767 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5263) );
  GTECH_AND2 C8769 ( .A(N5266), .B(a3stg_fracadd[2]), .Z(N5267) );
  GTECH_AND2 C8770 ( .A(N4409), .B(a6stg_step), .Z(N5266) );
  GTECH_AND2 C8772 ( .A(N5269), .B(a3stg_fracadd[1]), .Z(N5270) );
  GTECH_AND2 C8773 ( .A(N4413), .B(a6stg_step), .Z(N5269) );
  GTECH_AND2 C8775 ( .A(N5272), .B(a4stg_shl[2]), .Z(N5273) );
  GTECH_AND2 C8776 ( .A(N4417), .B(a6stg_step), .Z(N5272) );
  GTECH_AND2 C8778 ( .A(N5275), .B(a4stg_rnd_frac_2), .Z(N5276) );
  GTECH_NOT I_818 ( .A(a6stg_step), .Z(N5275) );
  GTECH_OR2 C8780 ( .A(N5288), .B(N5290), .Z(a4stg_rnd_frac_pre2_in[1]) );
  GTECH_OR2 C8781 ( .A(N5285), .B(N5287), .Z(N5288) );
  GTECH_OR2 C8782 ( .A(N5282), .B(N5284), .Z(N5285) );
  GTECH_OR2 C8783 ( .A(N5279), .B(N5281), .Z(N5282) );
  GTECH_AND2 C8784 ( .A(N5278), .B(a3stg_fracadd[1]), .Z(N5279) );
  GTECH_AND2 C8785 ( .A(N5277), .B(N4406), .Z(N5278) );
  GTECH_AND2 C8786 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5277) );
  GTECH_AND2 C8788 ( .A(N5280), .B(a3stg_fracadd[1]), .Z(N5281) );
  GTECH_AND2 C8789 ( .A(N4409), .B(a6stg_step), .Z(N5280) );
  GTECH_AND2 C8791 ( .A(N5283), .B(a3stg_fracadd[0]), .Z(N5284) );
  GTECH_AND2 C8792 ( .A(N4413), .B(a6stg_step), .Z(N5283) );
  GTECH_AND2 C8794 ( .A(N5286), .B(a4stg_shl[1]), .Z(N5287) );
  GTECH_AND2 C8795 ( .A(N4417), .B(a6stg_step), .Z(N5286) );
  GTECH_AND2 C8797 ( .A(N5289), .B(a4stg_rnd_frac_1), .Z(N5290) );
  GTECH_NOT I_819 ( .A(a6stg_step), .Z(N5289) );
  GTECH_OR2 C8799 ( .A(N5299), .B(N5301), .Z(a4stg_rnd_frac_pre2_in[0]) );
  GTECH_OR2 C8800 ( .A(N5296), .B(N5298), .Z(N5299) );
  GTECH_OR2 C8801 ( .A(N5293), .B(N5295), .Z(N5296) );
  GTECH_AND2 C8802 ( .A(N5292), .B(a3stg_fracadd[0]), .Z(N5293) );
  GTECH_AND2 C8803 ( .A(N5291), .B(N4406), .Z(N5292) );
  GTECH_AND2 C8804 ( .A(a3stg_faddsubopa[1]), .B(a6stg_step), .Z(N5291) );
  GTECH_AND2 C8806 ( .A(N5294), .B(a3stg_fracadd[0]), .Z(N5295) );
  GTECH_AND2 C8807 ( .A(N4409), .B(a6stg_step), .Z(N5294) );
  GTECH_AND2 C8809 ( .A(N5297), .B(a4stg_shl[0]), .Z(N5298) );
  GTECH_AND2 C8810 ( .A(N4417), .B(a6stg_step), .Z(N5297) );
  GTECH_AND2 C8812 ( .A(N5300), .B(a4stg_rnd_frac_0), .Z(N5301) );
  GTECH_NOT I_820 ( .A(a6stg_step), .Z(N5300) );
  GTECH_AND2 C8814 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[63]), .Z(
        a4stg_shl_data_in[63]) );
  GTECH_OR2 C8815 ( .A(N5302), .B(N5303), .Z(a4stg_shl_data_in[62]) );
  GTECH_AND2 C8816 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[62]), .Z(N5302)
         );
  GTECH_AND2 C8817 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[63]), .Z(N5303) );
  GTECH_OR2 C8818 ( .A(N5304), .B(N5305), .Z(a4stg_shl_data_in[61]) );
  GTECH_AND2 C8819 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[61]), .Z(N5304)
         );
  GTECH_AND2 C8820 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[62]), .Z(N5305) );
  GTECH_OR2 C8821 ( .A(N5306), .B(N5307), .Z(a4stg_shl_data_in[60]) );
  GTECH_AND2 C8822 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[60]), .Z(N5306)
         );
  GTECH_AND2 C8823 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[61]), .Z(N5307) );
  GTECH_OR2 C8824 ( .A(N5308), .B(N5309), .Z(a4stg_shl_data_in[59]) );
  GTECH_AND2 C8825 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[59]), .Z(N5308)
         );
  GTECH_AND2 C8826 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[60]), .Z(N5309) );
  GTECH_OR2 C8827 ( .A(N5310), .B(N5311), .Z(a4stg_shl_data_in[58]) );
  GTECH_AND2 C8828 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[58]), .Z(N5310)
         );
  GTECH_AND2 C8829 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[59]), .Z(N5311) );
  GTECH_OR2 C8830 ( .A(N5312), .B(N5313), .Z(a4stg_shl_data_in[57]) );
  GTECH_AND2 C8831 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[57]), .Z(N5312)
         );
  GTECH_AND2 C8832 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[58]), .Z(N5313) );
  GTECH_OR2 C8833 ( .A(N5314), .B(N5315), .Z(a4stg_shl_data_in[56]) );
  GTECH_AND2 C8834 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[56]), .Z(N5314)
         );
  GTECH_AND2 C8835 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[57]), .Z(N5315) );
  GTECH_OR2 C8836 ( .A(N5316), .B(N5317), .Z(a4stg_shl_data_in[55]) );
  GTECH_AND2 C8837 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[55]), .Z(N5316)
         );
  GTECH_AND2 C8838 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[56]), .Z(N5317) );
  GTECH_OR2 C8839 ( .A(N5318), .B(N5319), .Z(a4stg_shl_data_in[54]) );
  GTECH_AND2 C8840 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[54]), .Z(N5318)
         );
  GTECH_AND2 C8841 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[55]), .Z(N5319) );
  GTECH_OR2 C8842 ( .A(N5320), .B(N5321), .Z(a4stg_shl_data_in[53]) );
  GTECH_AND2 C8843 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[53]), .Z(N5320)
         );
  GTECH_AND2 C8844 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[54]), .Z(N5321) );
  GTECH_OR2 C8845 ( .A(N5322), .B(N5323), .Z(a4stg_shl_data_in[52]) );
  GTECH_AND2 C8846 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[52]), .Z(N5322)
         );
  GTECH_AND2 C8847 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[53]), .Z(N5323) );
  GTECH_OR2 C8848 ( .A(N5324), .B(N5325), .Z(a4stg_shl_data_in[51]) );
  GTECH_AND2 C8849 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[51]), .Z(N5324)
         );
  GTECH_AND2 C8850 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[52]), .Z(N5325) );
  GTECH_OR2 C8851 ( .A(N5326), .B(N5327), .Z(a4stg_shl_data_in[50]) );
  GTECH_AND2 C8852 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[50]), .Z(N5326)
         );
  GTECH_AND2 C8853 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[51]), .Z(N5327) );
  GTECH_OR2 C8854 ( .A(N5328), .B(N5329), .Z(a4stg_shl_data_in[49]) );
  GTECH_AND2 C8855 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[49]), .Z(N5328)
         );
  GTECH_AND2 C8856 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[50]), .Z(N5329) );
  GTECH_OR2 C8857 ( .A(N5330), .B(N5331), .Z(a4stg_shl_data_in[48]) );
  GTECH_AND2 C8858 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[48]), .Z(N5330)
         );
  GTECH_AND2 C8859 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[49]), .Z(N5331) );
  GTECH_OR2 C8860 ( .A(N5332), .B(N5333), .Z(a4stg_shl_data_in[47]) );
  GTECH_AND2 C8861 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[47]), .Z(N5332)
         );
  GTECH_AND2 C8862 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[48]), .Z(N5333) );
  GTECH_OR2 C8863 ( .A(N5334), .B(N5335), .Z(a4stg_shl_data_in[46]) );
  GTECH_AND2 C8864 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[46]), .Z(N5334)
         );
  GTECH_AND2 C8865 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[47]), .Z(N5335) );
  GTECH_OR2 C8866 ( .A(N5336), .B(N5337), .Z(a4stg_shl_data_in[45]) );
  GTECH_AND2 C8867 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[45]), .Z(N5336)
         );
  GTECH_AND2 C8868 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[46]), .Z(N5337) );
  GTECH_OR2 C8869 ( .A(N5338), .B(N5339), .Z(a4stg_shl_data_in[44]) );
  GTECH_AND2 C8870 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[44]), .Z(N5338)
         );
  GTECH_AND2 C8871 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[45]), .Z(N5339) );
  GTECH_OR2 C8872 ( .A(N5340), .B(N5341), .Z(a4stg_shl_data_in[43]) );
  GTECH_AND2 C8873 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[43]), .Z(N5340)
         );
  GTECH_AND2 C8874 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[44]), .Z(N5341) );
  GTECH_OR2 C8875 ( .A(N5342), .B(N5343), .Z(a4stg_shl_data_in[42]) );
  GTECH_AND2 C8876 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[42]), .Z(N5342)
         );
  GTECH_AND2 C8877 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[43]), .Z(N5343) );
  GTECH_OR2 C8878 ( .A(N5344), .B(N5345), .Z(a4stg_shl_data_in[41]) );
  GTECH_AND2 C8879 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[41]), .Z(N5344)
         );
  GTECH_AND2 C8880 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[42]), .Z(N5345) );
  GTECH_OR2 C8881 ( .A(N5346), .B(N5347), .Z(a4stg_shl_data_in[40]) );
  GTECH_AND2 C8882 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[40]), .Z(N5346)
         );
  GTECH_AND2 C8883 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[41]), .Z(N5347) );
  GTECH_OR2 C8884 ( .A(N5348), .B(N5349), .Z(a4stg_shl_data_in[39]) );
  GTECH_AND2 C8885 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[39]), .Z(N5348)
         );
  GTECH_AND2 C8886 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[40]), .Z(N5349) );
  GTECH_OR2 C8887 ( .A(N5350), .B(N5351), .Z(a4stg_shl_data_in[38]) );
  GTECH_AND2 C8888 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[38]), .Z(N5350)
         );
  GTECH_AND2 C8889 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[39]), .Z(N5351) );
  GTECH_OR2 C8890 ( .A(N5352), .B(N5353), .Z(a4stg_shl_data_in[37]) );
  GTECH_AND2 C8891 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[37]), .Z(N5352)
         );
  GTECH_AND2 C8892 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[38]), .Z(N5353) );
  GTECH_OR2 C8893 ( .A(N5354), .B(N5355), .Z(a4stg_shl_data_in[36]) );
  GTECH_AND2 C8894 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[36]), .Z(N5354)
         );
  GTECH_AND2 C8895 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[37]), .Z(N5355) );
  GTECH_OR2 C8896 ( .A(N5356), .B(N5357), .Z(a4stg_shl_data_in[35]) );
  GTECH_AND2 C8897 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[35]), .Z(N5356)
         );
  GTECH_AND2 C8898 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[36]), .Z(N5357) );
  GTECH_OR2 C8899 ( .A(N5358), .B(N5359), .Z(a4stg_shl_data_in[34]) );
  GTECH_AND2 C8900 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[34]), .Z(N5358)
         );
  GTECH_AND2 C8901 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[35]), .Z(N5359) );
  GTECH_OR2 C8902 ( .A(N5360), .B(N5361), .Z(a4stg_shl_data_in[33]) );
  GTECH_AND2 C8903 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[33]), .Z(N5360)
         );
  GTECH_AND2 C8904 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[34]), .Z(N5361) );
  GTECH_OR2 C8905 ( .A(N5362), .B(N5363), .Z(a4stg_shl_data_in[32]) );
  GTECH_AND2 C8906 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[32]), .Z(N5362)
         );
  GTECH_AND2 C8907 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[33]), .Z(N5363) );
  GTECH_OR2 C8908 ( .A(N5364), .B(N5365), .Z(a4stg_shl_data_in[31]) );
  GTECH_AND2 C8909 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[31]), .Z(N5364)
         );
  GTECH_AND2 C8910 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[32]), .Z(N5365) );
  GTECH_OR2 C8911 ( .A(N5366), .B(N5367), .Z(a4stg_shl_data_in[30]) );
  GTECH_AND2 C8912 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[30]), .Z(N5366)
         );
  GTECH_AND2 C8913 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[31]), .Z(N5367) );
  GTECH_OR2 C8914 ( .A(N5368), .B(N5369), .Z(a4stg_shl_data_in[29]) );
  GTECH_AND2 C8915 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[29]), .Z(N5368)
         );
  GTECH_AND2 C8916 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[30]), .Z(N5369) );
  GTECH_OR2 C8917 ( .A(N5370), .B(N5371), .Z(a4stg_shl_data_in[28]) );
  GTECH_AND2 C8918 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[28]), .Z(N5370)
         );
  GTECH_AND2 C8919 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[29]), .Z(N5371) );
  GTECH_OR2 C8920 ( .A(N5372), .B(N5373), .Z(a4stg_shl_data_in[27]) );
  GTECH_AND2 C8921 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[27]), .Z(N5372)
         );
  GTECH_AND2 C8922 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[28]), .Z(N5373) );
  GTECH_OR2 C8923 ( .A(N5374), .B(N5375), .Z(a4stg_shl_data_in[26]) );
  GTECH_AND2 C8924 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[26]), .Z(N5374)
         );
  GTECH_AND2 C8925 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[27]), .Z(N5375) );
  GTECH_OR2 C8926 ( .A(N5376), .B(N5377), .Z(a4stg_shl_data_in[25]) );
  GTECH_AND2 C8927 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[25]), .Z(N5376)
         );
  GTECH_AND2 C8928 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[26]), .Z(N5377) );
  GTECH_OR2 C8929 ( .A(N5378), .B(N5379), .Z(a4stg_shl_data_in[24]) );
  GTECH_AND2 C8930 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[24]), .Z(N5378)
         );
  GTECH_AND2 C8931 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[25]), .Z(N5379) );
  GTECH_OR2 C8932 ( .A(N5380), .B(N5381), .Z(a4stg_shl_data_in[23]) );
  GTECH_AND2 C8933 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[23]), .Z(N5380)
         );
  GTECH_AND2 C8934 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[24]), .Z(N5381) );
  GTECH_OR2 C8935 ( .A(N5382), .B(N5383), .Z(a4stg_shl_data_in[22]) );
  GTECH_AND2 C8936 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[22]), .Z(N5382)
         );
  GTECH_AND2 C8937 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[23]), .Z(N5383) );
  GTECH_OR2 C8938 ( .A(N5384), .B(N5385), .Z(a4stg_shl_data_in[21]) );
  GTECH_AND2 C8939 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[21]), .Z(N5384)
         );
  GTECH_AND2 C8940 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[22]), .Z(N5385) );
  GTECH_OR2 C8941 ( .A(N5386), .B(N5387), .Z(a4stg_shl_data_in[20]) );
  GTECH_AND2 C8942 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[20]), .Z(N5386)
         );
  GTECH_AND2 C8943 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[21]), .Z(N5387) );
  GTECH_OR2 C8944 ( .A(N5388), .B(N5389), .Z(a4stg_shl_data_in[19]) );
  GTECH_AND2 C8945 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[19]), .Z(N5388)
         );
  GTECH_AND2 C8946 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[20]), .Z(N5389) );
  GTECH_OR2 C8947 ( .A(N5390), .B(N5391), .Z(a4stg_shl_data_in[18]) );
  GTECH_AND2 C8948 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[18]), .Z(N5390)
         );
  GTECH_AND2 C8949 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[19]), .Z(N5391) );
  GTECH_OR2 C8950 ( .A(N5392), .B(N5393), .Z(a4stg_shl_data_in[17]) );
  GTECH_AND2 C8951 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[17]), .Z(N5392)
         );
  GTECH_AND2 C8952 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[18]), .Z(N5393) );
  GTECH_OR2 C8953 ( .A(N5394), .B(N5395), .Z(a4stg_shl_data_in[16]) );
  GTECH_AND2 C8954 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[16]), .Z(N5394)
         );
  GTECH_AND2 C8955 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[17]), .Z(N5395) );
  GTECH_OR2 C8956 ( .A(N5396), .B(N5397), .Z(a4stg_shl_data_in[15]) );
  GTECH_AND2 C8957 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[15]), .Z(N5396)
         );
  GTECH_AND2 C8958 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[16]), .Z(N5397) );
  GTECH_OR2 C8959 ( .A(N5398), .B(N5399), .Z(a4stg_shl_data_in[14]) );
  GTECH_AND2 C8960 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[14]), .Z(N5398)
         );
  GTECH_AND2 C8961 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[15]), .Z(N5399) );
  GTECH_OR2 C8962 ( .A(N5400), .B(N5401), .Z(a4stg_shl_data_in[13]) );
  GTECH_AND2 C8963 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[13]), .Z(N5400)
         );
  GTECH_AND2 C8964 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[14]), .Z(N5401) );
  GTECH_OR2 C8965 ( .A(N5402), .B(N5403), .Z(a4stg_shl_data_in[12]) );
  GTECH_AND2 C8966 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[12]), .Z(N5402)
         );
  GTECH_AND2 C8967 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[13]), .Z(N5403) );
  GTECH_OR2 C8968 ( .A(N5404), .B(N5405), .Z(a4stg_shl_data_in[11]) );
  GTECH_AND2 C8969 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[11]), .Z(N5404)
         );
  GTECH_AND2 C8970 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[12]), .Z(N5405) );
  GTECH_OR2 C8971 ( .A(N5406), .B(N5407), .Z(a4stg_shl_data_in[10]) );
  GTECH_AND2 C8972 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[10]), .Z(N5406)
         );
  GTECH_AND2 C8973 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[11]), .Z(N5407) );
  GTECH_OR2 C8974 ( .A(N5408), .B(N5409), .Z(a4stg_shl_data_in[9]) );
  GTECH_AND2 C8975 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[9]), .Z(N5408)
         );
  GTECH_AND2 C8976 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[10]), .Z(N5409) );
  GTECH_OR2 C8977 ( .A(N5410), .B(N5411), .Z(a4stg_shl_data_in[8]) );
  GTECH_AND2 C8978 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[8]), .Z(N5410)
         );
  GTECH_AND2 C8979 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[9]), .Z(N5411) );
  GTECH_OR2 C8980 ( .A(N5412), .B(N5413), .Z(a4stg_shl_data_in[7]) );
  GTECH_AND2 C8981 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[7]), .Z(N5412)
         );
  GTECH_AND2 C8982 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[8]), .Z(N5413) );
  GTECH_OR2 C8983 ( .A(N5414), .B(N5415), .Z(a4stg_shl_data_in[6]) );
  GTECH_AND2 C8984 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[6]), .Z(N5414)
         );
  GTECH_AND2 C8985 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[7]), .Z(N5415) );
  GTECH_OR2 C8986 ( .A(N5416), .B(N5417), .Z(a4stg_shl_data_in[5]) );
  GTECH_AND2 C8987 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[5]), .Z(N5416)
         );
  GTECH_AND2 C8988 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[6]), .Z(N5417) );
  GTECH_OR2 C8989 ( .A(N5418), .B(N5419), .Z(a4stg_shl_data_in[4]) );
  GTECH_AND2 C8990 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[4]), .Z(N5418)
         );
  GTECH_AND2 C8991 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[5]), .Z(N5419) );
  GTECH_OR2 C8992 ( .A(N5420), .B(N5421), .Z(a4stg_shl_data_in[3]) );
  GTECH_AND2 C8993 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[3]), .Z(N5420)
         );
  GTECH_AND2 C8994 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[4]), .Z(N5421) );
  GTECH_OR2 C8995 ( .A(N5422), .B(N5423), .Z(a4stg_shl_data_in[2]) );
  GTECH_AND2 C8996 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[2]), .Z(N5422)
         );
  GTECH_AND2 C8997 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[3]), .Z(N5423) );
  GTECH_OR2 C8998 ( .A(N5424), .B(N5425), .Z(a4stg_shl_data_in[1]) );
  GTECH_AND2 C8999 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[1]), .Z(N5424)
         );
  GTECH_AND2 C9000 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[2]), .Z(N5425) );
  GTECH_OR2 C9001 ( .A(N5426), .B(N5427), .Z(a4stg_shl_data_in[0]) );
  GTECH_AND2 C9002 ( .A(a3stg_denorm_inva), .B(a3stg_ld0_frac[0]), .Z(N5426)
         );
  GTECH_AND2 C9003 ( .A(a3stg_denorma), .B(a3stg_ld0_frac[1]), .Z(N5427) );
  GTECH_OR2 C9004 ( .A(N5428), .B(a4stg_rnd_frac_pre3[63]), .Z(
        a4stg_rnd_frac_63) );
  GTECH_OR2 C9005 ( .A(a4stg_rnd_frac_pre1[63]), .B(a4stg_rnd_frac_pre2[63]), 
        .Z(N5428) );
  GTECH_OR2 C9006 ( .A(N5429), .B(a4stg_rnd_frac_pre3[62]), .Z(
        a4stg_rnd_frac_62) );
  GTECH_OR2 C9007 ( .A(a4stg_rnd_frac_pre1[62]), .B(a4stg_rnd_frac_pre2[62]), 
        .Z(N5429) );
  GTECH_OR2 C9008 ( .A(N5430), .B(a4stg_rnd_frac_pre3[61]), .Z(
        a4stg_rnd_frac_61) );
  GTECH_OR2 C9009 ( .A(a4stg_rnd_frac_pre1[61]), .B(a4stg_rnd_frac_pre2[61]), 
        .Z(N5430) );
  GTECH_OR2 C9010 ( .A(N5431), .B(a4stg_rnd_frac_pre3[60]), .Z(
        a4stg_rnd_frac_60) );
  GTECH_OR2 C9011 ( .A(a4stg_rnd_frac_pre1[60]), .B(a4stg_rnd_frac_pre2[60]), 
        .Z(N5431) );
  GTECH_OR2 C9012 ( .A(N5432), .B(a4stg_rnd_frac_pre3[59]), .Z(
        a4stg_rnd_frac_59) );
  GTECH_OR2 C9013 ( .A(a4stg_rnd_frac_pre1[59]), .B(a4stg_rnd_frac_pre2[59]), 
        .Z(N5432) );
  GTECH_OR2 C9014 ( .A(N5433), .B(a4stg_rnd_frac_pre3[58]), .Z(
        a4stg_rnd_frac_58) );
  GTECH_OR2 C9015 ( .A(a4stg_rnd_frac_pre1[58]), .B(a4stg_rnd_frac_pre2[58]), 
        .Z(N5433) );
  GTECH_OR2 C9016 ( .A(N5434), .B(a4stg_rnd_frac_pre3[57]), .Z(
        a4stg_rnd_frac_57) );
  GTECH_OR2 C9017 ( .A(a4stg_rnd_frac_pre1[57]), .B(a4stg_rnd_frac_pre2[57]), 
        .Z(N5434) );
  GTECH_OR2 C9018 ( .A(N5435), .B(a4stg_rnd_frac_pre3[56]), .Z(
        a4stg_rnd_frac_56) );
  GTECH_OR2 C9019 ( .A(a4stg_rnd_frac_pre1[56]), .B(a4stg_rnd_frac_pre2[56]), 
        .Z(N5435) );
  GTECH_OR2 C9020 ( .A(N5436), .B(a4stg_rnd_frac_pre3[55]), .Z(
        a4stg_rnd_frac_55) );
  GTECH_OR2 C9021 ( .A(a4stg_rnd_frac_pre1[55]), .B(a4stg_rnd_frac_pre2[55]), 
        .Z(N5436) );
  GTECH_OR2 C9022 ( .A(N5437), .B(a4stg_rnd_frac_pre3[54]), .Z(
        a4stg_rnd_frac_54) );
  GTECH_OR2 C9023 ( .A(a4stg_rnd_frac_pre1[54]), .B(a4stg_rnd_frac_pre2[54]), 
        .Z(N5437) );
  GTECH_OR2 C9024 ( .A(N5438), .B(a4stg_rnd_frac_pre3[53]), .Z(
        a4stg_rnd_frac_53) );
  GTECH_OR2 C9025 ( .A(a4stg_rnd_frac_pre1[53]), .B(a4stg_rnd_frac_pre2[53]), 
        .Z(N5438) );
  GTECH_OR2 C9026 ( .A(N5439), .B(a4stg_rnd_frac_pre3[52]), .Z(
        a4stg_rnd_frac_52) );
  GTECH_OR2 C9027 ( .A(a4stg_rnd_frac_pre1[52]), .B(a4stg_rnd_frac_pre2[52]), 
        .Z(N5439) );
  GTECH_OR2 C9028 ( .A(N5440), .B(a4stg_rnd_frac_pre3[51]), .Z(
        a4stg_rnd_frac_51) );
  GTECH_OR2 C9029 ( .A(a4stg_rnd_frac_pre1[51]), .B(a4stg_rnd_frac_pre2[51]), 
        .Z(N5440) );
  GTECH_OR2 C9030 ( .A(N5441), .B(a4stg_rnd_frac_pre3[50]), .Z(
        a4stg_rnd_frac_50) );
  GTECH_OR2 C9031 ( .A(a4stg_rnd_frac_pre1[50]), .B(a4stg_rnd_frac_pre2[50]), 
        .Z(N5441) );
  GTECH_OR2 C9032 ( .A(N5442), .B(a4stg_rnd_frac_pre3[49]), .Z(
        a4stg_rnd_frac_49) );
  GTECH_OR2 C9033 ( .A(a4stg_rnd_frac_pre1[49]), .B(a4stg_rnd_frac_pre2[49]), 
        .Z(N5442) );
  GTECH_OR2 C9034 ( .A(N5443), .B(a4stg_rnd_frac_pre3[48]), .Z(
        a4stg_rnd_frac_48) );
  GTECH_OR2 C9035 ( .A(a4stg_rnd_frac_pre1[48]), .B(a4stg_rnd_frac_pre2[48]), 
        .Z(N5443) );
  GTECH_OR2 C9036 ( .A(N5444), .B(a4stg_rnd_frac_pre3[47]), .Z(
        a4stg_rnd_frac_47) );
  GTECH_OR2 C9037 ( .A(a4stg_rnd_frac_pre1[47]), .B(a4stg_rnd_frac_pre2[47]), 
        .Z(N5444) );
  GTECH_OR2 C9038 ( .A(N5445), .B(a4stg_rnd_frac_pre3[46]), .Z(
        a4stg_rnd_frac_46) );
  GTECH_OR2 C9039 ( .A(a4stg_rnd_frac_pre1[46]), .B(a4stg_rnd_frac_pre2[46]), 
        .Z(N5445) );
  GTECH_OR2 C9040 ( .A(N5446), .B(a4stg_rnd_frac_pre3[45]), .Z(
        a4stg_rnd_frac_45) );
  GTECH_OR2 C9041 ( .A(a4stg_rnd_frac_pre1[45]), .B(a4stg_rnd_frac_pre2[45]), 
        .Z(N5446) );
  GTECH_OR2 C9042 ( .A(N5447), .B(a4stg_rnd_frac_pre3[44]), .Z(
        a4stg_rnd_frac_44) );
  GTECH_OR2 C9043 ( .A(a4stg_rnd_frac_pre1[44]), .B(a4stg_rnd_frac_pre2[44]), 
        .Z(N5447) );
  GTECH_OR2 C9044 ( .A(N5448), .B(a4stg_rnd_frac_pre3[43]), .Z(
        a4stg_rnd_frac_43) );
  GTECH_OR2 C9045 ( .A(a4stg_rnd_frac_pre1[43]), .B(a4stg_rnd_frac_pre2[43]), 
        .Z(N5448) );
  GTECH_OR2 C9046 ( .A(N5449), .B(a4stg_rnd_frac_pre3[42]), .Z(
        a4stg_rnd_frac_42) );
  GTECH_OR2 C9047 ( .A(a4stg_rnd_frac_pre1[42]), .B(a4stg_rnd_frac_pre2[42]), 
        .Z(N5449) );
  GTECH_OR2 C9048 ( .A(N5450), .B(a4stg_rnd_frac_pre3[41]), .Z(
        a4stg_rnd_frac_41) );
  GTECH_OR2 C9049 ( .A(a4stg_rnd_frac_pre1[41]), .B(a4stg_rnd_frac_pre2[41]), 
        .Z(N5450) );
  GTECH_OR2 C9050 ( .A(N5451), .B(a4stg_rnd_frac_pre3[40]), .Z(
        a4stg_rnd_frac_40) );
  GTECH_OR2 C9051 ( .A(a4stg_rnd_frac_pre1[40]), .B(a4stg_rnd_frac_pre2[40]), 
        .Z(N5451) );
  GTECH_OR2 C9052 ( .A(N5452), .B(a4stg_rnd_frac_pre3[39]), .Z(
        a4stg_rnd_frac_39) );
  GTECH_OR2 C9053 ( .A(a4stg_rnd_frac_pre1[39]), .B(a4stg_rnd_frac_pre2[39]), 
        .Z(N5452) );
  GTECH_OR2 C9054 ( .A(N5453), .B(a4stg_rnd_frac_pre3[38]), .Z(
        a4stg_rnd_frac[38]) );
  GTECH_OR2 C9055 ( .A(a4stg_rnd_frac_pre1[38]), .B(a4stg_rnd_frac_pre2[38]), 
        .Z(N5453) );
  GTECH_OR2 C9056 ( .A(N5454), .B(a4stg_rnd_frac_pre3[37]), .Z(
        a4stg_rnd_frac[37]) );
  GTECH_OR2 C9057 ( .A(a4stg_rnd_frac_pre1[37]), .B(a4stg_rnd_frac_pre2[37]), 
        .Z(N5454) );
  GTECH_OR2 C9058 ( .A(N5455), .B(a4stg_rnd_frac_pre3[36]), .Z(
        a4stg_rnd_frac[36]) );
  GTECH_OR2 C9059 ( .A(a4stg_rnd_frac_pre1[36]), .B(a4stg_rnd_frac_pre2[36]), 
        .Z(N5455) );
  GTECH_OR2 C9060 ( .A(N5456), .B(a4stg_rnd_frac_pre3[35]), .Z(
        a4stg_rnd_frac[35]) );
  GTECH_OR2 C9061 ( .A(a4stg_rnd_frac_pre1[35]), .B(a4stg_rnd_frac_pre2[35]), 
        .Z(N5456) );
  GTECH_OR2 C9062 ( .A(N5457), .B(a4stg_rnd_frac_pre3[34]), .Z(
        a4stg_rnd_frac[34]) );
  GTECH_OR2 C9063 ( .A(a4stg_rnd_frac_pre1[34]), .B(a4stg_rnd_frac_pre2[34]), 
        .Z(N5457) );
  GTECH_OR2 C9064 ( .A(N5458), .B(a4stg_rnd_frac_pre3[33]), .Z(
        a4stg_rnd_frac[33]) );
  GTECH_OR2 C9065 ( .A(a4stg_rnd_frac_pre1[33]), .B(a4stg_rnd_frac_pre2[33]), 
        .Z(N5458) );
  GTECH_OR2 C9066 ( .A(N5459), .B(a4stg_rnd_frac_pre3[32]), .Z(
        a4stg_rnd_frac[32]) );
  GTECH_OR2 C9067 ( .A(a4stg_rnd_frac_pre1[32]), .B(a4stg_rnd_frac_pre2[32]), 
        .Z(N5459) );
  GTECH_OR2 C9068 ( .A(N5460), .B(a4stg_rnd_frac_pre3[31]), .Z(
        a4stg_rnd_frac[31]) );
  GTECH_OR2 C9069 ( .A(a4stg_rnd_frac_pre1[31]), .B(a4stg_rnd_frac_pre2[31]), 
        .Z(N5460) );
  GTECH_OR2 C9070 ( .A(N5461), .B(a4stg_rnd_frac_pre3[30]), .Z(
        a4stg_rnd_frac[30]) );
  GTECH_OR2 C9071 ( .A(a4stg_rnd_frac_pre1[30]), .B(a4stg_rnd_frac_pre2[30]), 
        .Z(N5461) );
  GTECH_OR2 C9072 ( .A(N5462), .B(a4stg_rnd_frac_pre3[29]), .Z(
        a4stg_rnd_frac[29]) );
  GTECH_OR2 C9073 ( .A(a4stg_rnd_frac_pre1[29]), .B(a4stg_rnd_frac_pre2[29]), 
        .Z(N5462) );
  GTECH_OR2 C9074 ( .A(N5463), .B(a4stg_rnd_frac_pre3[28]), .Z(
        a4stg_rnd_frac[28]) );
  GTECH_OR2 C9075 ( .A(a4stg_rnd_frac_pre1[28]), .B(a4stg_rnd_frac_pre2[28]), 
        .Z(N5463) );
  GTECH_OR2 C9076 ( .A(N5464), .B(a4stg_rnd_frac_pre3[27]), .Z(
        a4stg_rnd_frac[27]) );
  GTECH_OR2 C9077 ( .A(a4stg_rnd_frac_pre1[27]), .B(a4stg_rnd_frac_pre2[27]), 
        .Z(N5464) );
  GTECH_OR2 C9078 ( .A(N5465), .B(a4stg_rnd_frac_pre3[26]), .Z(
        a4stg_rnd_frac[26]) );
  GTECH_OR2 C9079 ( .A(a4stg_rnd_frac_pre1[26]), .B(a4stg_rnd_frac_pre2[26]), 
        .Z(N5465) );
  GTECH_OR2 C9080 ( .A(N5466), .B(a4stg_rnd_frac_pre3[25]), .Z(
        a4stg_rnd_frac[25]) );
  GTECH_OR2 C9081 ( .A(a4stg_rnd_frac_pre1[25]), .B(a4stg_rnd_frac_pre2[25]), 
        .Z(N5466) );
  GTECH_OR2 C9082 ( .A(N5467), .B(a4stg_rnd_frac_pre3[24]), .Z(
        a4stg_rnd_frac[24]) );
  GTECH_OR2 C9083 ( .A(a4stg_rnd_frac_pre1[24]), .B(a4stg_rnd_frac_pre2[24]), 
        .Z(N5467) );
  GTECH_OR2 C9084 ( .A(N5468), .B(a4stg_rnd_frac_pre3[23]), .Z(
        a4stg_rnd_frac[23]) );
  GTECH_OR2 C9085 ( .A(a4stg_rnd_frac_pre1[23]), .B(a4stg_rnd_frac_pre2[23]), 
        .Z(N5468) );
  GTECH_OR2 C9086 ( .A(N5469), .B(a4stg_rnd_frac_pre3[22]), .Z(
        a4stg_rnd_frac[22]) );
  GTECH_OR2 C9087 ( .A(a4stg_rnd_frac_pre1[22]), .B(a4stg_rnd_frac_pre2[22]), 
        .Z(N5469) );
  GTECH_OR2 C9088 ( .A(N5470), .B(a4stg_rnd_frac_pre3[21]), .Z(
        a4stg_rnd_frac[21]) );
  GTECH_OR2 C9089 ( .A(a4stg_rnd_frac_pre1[21]), .B(a4stg_rnd_frac_pre2[21]), 
        .Z(N5470) );
  GTECH_OR2 C9090 ( .A(N5471), .B(a4stg_rnd_frac_pre3[20]), .Z(
        a4stg_rnd_frac[20]) );
  GTECH_OR2 C9091 ( .A(a4stg_rnd_frac_pre1[20]), .B(a4stg_rnd_frac_pre2[20]), 
        .Z(N5471) );
  GTECH_OR2 C9092 ( .A(N5472), .B(a4stg_rnd_frac_pre3[19]), .Z(
        a4stg_rnd_frac[19]) );
  GTECH_OR2 C9093 ( .A(a4stg_rnd_frac_pre1[19]), .B(a4stg_rnd_frac_pre2[19]), 
        .Z(N5472) );
  GTECH_OR2 C9094 ( .A(N5473), .B(a4stg_rnd_frac_pre3[18]), .Z(
        a4stg_rnd_frac[18]) );
  GTECH_OR2 C9095 ( .A(a4stg_rnd_frac_pre1[18]), .B(a4stg_rnd_frac_pre2[18]), 
        .Z(N5473) );
  GTECH_OR2 C9096 ( .A(N5474), .B(a4stg_rnd_frac_pre3[17]), .Z(
        a4stg_rnd_frac[17]) );
  GTECH_OR2 C9097 ( .A(a4stg_rnd_frac_pre1[17]), .B(a4stg_rnd_frac_pre2[17]), 
        .Z(N5474) );
  GTECH_OR2 C9098 ( .A(N5475), .B(a4stg_rnd_frac_pre3[16]), .Z(
        a4stg_rnd_frac[16]) );
  GTECH_OR2 C9099 ( .A(a4stg_rnd_frac_pre1[16]), .B(a4stg_rnd_frac_pre2[16]), 
        .Z(N5475) );
  GTECH_OR2 C9100 ( .A(N5476), .B(a4stg_rnd_frac_pre3[15]), .Z(
        a4stg_rnd_frac[15]) );
  GTECH_OR2 C9101 ( .A(a4stg_rnd_frac_pre1[15]), .B(a4stg_rnd_frac_pre2[15]), 
        .Z(N5476) );
  GTECH_OR2 C9102 ( .A(N5477), .B(a4stg_rnd_frac_pre3[14]), .Z(
        a4stg_rnd_frac[14]) );
  GTECH_OR2 C9103 ( .A(a4stg_rnd_frac_pre1[14]), .B(a4stg_rnd_frac_pre2[14]), 
        .Z(N5477) );
  GTECH_OR2 C9104 ( .A(N5478), .B(a4stg_rnd_frac_pre3[13]), .Z(
        a4stg_rnd_frac[13]) );
  GTECH_OR2 C9105 ( .A(a4stg_rnd_frac_pre1[13]), .B(a4stg_rnd_frac_pre2[13]), 
        .Z(N5478) );
  GTECH_OR2 C9106 ( .A(N5479), .B(a4stg_rnd_frac_pre3[12]), .Z(
        a4stg_rnd_frac[12]) );
  GTECH_OR2 C9107 ( .A(a4stg_rnd_frac_pre1[12]), .B(a4stg_rnd_frac_pre2[12]), 
        .Z(N5479) );
  GTECH_OR2 C9108 ( .A(N5480), .B(a4stg_rnd_frac_pre3[11]), .Z(
        a4stg_rnd_frac_11) );
  GTECH_OR2 C9109 ( .A(a4stg_rnd_frac_pre1[11]), .B(a4stg_rnd_frac_pre2[11]), 
        .Z(N5480) );
  GTECH_OR2 C9110 ( .A(N5481), .B(a4stg_rnd_frac_pre3[10]), .Z(
        a4stg_rnd_frac_10) );
  GTECH_OR2 C9111 ( .A(a4stg_rnd_frac_pre1[10]), .B(a4stg_rnd_frac_pre2[10]), 
        .Z(N5481) );
  GTECH_OR2 C9112 ( .A(N5482), .B(a4stg_rnd_frac_pre3[9]), .Z(a4stg_rnd_frac_9) );
  GTECH_OR2 C9113 ( .A(a4stg_rnd_frac_pre1[9]), .B(a4stg_rnd_frac_pre2[9]), 
        .Z(N5482) );
  GTECH_OR2 C9114 ( .A(N5483), .B(a4stg_rnd_frac_pre3[8]), .Z(a4stg_rnd_frac_8) );
  GTECH_OR2 C9115 ( .A(a4stg_rnd_frac_pre1[8]), .B(a4stg_rnd_frac_pre2[8]), 
        .Z(N5483) );
  GTECH_OR2 C9116 ( .A(N5484), .B(a4stg_rnd_frac_pre3[7]), .Z(a4stg_rnd_frac_7) );
  GTECH_OR2 C9117 ( .A(a4stg_rnd_frac_pre1[7]), .B(a4stg_rnd_frac_pre2[7]), 
        .Z(N5484) );
  GTECH_OR2 C9118 ( .A(N5485), .B(a4stg_rnd_frac_pre3[6]), .Z(a4stg_rnd_frac_6) );
  GTECH_OR2 C9119 ( .A(a4stg_rnd_frac_pre1[6]), .B(a4stg_rnd_frac_pre2[6]), 
        .Z(N5485) );
  GTECH_OR2 C9120 ( .A(N5486), .B(a4stg_rnd_frac_pre3[5]), .Z(a4stg_rnd_frac_5) );
  GTECH_OR2 C9121 ( .A(a4stg_rnd_frac_pre1[5]), .B(a4stg_rnd_frac_pre2[5]), 
        .Z(N5486) );
  GTECH_OR2 C9122 ( .A(N5487), .B(a4stg_rnd_frac_pre3[4]), .Z(a4stg_rnd_frac_4) );
  GTECH_OR2 C9123 ( .A(a4stg_rnd_frac_pre1[4]), .B(a4stg_rnd_frac_pre2[4]), 
        .Z(N5487) );
  GTECH_OR2 C9124 ( .A(N5488), .B(a4stg_rnd_frac_pre3[3]), .Z(a4stg_rnd_frac_3) );
  GTECH_OR2 C9125 ( .A(a4stg_rnd_frac_pre1[3]), .B(a4stg_rnd_frac_pre2[3]), 
        .Z(N5488) );
  GTECH_OR2 C9126 ( .A(N5489), .B(a4stg_rnd_frac_pre3[2]), .Z(a4stg_rnd_frac_2) );
  GTECH_OR2 C9127 ( .A(a4stg_rnd_frac_pre1[2]), .B(a4stg_rnd_frac_pre2[2]), 
        .Z(N5489) );
  GTECH_OR2 C9128 ( .A(N5490), .B(a4stg_rnd_frac_pre3[1]), .Z(a4stg_rnd_frac_1) );
  GTECH_OR2 C9129 ( .A(a4stg_rnd_frac_pre1[1]), .B(a4stg_rnd_frac_pre2[1]), 
        .Z(N5490) );
  GTECH_OR2 C9130 ( .A(N5491), .B(a4stg_rnd_frac_pre3[0]), .Z(a4stg_rnd_frac_0) );
  GTECH_OR2 C9131 ( .A(a4stg_rnd_frac_pre1[0]), .B(a4stg_rnd_frac_pre2[0]), 
        .Z(N5491) );
  GTECH_OR2 C9132 ( .A(N5499), .B(a4stg_rnd_frac_0), .Z(a4stg_frac_9_0_nx) );
  GTECH_OR2 C9133 ( .A(N5498), .B(a4stg_rnd_frac_1), .Z(N5499) );
  GTECH_OR2 C9134 ( .A(N5497), .B(a4stg_rnd_frac_2), .Z(N5498) );
  GTECH_OR2 C9135 ( .A(N5496), .B(a4stg_rnd_frac_3), .Z(N5497) );
  GTECH_OR2 C9136 ( .A(N5495), .B(a4stg_rnd_frac_4), .Z(N5496) );
  GTECH_OR2 C9137 ( .A(N5494), .B(a4stg_rnd_frac_5), .Z(N5495) );
  GTECH_OR2 C9138 ( .A(N5493), .B(a4stg_rnd_frac_6), .Z(N5494) );
  GTECH_OR2 C9139 ( .A(N5492), .B(a4stg_rnd_frac_7), .Z(N5493) );
  GTECH_OR2 C9140 ( .A(a4stg_rnd_frac_9), .B(a4stg_rnd_frac_8), .Z(N5492) );
  GTECH_OR2 C9141 ( .A(a4stg_frac_9_0_nx), .B(a4stg_rnd_frac_10), .Z(
        a4stg_frac_dbl_nx) );
  GTECH_OR2 C9142 ( .A(a4stg_frac_dbl_nx), .B(N5526), .Z(a4stg_frac_38_0_nx)
         );
  GTECH_OR2 C9143 ( .A(N5525), .B(a4stg_rnd_frac_11), .Z(N5526) );
  GTECH_OR2 C9144 ( .A(N5524), .B(a4stg_rnd_frac[12]), .Z(N5525) );
  GTECH_OR2 C9145 ( .A(N5523), .B(a4stg_rnd_frac[13]), .Z(N5524) );
  GTECH_OR2 C9146 ( .A(N5522), .B(a4stg_rnd_frac[14]), .Z(N5523) );
  GTECH_OR2 C9147 ( .A(N5521), .B(a4stg_rnd_frac[15]), .Z(N5522) );
  GTECH_OR2 C9148 ( .A(N5520), .B(a4stg_rnd_frac[16]), .Z(N5521) );
  GTECH_OR2 C9149 ( .A(N5519), .B(a4stg_rnd_frac[17]), .Z(N5520) );
  GTECH_OR2 C9150 ( .A(N5518), .B(a4stg_rnd_frac[18]), .Z(N5519) );
  GTECH_OR2 C9151 ( .A(N5517), .B(a4stg_rnd_frac[19]), .Z(N5518) );
  GTECH_OR2 C9152 ( .A(N5516), .B(a4stg_rnd_frac[20]), .Z(N5517) );
  GTECH_OR2 C9153 ( .A(N5515), .B(a4stg_rnd_frac[21]), .Z(N5516) );
  GTECH_OR2 C9154 ( .A(N5514), .B(a4stg_rnd_frac[22]), .Z(N5515) );
  GTECH_OR2 C9155 ( .A(N5513), .B(a4stg_rnd_frac[23]), .Z(N5514) );
  GTECH_OR2 C9156 ( .A(N5512), .B(a4stg_rnd_frac[24]), .Z(N5513) );
  GTECH_OR2 C9157 ( .A(N5511), .B(a4stg_rnd_frac[25]), .Z(N5512) );
  GTECH_OR2 C9158 ( .A(N5510), .B(a4stg_rnd_frac[26]), .Z(N5511) );
  GTECH_OR2 C9159 ( .A(N5509), .B(a4stg_rnd_frac[27]), .Z(N5510) );
  GTECH_OR2 C9160 ( .A(N5508), .B(a4stg_rnd_frac[28]), .Z(N5509) );
  GTECH_OR2 C9161 ( .A(N5507), .B(a4stg_rnd_frac[29]), .Z(N5508) );
  GTECH_OR2 C9162 ( .A(N5506), .B(a4stg_rnd_frac[30]), .Z(N5507) );
  GTECH_OR2 C9163 ( .A(N5505), .B(a4stg_rnd_frac[31]), .Z(N5506) );
  GTECH_OR2 C9164 ( .A(N5504), .B(a4stg_rnd_frac[32]), .Z(N5505) );
  GTECH_OR2 C9165 ( .A(N5503), .B(a4stg_rnd_frac[33]), .Z(N5504) );
  GTECH_OR2 C9166 ( .A(N5502), .B(a4stg_rnd_frac[34]), .Z(N5503) );
  GTECH_OR2 C9167 ( .A(N5501), .B(a4stg_rnd_frac[35]), .Z(N5502) );
  GTECH_OR2 C9168 ( .A(N5500), .B(a4stg_rnd_frac[36]), .Z(N5501) );
  GTECH_OR2 C9169 ( .A(a4stg_rnd_frac[38]), .B(a4stg_rnd_frac[37]), .Z(N5500)
         );
  GTECH_OR2 C9170 ( .A(a4stg_frac_38_0_nx), .B(a4stg_rnd_frac_39), .Z(
        a4stg_frac_sng_nx) );
  GTECH_OR2 C9171 ( .A(a4stg_frac_sng_nx), .B(N5549), .Z(a4stg_frac_neq_0) );
  GTECH_OR2 C9172 ( .A(N5548), .B(a4stg_rnd_frac_40), .Z(N5549) );
  GTECH_OR2 C9173 ( .A(N5547), .B(a4stg_rnd_frac_41), .Z(N5548) );
  GTECH_OR2 C9174 ( .A(N5546), .B(a4stg_rnd_frac_42), .Z(N5547) );
  GTECH_OR2 C9175 ( .A(N5545), .B(a4stg_rnd_frac_43), .Z(N5546) );
  GTECH_OR2 C9176 ( .A(N5544), .B(a4stg_rnd_frac_44), .Z(N5545) );
  GTECH_OR2 C9177 ( .A(N5543), .B(a4stg_rnd_frac_45), .Z(N5544) );
  GTECH_OR2 C9178 ( .A(N5542), .B(a4stg_rnd_frac_46), .Z(N5543) );
  GTECH_OR2 C9179 ( .A(N5541), .B(a4stg_rnd_frac_47), .Z(N5542) );
  GTECH_OR2 C9180 ( .A(N5540), .B(a4stg_rnd_frac_48), .Z(N5541) );
  GTECH_OR2 C9181 ( .A(N5539), .B(a4stg_rnd_frac_49), .Z(N5540) );
  GTECH_OR2 C9182 ( .A(N5538), .B(a4stg_rnd_frac_50), .Z(N5539) );
  GTECH_OR2 C9183 ( .A(N5537), .B(a4stg_rnd_frac_51), .Z(N5538) );
  GTECH_OR2 C9184 ( .A(N5536), .B(a4stg_rnd_frac_52), .Z(N5537) );
  GTECH_OR2 C9185 ( .A(N5535), .B(a4stg_rnd_frac_53), .Z(N5536) );
  GTECH_OR2 C9186 ( .A(N5534), .B(a4stg_rnd_frac_54), .Z(N5535) );
  GTECH_OR2 C9187 ( .A(N5533), .B(a4stg_rnd_frac_55), .Z(N5534) );
  GTECH_OR2 C9188 ( .A(N5532), .B(a4stg_rnd_frac_56), .Z(N5533) );
  GTECH_OR2 C9189 ( .A(N5531), .B(a4stg_rnd_frac_57), .Z(N5532) );
  GTECH_OR2 C9190 ( .A(N5530), .B(a4stg_rnd_frac_58), .Z(N5531) );
  GTECH_OR2 C9191 ( .A(N5529), .B(a4stg_rnd_frac_59), .Z(N5530) );
  GTECH_OR2 C9192 ( .A(N5528), .B(a4stg_rnd_frac_60), .Z(N5529) );
  GTECH_OR2 C9193 ( .A(N5527), .B(a4stg_rnd_frac_61), .Z(N5528) );
  GTECH_OR2 C9194 ( .A(a4stg_rnd_frac_63), .B(a4stg_rnd_frac_62), .Z(N5527) );
  GTECH_OR2 C9195 ( .A(N5611), .B(a4stg_shl_data[0]), .Z(a4stg_shl_data_neq_0)
         );
  GTECH_OR2 C9196 ( .A(N5610), .B(a4stg_shl_data[1]), .Z(N5611) );
  GTECH_OR2 C9197 ( .A(N5609), .B(a4stg_shl_data[2]), .Z(N5610) );
  GTECH_OR2 C9198 ( .A(N5608), .B(a4stg_shl_data[3]), .Z(N5609) );
  GTECH_OR2 C9199 ( .A(N5607), .B(a4stg_shl_data[4]), .Z(N5608) );
  GTECH_OR2 C9200 ( .A(N5606), .B(a4stg_shl_data[5]), .Z(N5607) );
  GTECH_OR2 C9201 ( .A(N5605), .B(a4stg_shl_data[6]), .Z(N5606) );
  GTECH_OR2 C9202 ( .A(N5604), .B(a4stg_shl_data[7]), .Z(N5605) );
  GTECH_OR2 C9203 ( .A(N5603), .B(a4stg_shl_data[8]), .Z(N5604) );
  GTECH_OR2 C9204 ( .A(N5602), .B(a4stg_shl_data[9]), .Z(N5603) );
  GTECH_OR2 C9205 ( .A(N5601), .B(a4stg_shl_data[10]), .Z(N5602) );
  GTECH_OR2 C9206 ( .A(N5600), .B(a4stg_shl_data[11]), .Z(N5601) );
  GTECH_OR2 C9207 ( .A(N5599), .B(a4stg_shl_data[12]), .Z(N5600) );
  GTECH_OR2 C9208 ( .A(N5598), .B(a4stg_shl_data[13]), .Z(N5599) );
  GTECH_OR2 C9209 ( .A(N5597), .B(a4stg_shl_data[14]), .Z(N5598) );
  GTECH_OR2 C9210 ( .A(N5596), .B(a4stg_shl_data[15]), .Z(N5597) );
  GTECH_OR2 C9211 ( .A(N5595), .B(a4stg_shl_data[16]), .Z(N5596) );
  GTECH_OR2 C9212 ( .A(N5594), .B(a4stg_shl_data[17]), .Z(N5595) );
  GTECH_OR2 C9213 ( .A(N5593), .B(a4stg_shl_data[18]), .Z(N5594) );
  GTECH_OR2 C9214 ( .A(N5592), .B(a4stg_shl_data[19]), .Z(N5593) );
  GTECH_OR2 C9215 ( .A(N5591), .B(a4stg_shl_data[20]), .Z(N5592) );
  GTECH_OR2 C9216 ( .A(N5590), .B(a4stg_shl_data[21]), .Z(N5591) );
  GTECH_OR2 C9217 ( .A(N5589), .B(a4stg_shl_data[22]), .Z(N5590) );
  GTECH_OR2 C9218 ( .A(N5588), .B(a4stg_shl_data[23]), .Z(N5589) );
  GTECH_OR2 C9219 ( .A(N5587), .B(a4stg_shl_data[24]), .Z(N5588) );
  GTECH_OR2 C9220 ( .A(N5586), .B(a4stg_shl_data[25]), .Z(N5587) );
  GTECH_OR2 C9221 ( .A(N5585), .B(a4stg_shl_data[26]), .Z(N5586) );
  GTECH_OR2 C9222 ( .A(N5584), .B(a4stg_shl_data[27]), .Z(N5585) );
  GTECH_OR2 C9223 ( .A(N5583), .B(a4stg_shl_data[28]), .Z(N5584) );
  GTECH_OR2 C9224 ( .A(N5582), .B(a4stg_shl_data[29]), .Z(N5583) );
  GTECH_OR2 C9225 ( .A(N5581), .B(a4stg_shl_data[30]), .Z(N5582) );
  GTECH_OR2 C9226 ( .A(N5580), .B(a4stg_shl_data[31]), .Z(N5581) );
  GTECH_OR2 C9227 ( .A(N5579), .B(a4stg_shl_data[32]), .Z(N5580) );
  GTECH_OR2 C9228 ( .A(N5578), .B(a4stg_shl_data[33]), .Z(N5579) );
  GTECH_OR2 C9229 ( .A(N5577), .B(a4stg_shl_data[34]), .Z(N5578) );
  GTECH_OR2 C9230 ( .A(N5576), .B(a4stg_shl_data[35]), .Z(N5577) );
  GTECH_OR2 C9231 ( .A(N5575), .B(a4stg_shl_data[36]), .Z(N5576) );
  GTECH_OR2 C9232 ( .A(N5574), .B(a4stg_shl_data[37]), .Z(N5575) );
  GTECH_OR2 C9233 ( .A(N5573), .B(a4stg_shl_data[38]), .Z(N5574) );
  GTECH_OR2 C9234 ( .A(N5572), .B(a4stg_shl_data[39]), .Z(N5573) );
  GTECH_OR2 C9235 ( .A(N5571), .B(a4stg_shl_data[40]), .Z(N5572) );
  GTECH_OR2 C9236 ( .A(N5570), .B(a4stg_shl_data[41]), .Z(N5571) );
  GTECH_OR2 C9237 ( .A(N5569), .B(a4stg_shl_data[42]), .Z(N5570) );
  GTECH_OR2 C9238 ( .A(N5568), .B(a4stg_shl_data[43]), .Z(N5569) );
  GTECH_OR2 C9239 ( .A(N5567), .B(a4stg_shl_data[44]), .Z(N5568) );
  GTECH_OR2 C9240 ( .A(N5566), .B(a4stg_shl_data[45]), .Z(N5567) );
  GTECH_OR2 C9241 ( .A(N5565), .B(a4stg_shl_data[46]), .Z(N5566) );
  GTECH_OR2 C9242 ( .A(N5564), .B(a4stg_shl_data[47]), .Z(N5565) );
  GTECH_OR2 C9243 ( .A(N5563), .B(a4stg_shl_data[48]), .Z(N5564) );
  GTECH_OR2 C9244 ( .A(N5562), .B(a4stg_shl_data[49]), .Z(N5563) );
  GTECH_OR2 C9245 ( .A(N5561), .B(a4stg_shl_data[50]), .Z(N5562) );
  GTECH_OR2 C9246 ( .A(N5560), .B(a4stg_shl_data[51]), .Z(N5561) );
  GTECH_OR2 C9247 ( .A(N5559), .B(a4stg_shl_data[52]), .Z(N5560) );
  GTECH_OR2 C9248 ( .A(N5558), .B(a4stg_shl_data[53]), .Z(N5559) );
  GTECH_OR2 C9249 ( .A(N5557), .B(a4stg_shl_data[54]), .Z(N5558) );
  GTECH_OR2 C9250 ( .A(N5556), .B(a4stg_shl_data[55]), .Z(N5557) );
  GTECH_OR2 C9251 ( .A(N5555), .B(a4stg_shl_data[56]), .Z(N5556) );
  GTECH_OR2 C9252 ( .A(N5554), .B(a4stg_shl_data[57]), .Z(N5555) );
  GTECH_OR2 C9253 ( .A(N5553), .B(a4stg_shl_data[58]), .Z(N5554) );
  GTECH_OR2 C9254 ( .A(N5552), .B(a4stg_shl_data[59]), .Z(N5553) );
  GTECH_OR2 C9255 ( .A(N5551), .B(a4stg_shl_data[60]), .Z(N5552) );
  GTECH_OR2 C9256 ( .A(N5550), .B(a4stg_shl_data[61]), .Z(N5551) );
  GTECH_OR2 C9257 ( .A(a4stg_shl_data[63]), .B(a4stg_shl_data[62]), .Z(N5550)
         );
  GTECH_OR2 C9258 ( .A(N5616), .B(N5617), .Z(a4stg_shl_tmp4[63]) );
  GTECH_OR2 C9259 ( .A(N5614), .B(N5615), .Z(N5616) );
  GTECH_OR2 C9260 ( .A(N5612), .B(N5613), .Z(N5614) );
  GTECH_AND2 C9261 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[63]), .Z(
        N5612) );
  GTECH_AND2 C9262 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[47]), .Z(
        N5613) );
  GTECH_AND2 C9263 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[31]), .Z(
        N5615) );
  GTECH_AND2 C9264 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[15]), .Z(
        N5617) );
  GTECH_OR2 C9265 ( .A(N5622), .B(N5623), .Z(a4stg_shl_tmp4[62]) );
  GTECH_OR2 C9266 ( .A(N5620), .B(N5621), .Z(N5622) );
  GTECH_OR2 C9267 ( .A(N5618), .B(N5619), .Z(N5620) );
  GTECH_AND2 C9268 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[62]), .Z(
        N5618) );
  GTECH_AND2 C9269 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[46]), .Z(
        N5619) );
  GTECH_AND2 C9270 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[30]), .Z(
        N5621) );
  GTECH_AND2 C9271 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[14]), .Z(
        N5623) );
  GTECH_OR2 C9272 ( .A(N5628), .B(N5629), .Z(a4stg_shl_tmp4[61]) );
  GTECH_OR2 C9273 ( .A(N5626), .B(N5627), .Z(N5628) );
  GTECH_OR2 C9274 ( .A(N5624), .B(N5625), .Z(N5626) );
  GTECH_AND2 C9275 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[61]), .Z(
        N5624) );
  GTECH_AND2 C9276 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[45]), .Z(
        N5625) );
  GTECH_AND2 C9277 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[29]), .Z(
        N5627) );
  GTECH_AND2 C9278 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[13]), .Z(
        N5629) );
  GTECH_OR2 C9279 ( .A(N5634), .B(N5635), .Z(a4stg_shl_tmp4[60]) );
  GTECH_OR2 C9280 ( .A(N5632), .B(N5633), .Z(N5634) );
  GTECH_OR2 C9281 ( .A(N5630), .B(N5631), .Z(N5632) );
  GTECH_AND2 C9282 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[60]), .Z(
        N5630) );
  GTECH_AND2 C9283 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[44]), .Z(
        N5631) );
  GTECH_AND2 C9284 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[28]), .Z(
        N5633) );
  GTECH_AND2 C9285 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[12]), .Z(
        N5635) );
  GTECH_OR2 C9286 ( .A(N5640), .B(N5641), .Z(a4stg_shl_tmp4[59]) );
  GTECH_OR2 C9287 ( .A(N5638), .B(N5639), .Z(N5640) );
  GTECH_OR2 C9288 ( .A(N5636), .B(N5637), .Z(N5638) );
  GTECH_AND2 C9289 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[59]), .Z(
        N5636) );
  GTECH_AND2 C9290 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[43]), .Z(
        N5637) );
  GTECH_AND2 C9291 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[27]), .Z(
        N5639) );
  GTECH_AND2 C9292 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[11]), .Z(
        N5641) );
  GTECH_OR2 C9293 ( .A(N5646), .B(N5647), .Z(a4stg_shl_tmp4[58]) );
  GTECH_OR2 C9294 ( .A(N5644), .B(N5645), .Z(N5646) );
  GTECH_OR2 C9295 ( .A(N5642), .B(N5643), .Z(N5644) );
  GTECH_AND2 C9296 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[58]), .Z(
        N5642) );
  GTECH_AND2 C9297 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[42]), .Z(
        N5643) );
  GTECH_AND2 C9298 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[26]), .Z(
        N5645) );
  GTECH_AND2 C9299 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[10]), .Z(
        N5647) );
  GTECH_OR2 C9300 ( .A(N5652), .B(N5653), .Z(a4stg_shl_tmp4[57]) );
  GTECH_OR2 C9301 ( .A(N5650), .B(N5651), .Z(N5652) );
  GTECH_OR2 C9302 ( .A(N5648), .B(N5649), .Z(N5650) );
  GTECH_AND2 C9303 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[57]), .Z(
        N5648) );
  GTECH_AND2 C9304 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[41]), .Z(
        N5649) );
  GTECH_AND2 C9305 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[25]), .Z(
        N5651) );
  GTECH_AND2 C9306 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[9]), .Z(
        N5653) );
  GTECH_OR2 C9307 ( .A(N5658), .B(N5659), .Z(a4stg_shl_tmp4[56]) );
  GTECH_OR2 C9308 ( .A(N5656), .B(N5657), .Z(N5658) );
  GTECH_OR2 C9309 ( .A(N5654), .B(N5655), .Z(N5656) );
  GTECH_AND2 C9310 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[56]), .Z(
        N5654) );
  GTECH_AND2 C9311 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[40]), .Z(
        N5655) );
  GTECH_AND2 C9312 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[24]), .Z(
        N5657) );
  GTECH_AND2 C9313 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[8]), .Z(
        N5659) );
  GTECH_OR2 C9314 ( .A(N5664), .B(N5665), .Z(a4stg_shl_tmp4[55]) );
  GTECH_OR2 C9315 ( .A(N5662), .B(N5663), .Z(N5664) );
  GTECH_OR2 C9316 ( .A(N5660), .B(N5661), .Z(N5662) );
  GTECH_AND2 C9317 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[55]), .Z(
        N5660) );
  GTECH_AND2 C9318 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[39]), .Z(
        N5661) );
  GTECH_AND2 C9319 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[23]), .Z(
        N5663) );
  GTECH_AND2 C9320 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[7]), .Z(
        N5665) );
  GTECH_OR2 C9321 ( .A(N5670), .B(N5671), .Z(a4stg_shl_tmp4[54]) );
  GTECH_OR2 C9322 ( .A(N5668), .B(N5669), .Z(N5670) );
  GTECH_OR2 C9323 ( .A(N5666), .B(N5667), .Z(N5668) );
  GTECH_AND2 C9324 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[54]), .Z(
        N5666) );
  GTECH_AND2 C9325 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[38]), .Z(
        N5667) );
  GTECH_AND2 C9326 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[22]), .Z(
        N5669) );
  GTECH_AND2 C9327 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[6]), .Z(
        N5671) );
  GTECH_OR2 C9328 ( .A(N5676), .B(N5677), .Z(a4stg_shl_tmp4[53]) );
  GTECH_OR2 C9329 ( .A(N5674), .B(N5675), .Z(N5676) );
  GTECH_OR2 C9330 ( .A(N5672), .B(N5673), .Z(N5674) );
  GTECH_AND2 C9331 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[53]), .Z(
        N5672) );
  GTECH_AND2 C9332 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[37]), .Z(
        N5673) );
  GTECH_AND2 C9333 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[21]), .Z(
        N5675) );
  GTECH_AND2 C9334 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[5]), .Z(
        N5677) );
  GTECH_OR2 C9335 ( .A(N5682), .B(N5683), .Z(a4stg_shl_tmp4[52]) );
  GTECH_OR2 C9336 ( .A(N5680), .B(N5681), .Z(N5682) );
  GTECH_OR2 C9337 ( .A(N5678), .B(N5679), .Z(N5680) );
  GTECH_AND2 C9338 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[52]), .Z(
        N5678) );
  GTECH_AND2 C9339 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[36]), .Z(
        N5679) );
  GTECH_AND2 C9340 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[20]), .Z(
        N5681) );
  GTECH_AND2 C9341 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[4]), .Z(
        N5683) );
  GTECH_OR2 C9342 ( .A(N5688), .B(N5689), .Z(a4stg_shl_tmp4[51]) );
  GTECH_OR2 C9343 ( .A(N5686), .B(N5687), .Z(N5688) );
  GTECH_OR2 C9344 ( .A(N5684), .B(N5685), .Z(N5686) );
  GTECH_AND2 C9345 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[51]), .Z(
        N5684) );
  GTECH_AND2 C9346 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[35]), .Z(
        N5685) );
  GTECH_AND2 C9347 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[19]), .Z(
        N5687) );
  GTECH_AND2 C9348 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[3]), .Z(
        N5689) );
  GTECH_OR2 C9349 ( .A(N5694), .B(N5695), .Z(a4stg_shl_tmp4[50]) );
  GTECH_OR2 C9350 ( .A(N5692), .B(N5693), .Z(N5694) );
  GTECH_OR2 C9351 ( .A(N5690), .B(N5691), .Z(N5692) );
  GTECH_AND2 C9352 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[50]), .Z(
        N5690) );
  GTECH_AND2 C9353 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[34]), .Z(
        N5691) );
  GTECH_AND2 C9354 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[18]), .Z(
        N5693) );
  GTECH_AND2 C9355 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[2]), .Z(
        N5695) );
  GTECH_OR2 C9356 ( .A(N5700), .B(N5701), .Z(a4stg_shl_tmp4[49]) );
  GTECH_OR2 C9357 ( .A(N5698), .B(N5699), .Z(N5700) );
  GTECH_OR2 C9358 ( .A(N5696), .B(N5697), .Z(N5698) );
  GTECH_AND2 C9359 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[49]), .Z(
        N5696) );
  GTECH_AND2 C9360 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[33]), .Z(
        N5697) );
  GTECH_AND2 C9361 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[17]), .Z(
        N5699) );
  GTECH_AND2 C9362 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[1]), .Z(
        N5701) );
  GTECH_OR2 C9363 ( .A(N5706), .B(N5707), .Z(a4stg_shl_tmp4[48]) );
  GTECH_OR2 C9364 ( .A(N5704), .B(N5705), .Z(N5706) );
  GTECH_OR2 C9365 ( .A(N5702), .B(N5703), .Z(N5704) );
  GTECH_AND2 C9366 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[48]), .Z(
        N5702) );
  GTECH_AND2 C9367 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[32]), .Z(
        N5703) );
  GTECH_AND2 C9368 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[16]), .Z(
        N5705) );
  GTECH_AND2 C9369 ( .A(a4stg_shl_cnt_dec54_3[0]), .B(a4stg_shl_data[0]), .Z(
        N5707) );
  GTECH_OR2 C9370 ( .A(N5710), .B(N5711), .Z(a4stg_shl_tmp4[47]) );
  GTECH_OR2 C9371 ( .A(N5708), .B(N5709), .Z(N5710) );
  GTECH_AND2 C9372 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[47]), .Z(
        N5708) );
  GTECH_AND2 C9373 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[31]), .Z(
        N5709) );
  GTECH_AND2 C9374 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[15]), .Z(
        N5711) );
  GTECH_OR2 C9375 ( .A(N5714), .B(N5715), .Z(a4stg_shl_tmp4[46]) );
  GTECH_OR2 C9376 ( .A(N5712), .B(N5713), .Z(N5714) );
  GTECH_AND2 C9377 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[46]), .Z(
        N5712) );
  GTECH_AND2 C9378 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[30]), .Z(
        N5713) );
  GTECH_AND2 C9379 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[14]), .Z(
        N5715) );
  GTECH_OR2 C9380 ( .A(N5718), .B(N5719), .Z(a4stg_shl_tmp4[45]) );
  GTECH_OR2 C9381 ( .A(N5716), .B(N5717), .Z(N5718) );
  GTECH_AND2 C9382 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[45]), .Z(
        N5716) );
  GTECH_AND2 C9383 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[29]), .Z(
        N5717) );
  GTECH_AND2 C9384 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[13]), .Z(
        N5719) );
  GTECH_OR2 C9385 ( .A(N5722), .B(N5723), .Z(a4stg_shl_tmp4[44]) );
  GTECH_OR2 C9386 ( .A(N5720), .B(N5721), .Z(N5722) );
  GTECH_AND2 C9387 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[44]), .Z(
        N5720) );
  GTECH_AND2 C9388 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[28]), .Z(
        N5721) );
  GTECH_AND2 C9389 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[12]), .Z(
        N5723) );
  GTECH_OR2 C9390 ( .A(N5726), .B(N5727), .Z(a4stg_shl_tmp4[43]) );
  GTECH_OR2 C9391 ( .A(N5724), .B(N5725), .Z(N5726) );
  GTECH_AND2 C9392 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[43]), .Z(
        N5724) );
  GTECH_AND2 C9393 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[27]), .Z(
        N5725) );
  GTECH_AND2 C9394 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[11]), .Z(
        N5727) );
  GTECH_OR2 C9395 ( .A(N5730), .B(N5731), .Z(a4stg_shl_tmp4[42]) );
  GTECH_OR2 C9396 ( .A(N5728), .B(N5729), .Z(N5730) );
  GTECH_AND2 C9397 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[42]), .Z(
        N5728) );
  GTECH_AND2 C9398 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[26]), .Z(
        N5729) );
  GTECH_AND2 C9399 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[10]), .Z(
        N5731) );
  GTECH_OR2 C9400 ( .A(N5734), .B(N5735), .Z(a4stg_shl_tmp4[41]) );
  GTECH_OR2 C9401 ( .A(N5732), .B(N5733), .Z(N5734) );
  GTECH_AND2 C9402 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[41]), .Z(
        N5732) );
  GTECH_AND2 C9403 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[25]), .Z(
        N5733) );
  GTECH_AND2 C9404 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[9]), .Z(
        N5735) );
  GTECH_OR2 C9405 ( .A(N5738), .B(N5739), .Z(a4stg_shl_tmp4[40]) );
  GTECH_OR2 C9406 ( .A(N5736), .B(N5737), .Z(N5738) );
  GTECH_AND2 C9407 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[40]), .Z(
        N5736) );
  GTECH_AND2 C9408 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[24]), .Z(
        N5737) );
  GTECH_AND2 C9409 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[8]), .Z(
        N5739) );
  GTECH_OR2 C9410 ( .A(N5742), .B(N5743), .Z(a4stg_shl_tmp4[39]) );
  GTECH_OR2 C9411 ( .A(N5740), .B(N5741), .Z(N5742) );
  GTECH_AND2 C9412 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[39]), .Z(
        N5740) );
  GTECH_AND2 C9413 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[23]), .Z(
        N5741) );
  GTECH_AND2 C9414 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[7]), .Z(
        N5743) );
  GTECH_OR2 C9415 ( .A(N5746), .B(N5747), .Z(a4stg_shl_tmp4[38]) );
  GTECH_OR2 C9416 ( .A(N5744), .B(N5745), .Z(N5746) );
  GTECH_AND2 C9417 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[38]), .Z(
        N5744) );
  GTECH_AND2 C9418 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[22]), .Z(
        N5745) );
  GTECH_AND2 C9419 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[6]), .Z(
        N5747) );
  GTECH_OR2 C9420 ( .A(N5750), .B(N5751), .Z(a4stg_shl_tmp4[37]) );
  GTECH_OR2 C9421 ( .A(N5748), .B(N5749), .Z(N5750) );
  GTECH_AND2 C9422 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[37]), .Z(
        N5748) );
  GTECH_AND2 C9423 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[21]), .Z(
        N5749) );
  GTECH_AND2 C9424 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[5]), .Z(
        N5751) );
  GTECH_OR2 C9425 ( .A(N5754), .B(N5755), .Z(a4stg_shl_tmp4[36]) );
  GTECH_OR2 C9426 ( .A(N5752), .B(N5753), .Z(N5754) );
  GTECH_AND2 C9427 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[36]), .Z(
        N5752) );
  GTECH_AND2 C9428 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[20]), .Z(
        N5753) );
  GTECH_AND2 C9429 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[4]), .Z(
        N5755) );
  GTECH_OR2 C9430 ( .A(N5758), .B(N5759), .Z(a4stg_shl_tmp4[35]) );
  GTECH_OR2 C9431 ( .A(N5756), .B(N5757), .Z(N5758) );
  GTECH_AND2 C9432 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[35]), .Z(
        N5756) );
  GTECH_AND2 C9433 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[19]), .Z(
        N5757) );
  GTECH_AND2 C9434 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[3]), .Z(
        N5759) );
  GTECH_OR2 C9435 ( .A(N5762), .B(N5763), .Z(a4stg_shl_tmp4[34]) );
  GTECH_OR2 C9436 ( .A(N5760), .B(N5761), .Z(N5762) );
  GTECH_AND2 C9437 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[34]), .Z(
        N5760) );
  GTECH_AND2 C9438 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[18]), .Z(
        N5761) );
  GTECH_AND2 C9439 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[2]), .Z(
        N5763) );
  GTECH_OR2 C9440 ( .A(N5766), .B(N5767), .Z(a4stg_shl_tmp4[33]) );
  GTECH_OR2 C9441 ( .A(N5764), .B(N5765), .Z(N5766) );
  GTECH_AND2 C9442 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[33]), .Z(
        N5764) );
  GTECH_AND2 C9443 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[17]), .Z(
        N5765) );
  GTECH_AND2 C9444 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[1]), .Z(
        N5767) );
  GTECH_OR2 C9445 ( .A(N5770), .B(N5771), .Z(a4stg_shl_tmp4[32]) );
  GTECH_OR2 C9446 ( .A(N5768), .B(N5769), .Z(N5770) );
  GTECH_AND2 C9447 ( .A(a4stg_shl_cnt_dec54_0[0]), .B(a4stg_shl_data[32]), .Z(
        N5768) );
  GTECH_AND2 C9448 ( .A(a4stg_shl_cnt_dec54_1[0]), .B(a4stg_shl_data[16]), .Z(
        N5769) );
  GTECH_AND2 C9449 ( .A(a4stg_shl_cnt_dec54_2[0]), .B(a4stg_shl_data[0]), .Z(
        N5771) );
  GTECH_OR2 C9450 ( .A(N5772), .B(N5773), .Z(a4stg_shl_tmp4[31]) );
  GTECH_AND2 C9451 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[31]), .Z(
        N5772) );
  GTECH_AND2 C9452 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[15]), .Z(
        N5773) );
  GTECH_OR2 C9453 ( .A(N5774), .B(N5775), .Z(a4stg_shl_tmp4[30]) );
  GTECH_AND2 C9454 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[30]), .Z(
        N5774) );
  GTECH_AND2 C9455 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[14]), .Z(
        N5775) );
  GTECH_OR2 C9456 ( .A(N5776), .B(N5777), .Z(a4stg_shl_tmp4[29]) );
  GTECH_AND2 C9457 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[29]), .Z(
        N5776) );
  GTECH_AND2 C9458 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[13]), .Z(
        N5777) );
  GTECH_OR2 C9459 ( .A(N5778), .B(N5779), .Z(a4stg_shl_tmp4[28]) );
  GTECH_AND2 C9460 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[28]), .Z(
        N5778) );
  GTECH_AND2 C9461 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[12]), .Z(
        N5779) );
  GTECH_OR2 C9462 ( .A(N5780), .B(N5781), .Z(a4stg_shl_tmp4[27]) );
  GTECH_AND2 C9463 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[27]), .Z(
        N5780) );
  GTECH_AND2 C9464 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[11]), .Z(
        N5781) );
  GTECH_OR2 C9465 ( .A(N5782), .B(N5783), .Z(a4stg_shl_tmp4[26]) );
  GTECH_AND2 C9466 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[26]), .Z(
        N5782) );
  GTECH_AND2 C9467 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[10]), .Z(
        N5783) );
  GTECH_OR2 C9468 ( .A(N5784), .B(N5785), .Z(a4stg_shl_tmp4[25]) );
  GTECH_AND2 C9469 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[25]), .Z(
        N5784) );
  GTECH_AND2 C9470 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[9]), .Z(
        N5785) );
  GTECH_OR2 C9471 ( .A(N5786), .B(N5787), .Z(a4stg_shl_tmp4[24]) );
  GTECH_AND2 C9472 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[24]), .Z(
        N5786) );
  GTECH_AND2 C9473 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[8]), .Z(
        N5787) );
  GTECH_OR2 C9474 ( .A(N5788), .B(N5789), .Z(a4stg_shl_tmp4[23]) );
  GTECH_AND2 C9475 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[23]), .Z(
        N5788) );
  GTECH_AND2 C9476 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[7]), .Z(
        N5789) );
  GTECH_OR2 C9477 ( .A(N5790), .B(N5791), .Z(a4stg_shl_tmp4[22]) );
  GTECH_AND2 C9478 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[22]), .Z(
        N5790) );
  GTECH_AND2 C9479 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[6]), .Z(
        N5791) );
  GTECH_OR2 C9480 ( .A(N5792), .B(N5793), .Z(a4stg_shl_tmp4[21]) );
  GTECH_AND2 C9481 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[21]), .Z(
        N5792) );
  GTECH_AND2 C9482 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[5]), .Z(
        N5793) );
  GTECH_OR2 C9483 ( .A(N5794), .B(N5795), .Z(a4stg_shl_tmp4[20]) );
  GTECH_AND2 C9484 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[20]), .Z(
        N5794) );
  GTECH_AND2 C9485 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[4]), .Z(
        N5795) );
  GTECH_OR2 C9486 ( .A(N5796), .B(N5797), .Z(a4stg_shl_tmp4[19]) );
  GTECH_AND2 C9487 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[19]), .Z(
        N5796) );
  GTECH_AND2 C9488 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[3]), .Z(
        N5797) );
  GTECH_OR2 C9489 ( .A(N5798), .B(N5799), .Z(a4stg_shl_tmp4[18]) );
  GTECH_AND2 C9490 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[18]), .Z(
        N5798) );
  GTECH_AND2 C9491 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[2]), .Z(
        N5799) );
  GTECH_OR2 C9492 ( .A(N5800), .B(N5801), .Z(a4stg_shl_tmp4[17]) );
  GTECH_AND2 C9493 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[17]), .Z(
        N5800) );
  GTECH_AND2 C9494 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[1]), .Z(
        N5801) );
  GTECH_OR2 C9495 ( .A(N5802), .B(N5803), .Z(a4stg_shl_tmp4[16]) );
  GTECH_AND2 C9496 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[16]), .Z(
        N5802) );
  GTECH_AND2 C9497 ( .A(a4stg_shl_cnt_dec54_1[1]), .B(a4stg_shl_data[0]), .Z(
        N5803) );
  GTECH_AND2 C9498 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[15]), .Z(
        a4stg_shl_tmp4[15]) );
  GTECH_AND2 C9499 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[14]), .Z(
        a4stg_shl_tmp4[14]) );
  GTECH_AND2 C9500 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[13]), .Z(
        a4stg_shl_tmp4[13]) );
  GTECH_AND2 C9501 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[12]), .Z(
        a4stg_shl_tmp4[12]) );
  GTECH_AND2 C9502 ( .A(a4stg_shl_cnt_dec54_0[1]), .B(a4stg_shl_data[11]), .Z(
        a4stg_shl_tmp4[11]) );
  GTECH_AND2 C9503 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[10]), .Z(
        a4stg_shl_tmp4[10]) );
  GTECH_AND2 C9504 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[9]), .Z(
        a4stg_shl_tmp4[9]) );
  GTECH_AND2 C9505 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[8]), .Z(
        a4stg_shl_tmp4[8]) );
  GTECH_AND2 C9506 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[7]), .Z(
        a4stg_shl_tmp4[7]) );
  GTECH_AND2 C9507 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[6]), .Z(
        a4stg_shl_tmp4[6]) );
  GTECH_AND2 C9508 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[5]), .Z(
        a4stg_shl_tmp4[5]) );
  GTECH_AND2 C9509 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[4]), .Z(
        a4stg_shl_tmp4[4]) );
  GTECH_AND2 C9510 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[3]), .Z(
        a4stg_shl_tmp4[3]) );
  GTECH_AND2 C9511 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[2]), .Z(
        a4stg_shl_tmp4[2]) );
  GTECH_AND2 C9512 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[1]), .Z(
        a4stg_shl_tmp4[1]) );
  GTECH_AND2 C9513 ( .A(a4stg_shl_cnt_dec54_0[2]), .B(a4stg_shl_data[0]), .Z(
        a4stg_shl_tmp4[0]) );
  GTECH_OR2 C9514 ( .A(N5806), .B(N5807), .Z(add_frac_out[63]) );
  GTECH_OR2 C9515 ( .A(N5804), .B(N5805), .Z(N5806) );
  GTECH_AND2 C9516 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[63]), .Z(
        N5804) );
  GTECH_AND2 C9517 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5805) );
  GTECH_AND2 C9518 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[63]), .Z(N5807) );
  GTECH_OR2 C9519 ( .A(N5812), .B(N5813), .Z(add_frac_out[62]) );
  GTECH_OR2 C9520 ( .A(N5810), .B(N5811), .Z(N5812) );
  GTECH_OR2 C9521 ( .A(N5808), .B(N5809), .Z(N5810) );
  GTECH_AND2 C9522 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[51]), .Z(N5808) );
  GTECH_AND2 C9523 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[62]), .Z(
        N5809) );
  GTECH_AND2 C9524 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5811) );
  GTECH_AND2 C9525 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[62]), .Z(N5813) );
  GTECH_OR2 C9526 ( .A(N5818), .B(N5819), .Z(add_frac_out[61]) );
  GTECH_OR2 C9527 ( .A(N5816), .B(N5817), .Z(N5818) );
  GTECH_OR2 C9528 ( .A(N5814), .B(N5815), .Z(N5816) );
  GTECH_AND2 C9529 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[50]), .Z(N5814) );
  GTECH_AND2 C9530 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[61]), .Z(
        N5815) );
  GTECH_AND2 C9531 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5817) );
  GTECH_AND2 C9532 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[61]), .Z(N5819) );
  GTECH_OR2 C9533 ( .A(N5824), .B(N5825), .Z(add_frac_out[60]) );
  GTECH_OR2 C9534 ( .A(N5822), .B(N5823), .Z(N5824) );
  GTECH_OR2 C9535 ( .A(N5820), .B(N5821), .Z(N5822) );
  GTECH_AND2 C9536 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[49]), .Z(N5820) );
  GTECH_AND2 C9537 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[60]), .Z(
        N5821) );
  GTECH_AND2 C9538 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5823) );
  GTECH_AND2 C9539 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[60]), .Z(N5825) );
  GTECH_OR2 C9540 ( .A(N5830), .B(N5831), .Z(add_frac_out[59]) );
  GTECH_OR2 C9541 ( .A(N5828), .B(N5829), .Z(N5830) );
  GTECH_OR2 C9542 ( .A(N5826), .B(N5827), .Z(N5828) );
  GTECH_AND2 C9543 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[48]), .Z(N5826) );
  GTECH_AND2 C9544 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[59]), .Z(
        N5827) );
  GTECH_AND2 C9545 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5829) );
  GTECH_AND2 C9546 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[59]), .Z(N5831) );
  GTECH_OR2 C9547 ( .A(N5836), .B(N5837), .Z(add_frac_out[58]) );
  GTECH_OR2 C9548 ( .A(N5834), .B(N5835), .Z(N5836) );
  GTECH_OR2 C9549 ( .A(N5832), .B(N5833), .Z(N5834) );
  GTECH_AND2 C9550 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[47]), .Z(N5832) );
  GTECH_AND2 C9551 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[58]), .Z(
        N5833) );
  GTECH_AND2 C9552 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5835) );
  GTECH_AND2 C9553 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[58]), .Z(N5837) );
  GTECH_OR2 C9554 ( .A(N5842), .B(N5843), .Z(add_frac_out[57]) );
  GTECH_OR2 C9555 ( .A(N5840), .B(N5841), .Z(N5842) );
  GTECH_OR2 C9556 ( .A(N5838), .B(N5839), .Z(N5840) );
  GTECH_AND2 C9557 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[46]), .Z(N5838) );
  GTECH_AND2 C9558 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[57]), .Z(
        N5839) );
  GTECH_AND2 C9559 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5841) );
  GTECH_AND2 C9560 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[57]), .Z(N5843) );
  GTECH_OR2 C9561 ( .A(N5848), .B(N5849), .Z(add_frac_out[56]) );
  GTECH_OR2 C9562 ( .A(N5846), .B(N5847), .Z(N5848) );
  GTECH_OR2 C9563 ( .A(N5844), .B(N5845), .Z(N5846) );
  GTECH_AND2 C9564 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[45]), .Z(N5844) );
  GTECH_AND2 C9565 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[56]), .Z(
        N5845) );
  GTECH_AND2 C9566 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5847) );
  GTECH_AND2 C9567 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[56]), .Z(N5849) );
  GTECH_OR2 C9568 ( .A(N5854), .B(N5855), .Z(add_frac_out[55]) );
  GTECH_OR2 C9569 ( .A(N5852), .B(N5853), .Z(N5854) );
  GTECH_OR2 C9570 ( .A(N5850), .B(N5851), .Z(N5852) );
  GTECH_AND2 C9571 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[44]), .Z(N5850) );
  GTECH_AND2 C9572 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[55]), .Z(
        N5851) );
  GTECH_AND2 C9573 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5853) );
  GTECH_AND2 C9574 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[55]), .Z(N5855) );
  GTECH_OR2 C9575 ( .A(N5860), .B(N5861), .Z(add_frac_out[54]) );
  GTECH_OR2 C9576 ( .A(N5858), .B(N5859), .Z(N5860) );
  GTECH_OR2 C9577 ( .A(N5856), .B(N5857), .Z(N5858) );
  GTECH_AND2 C9578 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[43]), .Z(N5856) );
  GTECH_AND2 C9579 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[54]), .Z(
        N5857) );
  GTECH_AND2 C9580 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5859) );
  GTECH_AND2 C9581 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[54]), .Z(N5861) );
  GTECH_OR2 C9582 ( .A(N5866), .B(N5867), .Z(add_frac_out[53]) );
  GTECH_OR2 C9583 ( .A(N5864), .B(N5865), .Z(N5866) );
  GTECH_OR2 C9584 ( .A(N5862), .B(N5863), .Z(N5864) );
  GTECH_AND2 C9585 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[42]), .Z(N5862) );
  GTECH_AND2 C9586 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[53]), .Z(
        N5863) );
  GTECH_AND2 C9587 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5865) );
  GTECH_AND2 C9588 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[53]), .Z(N5867) );
  GTECH_OR2 C9589 ( .A(N5872), .B(N5873), .Z(add_frac_out[52]) );
  GTECH_OR2 C9590 ( .A(N5870), .B(N5871), .Z(N5872) );
  GTECH_OR2 C9591 ( .A(N5868), .B(N5869), .Z(N5870) );
  GTECH_AND2 C9592 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[41]), .Z(N5868) );
  GTECH_AND2 C9593 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[52]), .Z(
        N5869) );
  GTECH_AND2 C9594 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5871) );
  GTECH_AND2 C9595 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[52]), .Z(N5873) );
  GTECH_OR2 C9596 ( .A(N5878), .B(N5879), .Z(add_frac_out[51]) );
  GTECH_OR2 C9597 ( .A(N5876), .B(N5877), .Z(N5878) );
  GTECH_OR2 C9598 ( .A(N5874), .B(N5875), .Z(N5876) );
  GTECH_AND2 C9599 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[40]), .Z(N5874) );
  GTECH_AND2 C9600 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[51]), .Z(
        N5875) );
  GTECH_AND2 C9601 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5877) );
  GTECH_AND2 C9602 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[51]), .Z(N5879) );
  GTECH_OR2 C9603 ( .A(N5884), .B(N5885), .Z(add_frac_out[50]) );
  GTECH_OR2 C9604 ( .A(N5882), .B(N5883), .Z(N5884) );
  GTECH_OR2 C9605 ( .A(N5880), .B(N5881), .Z(N5882) );
  GTECH_AND2 C9606 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[39]), .Z(N5880) );
  GTECH_AND2 C9607 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[50]), .Z(
        N5881) );
  GTECH_AND2 C9608 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5883) );
  GTECH_AND2 C9609 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[50]), .Z(N5885) );
  GTECH_OR2 C9610 ( .A(N5890), .B(N5891), .Z(add_frac_out[49]) );
  GTECH_OR2 C9611 ( .A(N5888), .B(N5889), .Z(N5890) );
  GTECH_OR2 C9612 ( .A(N5886), .B(N5887), .Z(N5888) );
  GTECH_AND2 C9613 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[38]), .Z(N5886) );
  GTECH_AND2 C9614 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[49]), .Z(
        N5887) );
  GTECH_AND2 C9615 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5889) );
  GTECH_AND2 C9616 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[49]), .Z(N5891) );
  GTECH_OR2 C9617 ( .A(N5896), .B(N5897), .Z(add_frac_out[48]) );
  GTECH_OR2 C9618 ( .A(N5894), .B(N5895), .Z(N5896) );
  GTECH_OR2 C9619 ( .A(N5892), .B(N5893), .Z(N5894) );
  GTECH_AND2 C9620 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[37]), .Z(N5892) );
  GTECH_AND2 C9621 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[48]), .Z(
        N5893) );
  GTECH_AND2 C9622 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5895) );
  GTECH_AND2 C9623 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[48]), .Z(N5897) );
  GTECH_OR2 C9624 ( .A(N5902), .B(N5903), .Z(add_frac_out[47]) );
  GTECH_OR2 C9625 ( .A(N5900), .B(N5901), .Z(N5902) );
  GTECH_OR2 C9626 ( .A(N5898), .B(N5899), .Z(N5900) );
  GTECH_AND2 C9627 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[36]), .Z(N5898) );
  GTECH_AND2 C9628 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[47]), .Z(
        N5899) );
  GTECH_AND2 C9629 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5901) );
  GTECH_AND2 C9630 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[47]), .Z(N5903) );
  GTECH_OR2 C9631 ( .A(N5908), .B(N5909), .Z(add_frac_out[46]) );
  GTECH_OR2 C9632 ( .A(N5906), .B(N5907), .Z(N5908) );
  GTECH_OR2 C9633 ( .A(N5904), .B(N5905), .Z(N5906) );
  GTECH_AND2 C9634 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[35]), .Z(N5904) );
  GTECH_AND2 C9635 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[46]), .Z(
        N5905) );
  GTECH_AND2 C9636 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5907) );
  GTECH_AND2 C9637 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[46]), .Z(N5909) );
  GTECH_OR2 C9638 ( .A(N5914), .B(N5915), .Z(add_frac_out[45]) );
  GTECH_OR2 C9639 ( .A(N5912), .B(N5913), .Z(N5914) );
  GTECH_OR2 C9640 ( .A(N5910), .B(N5911), .Z(N5912) );
  GTECH_AND2 C9641 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[34]), .Z(N5910) );
  GTECH_AND2 C9642 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[45]), .Z(
        N5911) );
  GTECH_AND2 C9643 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5913) );
  GTECH_AND2 C9644 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[45]), .Z(N5915) );
  GTECH_OR2 C9645 ( .A(N5920), .B(N5921), .Z(add_frac_out[44]) );
  GTECH_OR2 C9646 ( .A(N5918), .B(N5919), .Z(N5920) );
  GTECH_OR2 C9647 ( .A(N5916), .B(N5917), .Z(N5918) );
  GTECH_AND2 C9648 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[33]), .Z(N5916) );
  GTECH_AND2 C9649 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[44]), .Z(
        N5917) );
  GTECH_AND2 C9650 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5919) );
  GTECH_AND2 C9651 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[44]), .Z(N5921) );
  GTECH_OR2 C9652 ( .A(N5926), .B(N5927), .Z(add_frac_out[43]) );
  GTECH_OR2 C9653 ( .A(N5924), .B(N5925), .Z(N5926) );
  GTECH_OR2 C9654 ( .A(N5922), .B(N5923), .Z(N5924) );
  GTECH_AND2 C9655 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[32]), .Z(N5922) );
  GTECH_AND2 C9656 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[43]), .Z(
        N5923) );
  GTECH_AND2 C9657 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5925) );
  GTECH_AND2 C9658 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[43]), .Z(N5927) );
  GTECH_OR2 C9659 ( .A(N5932), .B(N5933), .Z(add_frac_out[42]) );
  GTECH_OR2 C9660 ( .A(N5930), .B(N5931), .Z(N5932) );
  GTECH_OR2 C9661 ( .A(N5928), .B(N5929), .Z(N5930) );
  GTECH_AND2 C9662 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[31]), .Z(N5928) );
  GTECH_AND2 C9663 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[42]), .Z(
        N5929) );
  GTECH_AND2 C9664 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5931) );
  GTECH_AND2 C9665 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[42]), .Z(N5933) );
  GTECH_OR2 C9666 ( .A(N5938), .B(N5939), .Z(add_frac_out[41]) );
  GTECH_OR2 C9667 ( .A(N5936), .B(N5937), .Z(N5938) );
  GTECH_OR2 C9668 ( .A(N5934), .B(N5935), .Z(N5936) );
  GTECH_AND2 C9669 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[30]), .Z(N5934) );
  GTECH_AND2 C9670 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[41]), .Z(
        N5935) );
  GTECH_AND2 C9671 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5937) );
  GTECH_AND2 C9672 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[41]), .Z(N5939) );
  GTECH_OR2 C9673 ( .A(N5944), .B(N5945), .Z(add_frac_out[40]) );
  GTECH_OR2 C9674 ( .A(N5942), .B(N5943), .Z(N5944) );
  GTECH_OR2 C9675 ( .A(N5940), .B(N5941), .Z(N5942) );
  GTECH_AND2 C9676 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[29]), .Z(N5940) );
  GTECH_AND2 C9677 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[40]), .Z(
        N5941) );
  GTECH_AND2 C9678 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5943) );
  GTECH_AND2 C9679 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[40]), .Z(N5945) );
  GTECH_OR2 C9680 ( .A(N5950), .B(N5951), .Z(add_frac_out[39]) );
  GTECH_OR2 C9681 ( .A(N5948), .B(N5949), .Z(N5950) );
  GTECH_OR2 C9682 ( .A(N5946), .B(N5947), .Z(N5948) );
  GTECH_AND2 C9683 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[28]), .Z(N5946) );
  GTECH_AND2 C9684 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[39]), .Z(
        N5947) );
  GTECH_AND2 C9685 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5949) );
  GTECH_AND2 C9686 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[39]), .Z(N5951) );
  GTECH_OR2 C9687 ( .A(N5956), .B(N5957), .Z(add_frac_out[38]) );
  GTECH_OR2 C9688 ( .A(N5954), .B(N5955), .Z(N5956) );
  GTECH_OR2 C9689 ( .A(N5952), .B(N5953), .Z(N5954) );
  GTECH_AND2 C9690 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[27]), .Z(N5952) );
  GTECH_AND2 C9691 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[38]), .Z(
        N5953) );
  GTECH_AND2 C9692 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5955) );
  GTECH_AND2 C9693 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[38]), .Z(N5957) );
  GTECH_OR2 C9694 ( .A(N5962), .B(N5963), .Z(add_frac_out[37]) );
  GTECH_OR2 C9695 ( .A(N5960), .B(N5961), .Z(N5962) );
  GTECH_OR2 C9696 ( .A(N5958), .B(N5959), .Z(N5960) );
  GTECH_AND2 C9697 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[26]), .Z(N5958) );
  GTECH_AND2 C9698 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[37]), .Z(
        N5959) );
  GTECH_AND2 C9699 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5961) );
  GTECH_AND2 C9700 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[37]), .Z(N5963) );
  GTECH_OR2 C9701 ( .A(N5968), .B(N5969), .Z(add_frac_out[36]) );
  GTECH_OR2 C9702 ( .A(N5966), .B(N5967), .Z(N5968) );
  GTECH_OR2 C9703 ( .A(N5964), .B(N5965), .Z(N5966) );
  GTECH_AND2 C9704 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[25]), .Z(N5964) );
  GTECH_AND2 C9705 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[36]), .Z(
        N5965) );
  GTECH_AND2 C9706 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5967) );
  GTECH_AND2 C9707 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[36]), .Z(N5969) );
  GTECH_OR2 C9708 ( .A(N5974), .B(N5975), .Z(add_frac_out[35]) );
  GTECH_OR2 C9709 ( .A(N5972), .B(N5973), .Z(N5974) );
  GTECH_OR2 C9710 ( .A(N5970), .B(N5971), .Z(N5972) );
  GTECH_AND2 C9711 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[24]), .Z(N5970) );
  GTECH_AND2 C9712 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[35]), .Z(
        N5971) );
  GTECH_AND2 C9713 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5973) );
  GTECH_AND2 C9714 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[35]), .Z(N5975) );
  GTECH_OR2 C9715 ( .A(N5980), .B(N5981), .Z(add_frac_out[34]) );
  GTECH_OR2 C9716 ( .A(N5978), .B(N5979), .Z(N5980) );
  GTECH_OR2 C9717 ( .A(N5976), .B(N5977), .Z(N5978) );
  GTECH_AND2 C9718 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[23]), .Z(N5976) );
  GTECH_AND2 C9719 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[34]), .Z(
        N5977) );
  GTECH_AND2 C9720 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5979) );
  GTECH_AND2 C9721 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[34]), .Z(N5981) );
  GTECH_OR2 C9722 ( .A(N5986), .B(N5987), .Z(add_frac_out[33]) );
  GTECH_OR2 C9723 ( .A(N5984), .B(N5985), .Z(N5986) );
  GTECH_OR2 C9724 ( .A(N5982), .B(N5983), .Z(N5984) );
  GTECH_AND2 C9725 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[22]), .Z(N5982) );
  GTECH_AND2 C9726 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[33]), .Z(
        N5983) );
  GTECH_AND2 C9727 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5985) );
  GTECH_AND2 C9728 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[33]), .Z(N5987) );
  GTECH_OR2 C9729 ( .A(N5992), .B(N5993), .Z(add_frac_out[32]) );
  GTECH_OR2 C9730 ( .A(N5990), .B(N5991), .Z(N5992) );
  GTECH_OR2 C9731 ( .A(N5988), .B(N5989), .Z(N5990) );
  GTECH_AND2 C9732 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[21]), .Z(N5988) );
  GTECH_AND2 C9733 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[32]), .Z(
        N5989) );
  GTECH_AND2 C9734 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5991) );
  GTECH_AND2 C9735 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[32]), .Z(N5993) );
  GTECH_OR2 C9736 ( .A(N5998), .B(N5999), .Z(add_frac_out[31]) );
  GTECH_OR2 C9737 ( .A(N5996), .B(N5997), .Z(N5998) );
  GTECH_OR2 C9738 ( .A(N5994), .B(N5995), .Z(N5996) );
  GTECH_AND2 C9739 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[20]), .Z(N5994) );
  GTECH_AND2 C9740 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[31]), .Z(
        N5995) );
  GTECH_AND2 C9741 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N5997) );
  GTECH_AND2 C9742 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[31]), .Z(N5999) );
  GTECH_OR2 C9743 ( .A(N6004), .B(N6005), .Z(add_frac_out[30]) );
  GTECH_OR2 C9744 ( .A(N6002), .B(N6003), .Z(N6004) );
  GTECH_OR2 C9745 ( .A(N6000), .B(N6001), .Z(N6002) );
  GTECH_AND2 C9746 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[19]), .Z(N6000) );
  GTECH_AND2 C9747 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[30]), .Z(
        N6001) );
  GTECH_AND2 C9748 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6003) );
  GTECH_AND2 C9749 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[30]), .Z(N6005) );
  GTECH_OR2 C9750 ( .A(N6010), .B(N6011), .Z(add_frac_out[29]) );
  GTECH_OR2 C9751 ( .A(N6008), .B(N6009), .Z(N6010) );
  GTECH_OR2 C9752 ( .A(N6006), .B(N6007), .Z(N6008) );
  GTECH_AND2 C9753 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[18]), .Z(N6006) );
  GTECH_AND2 C9754 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[29]), .Z(
        N6007) );
  GTECH_AND2 C9755 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6009) );
  GTECH_AND2 C9756 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[29]), .Z(N6011) );
  GTECH_OR2 C9757 ( .A(N6016), .B(N6017), .Z(add_frac_out[28]) );
  GTECH_OR2 C9758 ( .A(N6014), .B(N6015), .Z(N6016) );
  GTECH_OR2 C9759 ( .A(N6012), .B(N6013), .Z(N6014) );
  GTECH_AND2 C9760 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[17]), .Z(N6012) );
  GTECH_AND2 C9761 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[28]), .Z(
        N6013) );
  GTECH_AND2 C9762 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6015) );
  GTECH_AND2 C9763 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[28]), .Z(N6017) );
  GTECH_OR2 C9764 ( .A(N6022), .B(N6023), .Z(add_frac_out[27]) );
  GTECH_OR2 C9765 ( .A(N6020), .B(N6021), .Z(N6022) );
  GTECH_OR2 C9766 ( .A(N6018), .B(N6019), .Z(N6020) );
  GTECH_AND2 C9767 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[16]), .Z(N6018) );
  GTECH_AND2 C9768 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[27]), .Z(
        N6019) );
  GTECH_AND2 C9769 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6021) );
  GTECH_AND2 C9770 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[27]), .Z(N6023) );
  GTECH_OR2 C9771 ( .A(N6028), .B(N6029), .Z(add_frac_out[26]) );
  GTECH_OR2 C9772 ( .A(N6026), .B(N6027), .Z(N6028) );
  GTECH_OR2 C9773 ( .A(N6024), .B(N6025), .Z(N6026) );
  GTECH_AND2 C9774 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[15]), .Z(N6024) );
  GTECH_AND2 C9775 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[26]), .Z(
        N6025) );
  GTECH_AND2 C9776 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6027) );
  GTECH_AND2 C9777 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[26]), .Z(N6029) );
  GTECH_OR2 C9778 ( .A(N6034), .B(N6035), .Z(add_frac_out[25]) );
  GTECH_OR2 C9779 ( .A(N6032), .B(N6033), .Z(N6034) );
  GTECH_OR2 C9780 ( .A(N6030), .B(N6031), .Z(N6032) );
  GTECH_AND2 C9781 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[14]), .Z(N6030) );
  GTECH_AND2 C9782 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[25]), .Z(
        N6031) );
  GTECH_AND2 C9783 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6033) );
  GTECH_AND2 C9784 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[25]), .Z(N6035) );
  GTECH_OR2 C9785 ( .A(N6040), .B(N6041), .Z(add_frac_out[24]) );
  GTECH_OR2 C9786 ( .A(N6038), .B(N6039), .Z(N6040) );
  GTECH_OR2 C9787 ( .A(N6036), .B(N6037), .Z(N6038) );
  GTECH_AND2 C9788 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[13]), .Z(N6036) );
  GTECH_AND2 C9789 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[24]), .Z(
        N6037) );
  GTECH_AND2 C9790 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6039) );
  GTECH_AND2 C9791 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[24]), .Z(N6041) );
  GTECH_OR2 C9792 ( .A(N6046), .B(N6047), .Z(add_frac_out[23]) );
  GTECH_OR2 C9793 ( .A(N6044), .B(N6045), .Z(N6046) );
  GTECH_OR2 C9794 ( .A(N6042), .B(N6043), .Z(N6044) );
  GTECH_AND2 C9795 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[12]), .Z(N6042) );
  GTECH_AND2 C9796 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[23]), .Z(
        N6043) );
  GTECH_AND2 C9797 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6045) );
  GTECH_AND2 C9798 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[23]), .Z(N6047) );
  GTECH_OR2 C9799 ( .A(N6052), .B(N6053), .Z(add_frac_out[22]) );
  GTECH_OR2 C9800 ( .A(N6050), .B(N6051), .Z(N6052) );
  GTECH_OR2 C9801 ( .A(N6048), .B(N6049), .Z(N6050) );
  GTECH_AND2 C9802 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[11]), .Z(N6048) );
  GTECH_AND2 C9803 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[22]), .Z(
        N6049) );
  GTECH_AND2 C9804 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6051) );
  GTECH_AND2 C9805 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[22]), .Z(N6053) );
  GTECH_OR2 C9806 ( .A(N6058), .B(N6059), .Z(add_frac_out[21]) );
  GTECH_OR2 C9807 ( .A(N6056), .B(N6057), .Z(N6058) );
  GTECH_OR2 C9808 ( .A(N6054), .B(N6055), .Z(N6056) );
  GTECH_AND2 C9809 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[10]), .Z(N6054) );
  GTECH_AND2 C9810 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[21]), .Z(
        N6055) );
  GTECH_AND2 C9811 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6057) );
  GTECH_AND2 C9812 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[21]), .Z(N6059) );
  GTECH_OR2 C9813 ( .A(N6064), .B(N6065), .Z(add_frac_out[20]) );
  GTECH_OR2 C9814 ( .A(N6062), .B(N6063), .Z(N6064) );
  GTECH_OR2 C9815 ( .A(N6060), .B(N6061), .Z(N6062) );
  GTECH_AND2 C9816 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[9]), .Z(N6060)
         );
  GTECH_AND2 C9817 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[20]), .Z(
        N6061) );
  GTECH_AND2 C9818 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6063) );
  GTECH_AND2 C9819 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[20]), .Z(N6065) );
  GTECH_OR2 C9820 ( .A(N6070), .B(N6071), .Z(add_frac_out[19]) );
  GTECH_OR2 C9821 ( .A(N6068), .B(N6069), .Z(N6070) );
  GTECH_OR2 C9822 ( .A(N6066), .B(N6067), .Z(N6068) );
  GTECH_AND2 C9823 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[8]), .Z(N6066)
         );
  GTECH_AND2 C9824 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[19]), .Z(
        N6067) );
  GTECH_AND2 C9825 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6069) );
  GTECH_AND2 C9826 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[19]), .Z(N6071) );
  GTECH_OR2 C9827 ( .A(N6076), .B(N6077), .Z(add_frac_out[18]) );
  GTECH_OR2 C9828 ( .A(N6074), .B(N6075), .Z(N6076) );
  GTECH_OR2 C9829 ( .A(N6072), .B(N6073), .Z(N6074) );
  GTECH_AND2 C9830 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[7]), .Z(N6072)
         );
  GTECH_AND2 C9831 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[18]), .Z(
        N6073) );
  GTECH_AND2 C9832 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6075) );
  GTECH_AND2 C9833 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[18]), .Z(N6077) );
  GTECH_OR2 C9834 ( .A(N6082), .B(N6083), .Z(add_frac_out[17]) );
  GTECH_OR2 C9835 ( .A(N6080), .B(N6081), .Z(N6082) );
  GTECH_OR2 C9836 ( .A(N6078), .B(N6079), .Z(N6080) );
  GTECH_AND2 C9837 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[6]), .Z(N6078)
         );
  GTECH_AND2 C9838 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[17]), .Z(
        N6079) );
  GTECH_AND2 C9839 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6081) );
  GTECH_AND2 C9840 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[17]), .Z(N6083) );
  GTECH_OR2 C9841 ( .A(N6088), .B(N6089), .Z(add_frac_out[16]) );
  GTECH_OR2 C9842 ( .A(N6086), .B(N6087), .Z(N6088) );
  GTECH_OR2 C9843 ( .A(N6084), .B(N6085), .Z(N6086) );
  GTECH_AND2 C9844 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[5]), .Z(N6084)
         );
  GTECH_AND2 C9845 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[16]), .Z(
        N6085) );
  GTECH_AND2 C9846 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6087) );
  GTECH_AND2 C9847 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[16]), .Z(N6089) );
  GTECH_OR2 C9848 ( .A(N6094), .B(N6095), .Z(add_frac_out[15]) );
  GTECH_OR2 C9849 ( .A(N6092), .B(N6093), .Z(N6094) );
  GTECH_OR2 C9850 ( .A(N6090), .B(N6091), .Z(N6092) );
  GTECH_AND2 C9851 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[4]), .Z(N6090)
         );
  GTECH_AND2 C9852 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[15]), .Z(
        N6091) );
  GTECH_AND2 C9853 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6093) );
  GTECH_AND2 C9854 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[15]), .Z(N6095) );
  GTECH_OR2 C9855 ( .A(N6100), .B(N6101), .Z(add_frac_out[14]) );
  GTECH_OR2 C9856 ( .A(N6098), .B(N6099), .Z(N6100) );
  GTECH_OR2 C9857 ( .A(N6096), .B(N6097), .Z(N6098) );
  GTECH_AND2 C9858 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[3]), .Z(N6096)
         );
  GTECH_AND2 C9859 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[14]), .Z(
        N6097) );
  GTECH_AND2 C9860 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6099) );
  GTECH_AND2 C9861 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[14]), .Z(N6101) );
  GTECH_OR2 C9862 ( .A(N6106), .B(N6107), .Z(add_frac_out[13]) );
  GTECH_OR2 C9863 ( .A(N6104), .B(N6105), .Z(N6106) );
  GTECH_OR2 C9864 ( .A(N6102), .B(N6103), .Z(N6104) );
  GTECH_AND2 C9865 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[2]), .Z(N6102)
         );
  GTECH_AND2 C9866 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[13]), .Z(
        N6103) );
  GTECH_AND2 C9867 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6105) );
  GTECH_AND2 C9868 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[13]), .Z(N6107) );
  GTECH_OR2 C9869 ( .A(N6112), .B(N6113), .Z(add_frac_out[12]) );
  GTECH_OR2 C9870 ( .A(N6110), .B(N6111), .Z(N6112) );
  GTECH_OR2 C9871 ( .A(N6108), .B(N6109), .Z(N6110) );
  GTECH_AND2 C9872 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[1]), .Z(N6108)
         );
  GTECH_AND2 C9873 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[12]), .Z(
        N6109) );
  GTECH_AND2 C9874 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6111) );
  GTECH_AND2 C9875 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[12]), .Z(N6113) );
  GTECH_OR2 C9876 ( .A(N6118), .B(N6119), .Z(add_frac_out[11]) );
  GTECH_OR2 C9877 ( .A(N6116), .B(N6117), .Z(N6118) );
  GTECH_OR2 C9878 ( .A(N6114), .B(N6115), .Z(N6116) );
  GTECH_AND2 C9879 ( .A(a5stg_frac_out_rndadd), .B(a5stg_rndadd[0]), .Z(N6114)
         );
  GTECH_AND2 C9880 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[11]), .Z(
        N6115) );
  GTECH_AND2 C9881 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6117) );
  GTECH_AND2 C9882 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[11]), .Z(N6119) );
  GTECH_OR2 C9883 ( .A(N6122), .B(N6123), .Z(add_frac_out[10]) );
  GTECH_OR2 C9884 ( .A(N6120), .B(N6121), .Z(N6122) );
  GTECH_AND2 C9885 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[10]), .Z(
        N6120) );
  GTECH_AND2 C9886 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6121) );
  GTECH_AND2 C9887 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[10]), .Z(N6123) );
  GTECH_OR2 C9888 ( .A(N6126), .B(N6127), .Z(add_frac_out[9]) );
  GTECH_OR2 C9889 ( .A(N6124), .B(N6125), .Z(N6126) );
  GTECH_AND2 C9890 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[9]), .Z(
        N6124) );
  GTECH_AND2 C9891 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6125) );
  GTECH_AND2 C9892 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[9]), .Z(N6127) );
  GTECH_OR2 C9893 ( .A(N6130), .B(N6131), .Z(add_frac_out[8]) );
  GTECH_OR2 C9894 ( .A(N6128), .B(N6129), .Z(N6130) );
  GTECH_AND2 C9895 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[8]), .Z(
        N6128) );
  GTECH_AND2 C9896 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6129) );
  GTECH_AND2 C9897 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[8]), .Z(N6131) );
  GTECH_OR2 C9898 ( .A(N6134), .B(N6135), .Z(add_frac_out[7]) );
  GTECH_OR2 C9899 ( .A(N6132), .B(N6133), .Z(N6134) );
  GTECH_AND2 C9900 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[7]), .Z(
        N6132) );
  GTECH_AND2 C9901 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6133) );
  GTECH_AND2 C9902 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[7]), .Z(N6135) );
  GTECH_OR2 C9903 ( .A(N6138), .B(N6139), .Z(add_frac_out[6]) );
  GTECH_OR2 C9904 ( .A(N6136), .B(N6137), .Z(N6138) );
  GTECH_AND2 C9905 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[6]), .Z(
        N6136) );
  GTECH_AND2 C9906 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6137) );
  GTECH_AND2 C9907 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[6]), .Z(N6139) );
  GTECH_OR2 C9908 ( .A(N6142), .B(N6143), .Z(add_frac_out[5]) );
  GTECH_OR2 C9909 ( .A(N6140), .B(N6141), .Z(N6142) );
  GTECH_AND2 C9910 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[5]), .Z(
        N6140) );
  GTECH_AND2 C9911 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6141) );
  GTECH_AND2 C9912 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[5]), .Z(N6143) );
  GTECH_OR2 C9913 ( .A(N6146), .B(N6147), .Z(add_frac_out[4]) );
  GTECH_OR2 C9914 ( .A(N6144), .B(N6145), .Z(N6146) );
  GTECH_AND2 C9915 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[4]), .Z(
        N6144) );
  GTECH_AND2 C9916 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6145) );
  GTECH_AND2 C9917 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[4]), .Z(N6147) );
  GTECH_OR2 C9918 ( .A(N6150), .B(N6151), .Z(add_frac_out[3]) );
  GTECH_OR2 C9919 ( .A(N6148), .B(N6149), .Z(N6150) );
  GTECH_AND2 C9920 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[3]), .Z(
        N6148) );
  GTECH_AND2 C9921 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6149) );
  GTECH_AND2 C9922 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[3]), .Z(N6151) );
  GTECH_OR2 C9923 ( .A(N6154), .B(N6155), .Z(add_frac_out[2]) );
  GTECH_OR2 C9924 ( .A(N6152), .B(N6153), .Z(N6154) );
  GTECH_AND2 C9925 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[2]), .Z(
        N6152) );
  GTECH_AND2 C9926 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6153) );
  GTECH_AND2 C9927 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[2]), .Z(N6155) );
  GTECH_OR2 C9928 ( .A(N6158), .B(N6159), .Z(add_frac_out[1]) );
  GTECH_OR2 C9929 ( .A(N6156), .B(N6157), .Z(N6158) );
  GTECH_AND2 C9930 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[1]), .Z(
        N6156) );
  GTECH_AND2 C9931 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6157) );
  GTECH_AND2 C9932 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[1]), .Z(N6159) );
  GTECH_OR2 C9933 ( .A(N6162), .B(N6163), .Z(add_frac_out[0]) );
  GTECH_OR2 C9934 ( .A(N6160), .B(N6161), .Z(N6162) );
  GTECH_AND2 C9935 ( .A(a5stg_frac_out_rnd_frac), .B(a5stg_rnd_frac[0]), .Z(
        N6160) );
  GTECH_AND2 C9936 ( .A(a5stg_in_of), .B(a5stg_to_0), .Z(N6161) );
  GTECH_AND2 C9937 ( .A(a5stg_frac_out_shl), .B(a5stg_shl[0]), .Z(N6163) );
endmodule


module fpu_add ( inq_op, inq_rnd_mode, inq_id, inq_fcc, inq_in1, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, add_dest_rdy, 
        fadd_clken_l, arst_l, grst_l, rclk, add_pipe_active, a1stg_step, 
        a6stg_fadd_in, add_id_out_in, a6stg_fcmpop, add_exc_out, a6stg_dbl_dst, 
        a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, add_sign_out, 
        add_exp_out, add_frac_out, add_cc_out, add_fcc_out, se_add_exp, 
        se_add_frac, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [1:0] inq_fcc;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] add_id_out_in;
  output [4:0] add_exc_out;
  output [10:0] add_exp_out;
  output [63:0] add_frac_out;
  output [1:0] add_cc_out;
  output [1:0] add_fcc_out;
  input inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0,
         inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0,
         inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, add_dest_rdy,
         fadd_clken_l, arst_l, grst_l, rclk, se_add_exp, se_add_frac, si;
  output add_pipe_active, a1stg_step, a6stg_fadd_in, a6stg_fcmpop,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         add_sign_out, so;
  wire   a1stg_in2_neq_in1_frac, a1stg_in2_gt_in1_frac, a1stg_in2_eq_in1_exp,
         a2stg_frac2hi_neq_0, a2stg_frac2lo_neq_0, a3stg_fsdtoix_nx,
         a3stg_fsdtoi_nx, a2stg_frac2_63, add_of_out_cout, a4stg_frac_neq_0,
         a4stg_shl_data_neq_0, a4stg_frac_dbl_nx, a4stg_frac_sng_nx,
         a3stg_denorm, a3stg_denorm_inv, a4stg_denorm_inv, a4stg_round,
         a4stg_rnd_frac_40, a4stg_rnd_frac_39, a4stg_rnd_frac_11,
         a4stg_rnd_frac_10, a4stg_frac_38_0_nx, a4stg_frac_9_0_nx,
         a1stg_denorm_sng_in1, a1stg_denorm_dbl_in1, a1stg_denorm_sng_in2,
         a1stg_denorm_dbl_in2, a1stg_norm_sng_in1, a1stg_norm_dbl_in1,
         a1stg_norm_sng_in2, a1stg_norm_dbl_in2, a1stg_stepa, a1stg_sngop,
         a1stg_intlngop, a1stg_fsdtoix, a1stg_fstod, a1stg_fstoi, a1stg_fstox,
         a1stg_fdtoi, a1stg_fdtox, a1stg_faddsubs, a1stg_faddsubd, a1stg_fdtos,
         a2stg_faddsubop, a2stg_fsdtoix_fdtos, a2stg_fitos, a2stg_fitod,
         a2stg_fxtos, a2stg_fxtod, a3stg_faddsubop, a4stg_dblop, a6stg_step,
         a3stg_sub_in, a4stg_in_of, a2stg_frac1_in_frac1, a2stg_frac1_in_frac2,
         a1stg_2nan_in_inv, a1stg_faddsubop_inv, a2stg_frac1_in_qnan,
         a2stg_frac1_in_nv, a2stg_frac1_in_nv_dbl, a2stg_frac2_in_frac1,
         a2stg_frac2_in_qnan, a2stg_shr_cnt_5_inv_in, a2stg_shr_frac2_shr_int,
         a2stg_shr_frac2_shr_dbl, a2stg_shr_frac2_shr_sng, a2stg_shr_frac2_max,
         a2stg_sub_step, a2stg_fracadd_frac2_inv_in,
         a2stg_fracadd_frac2_inv_shr1_in, a2stg_fracadd_frac2,
         a2stg_fracadd_cin_in, a3stg_exp_7ff, a3stg_exp_ff, a3stg_exp_add,
         a2stg_expdec_neq_0, a3stg_exp10_0_eq0, a3stg_exp10_1_eq0,
         a3stg_fdtos_inv, a4stg_fixtos_fxtod_inv, a4stg_rnd_frac_add_inv,
         a4stg_rnd_sng, a4stg_rnd_dbl, add_frac_out_rndadd,
         add_frac_out_rnd_frac, add_frac_out_shl, a4stg_to_0,
         add_exp_out_expinc, add_exp_out_exp, add_exp_out_exp1,
         add_exp_out_expadd, a4stg_to_0_inv, scan_out_fpu_add_ctl,
         a3stg_inc_exp_inv, a3stg_same_exp_inv, a3stg_dec_exp_inv,
         a4stg_rndadd_cout, a1stg_expadd3_11, scan_out_fpu_add_exp_dp;
  wire   [11:0] a1stg_expadd1_11_0;
  wire   [12:0] a2stg_expadd;
  wire   [11:0] a2stg_exp;
  wire   [11:0] a4stg_exp_11_0;
  wire   [5:0] a1stg_expadd2_5_0;
  wire   [10:0] a1stg_expadd4_inv;
  wire   [10:0] a3stg_exp_10_0;
  wire   [5:0] a3stg_lead0;
  wire   [1:0] a3stg_faddsubopa;
  wire   [5:0] a2stg_shr_cnt_in;
  wire   [9:0] a4stg_shl_cnt_in;
  wire   [5:0] a4stg_shl_cnt;

  fpu_add_ctl fpu_add_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_63(inq_in1[63]), .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(inq_in1_exp_neq_ffs), 
        .inq_in2_51(inq_in2[51]), .inq_in2_54(inq_in2[54]), .inq_in2_63(
        inq_in2[63]), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0), .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(
        inq_op), .inq_rnd_mode(inq_rnd_mode), .inq_id(inq_id), .inq_fcc(
        inq_fcc), .inq_add(inq_add), .add_dest_rdy(add_dest_rdy), 
        .a1stg_in2_neq_in1_frac(a1stg_in2_neq_in1_frac), 
        .a1stg_in2_gt_in1_frac(a1stg_in2_gt_in1_frac), .a1stg_in2_eq_in1_exp(
        a1stg_in2_eq_in1_exp), .a1stg_expadd1(a1stg_expadd1_11_0), 
        .a2stg_expadd(a2stg_expadd[11:0]), .a2stg_frac2hi_neq_0(
        a2stg_frac2hi_neq_0), .a2stg_frac2lo_neq_0(a2stg_frac2lo_neq_0), 
        .a2stg_exp(a2stg_exp), .a3stg_fsdtoix_nx(a3stg_fsdtoix_nx), 
        .a3stg_fsdtoi_nx(a3stg_fsdtoi_nx), .a2stg_frac2_63(a2stg_frac2_63), 
        .a4stg_exp(a4stg_exp_11_0), .add_of_out_cout(add_of_out_cout), 
        .a4stg_frac_neq_0(a4stg_frac_neq_0), .a4stg_shl_data_neq_0(
        a4stg_shl_data_neq_0), .a4stg_frac_dbl_nx(a4stg_frac_dbl_nx), 
        .a4stg_frac_sng_nx(a4stg_frac_sng_nx), .a1stg_expadd2(
        a1stg_expadd2_5_0), .a1stg_expadd4_inv(a1stg_expadd4_inv), 
        .a3stg_denorm(a3stg_denorm), .a3stg_denorm_inv(a3stg_denorm_inv), 
        .a4stg_denorm_inv(a4stg_denorm_inv), .a3stg_exp(a3stg_exp_10_0), 
        .a4stg_round(a4stg_round), .a3stg_lead0(a3stg_lead0), 
        .a4stg_rnd_frac_40(a4stg_rnd_frac_40), .a4stg_rnd_frac_39(
        a4stg_rnd_frac_39), .a4stg_rnd_frac_11(a4stg_rnd_frac_11), 
        .a4stg_rnd_frac_10(a4stg_rnd_frac_10), .a4stg_frac_38_0_nx(
        a4stg_frac_38_0_nx), .a4stg_frac_9_0_nx(a4stg_frac_9_0_nx), .arst_l(
        arst_l), .grst_l(grst_l), .rclk(rclk), .add_pipe_active(
        add_pipe_active), .a1stg_denorm_sng_in1(a1stg_denorm_sng_in1), 
        .a1stg_denorm_dbl_in1(a1stg_denorm_dbl_in1), .a1stg_denorm_sng_in2(
        a1stg_denorm_sng_in2), .a1stg_denorm_dbl_in2(a1stg_denorm_dbl_in2), 
        .a1stg_norm_sng_in1(a1stg_norm_sng_in1), .a1stg_norm_dbl_in1(
        a1stg_norm_dbl_in1), .a1stg_norm_sng_in2(a1stg_norm_sng_in2), 
        .a1stg_norm_dbl_in2(a1stg_norm_dbl_in2), .a1stg_step(a1stg_step), 
        .a1stg_stepa(a1stg_stepa), .a1stg_sngop(a1stg_sngop), .a1stg_intlngop(
        a1stg_intlngop), .a1stg_fsdtoix(a1stg_fsdtoix), .a1stg_fstod(
        a1stg_fstod), .a1stg_fstoi(a1stg_fstoi), .a1stg_fstox(a1stg_fstox), 
        .a1stg_fdtoi(a1stg_fdtoi), .a1stg_fdtox(a1stg_fdtox), .a1stg_faddsubs(
        a1stg_faddsubs), .a1stg_faddsubd(a1stg_faddsubd), .a1stg_fdtos(
        a1stg_fdtos), .a2stg_faddsubop(a2stg_faddsubop), .a2stg_fsdtoix_fdtos(
        a2stg_fsdtoix_fdtos), .a2stg_fitos(a2stg_fitos), .a2stg_fitod(
        a2stg_fitod), .a2stg_fxtos(a2stg_fxtos), .a2stg_fxtod(a2stg_fxtod), 
        .a3stg_faddsubop(a3stg_faddsubop), .a3stg_faddsubopa(a3stg_faddsubopa), 
        .a4stg_dblop(a4stg_dblop), .a6stg_fadd_in(a6stg_fadd_in), 
        .add_id_out_in(add_id_out_in), .add_fcc_out(add_fcc_out), 
        .a6stg_dbl_dst(a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), 
        .a6stg_long_dst(a6stg_long_dst), .a6stg_int_dst(a6stg_int_dst), 
        .a6stg_fcmpop(a6stg_fcmpop), .a6stg_step(a6stg_step), .a3stg_sub_in(
        a3stg_sub_in), .add_sign_out(add_sign_out), .add_cc_out(add_cc_out), 
        .a4stg_in_of(a4stg_in_of), .add_exc_out(add_exc_out), 
        .a2stg_frac1_in_frac1(a2stg_frac1_in_frac1), .a2stg_frac1_in_frac2(
        a2stg_frac1_in_frac2), .a1stg_2nan_in_inv(a1stg_2nan_in_inv), 
        .a1stg_faddsubop_inv(a1stg_faddsubop_inv), .a2stg_frac1_in_qnan(
        a2stg_frac1_in_qnan), .a2stg_frac1_in_nv(a2stg_frac1_in_nv), 
        .a2stg_frac1_in_nv_dbl(a2stg_frac1_in_nv_dbl), .a2stg_frac2_in_frac1(
        a2stg_frac2_in_frac1), .a2stg_frac2_in_qnan(a2stg_frac2_in_qnan), 
        .a2stg_shr_cnt_in(a2stg_shr_cnt_in), .a2stg_shr_cnt_5_inv_in(
        a2stg_shr_cnt_5_inv_in), .a2stg_shr_frac2_shr_int(
        a2stg_shr_frac2_shr_int), .a2stg_shr_frac2_shr_dbl(
        a2stg_shr_frac2_shr_dbl), .a2stg_shr_frac2_shr_sng(
        a2stg_shr_frac2_shr_sng), .a2stg_shr_frac2_max(a2stg_shr_frac2_max), 
        .a2stg_sub_step(a2stg_sub_step), .a2stg_fracadd_frac2_inv_in(
        a2stg_fracadd_frac2_inv_in), .a2stg_fracadd_frac2_inv_shr1_in(
        a2stg_fracadd_frac2_inv_shr1_in), .a2stg_fracadd_frac2(
        a2stg_fracadd_frac2), .a2stg_fracadd_cin_in(a2stg_fracadd_cin_in), 
        .a3stg_exp_7ff(a3stg_exp_7ff), .a3stg_exp_ff(a3stg_exp_ff), 
        .a3stg_exp_add(a3stg_exp_add), .a2stg_expdec_neq_0(a2stg_expdec_neq_0), 
        .a3stg_exp10_0_eq0(a3stg_exp10_0_eq0), .a3stg_exp10_1_eq0(
        a3stg_exp10_1_eq0), .a3stg_fdtos_inv(a3stg_fdtos_inv), 
        .a4stg_fixtos_fxtod_inv(a4stg_fixtos_fxtod_inv), 
        .a4stg_rnd_frac_add_inv(a4stg_rnd_frac_add_inv), .a4stg_shl_cnt_in(
        a4stg_shl_cnt_in), .a4stg_rnd_sng(a4stg_rnd_sng), .a4stg_rnd_dbl(
        a4stg_rnd_dbl), .add_frac_out_rndadd(add_frac_out_rndadd), 
        .add_frac_out_rnd_frac(add_frac_out_rnd_frac), .add_frac_out_shl(
        add_frac_out_shl), .a4stg_to_0(a4stg_to_0), .add_exp_out_expinc(
        add_exp_out_expinc), .add_exp_out_exp(add_exp_out_exp), 
        .add_exp_out_exp1(add_exp_out_exp1), .add_exp_out_expadd(
        add_exp_out_expadd), .a4stg_to_0_inv(a4stg_to_0_inv), .se(se_add_exp), 
        .si(si), .so(scan_out_fpu_add_ctl) );
  fpu_add_exp_dp fpu_add_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .inq_op(inq_op[1:0]), .inq_op_7(inq_op[7]), 
        .a1stg_step(a1stg_stepa), .a1stg_faddsubd(a1stg_faddsubd), 
        .a1stg_faddsubs(a1stg_faddsubs), .a1stg_fsdtoix(a1stg_fsdtoix), 
        .a6stg_step(a6stg_step), .a1stg_fstod(a1stg_fstod), .a1stg_fdtos(
        a1stg_fdtos), .a1stg_fstoi(a1stg_fstoi), .a1stg_fstox(a1stg_fstox), 
        .a1stg_fdtoi(a1stg_fdtoi), .a1stg_fdtox(a1stg_fdtox), 
        .a2stg_fsdtoix_fdtos(a2stg_fsdtoix_fdtos), .a2stg_faddsubop(
        a2stg_faddsubop), .a2stg_fitos(a2stg_fitos), .a2stg_fitod(a2stg_fitod), 
        .a2stg_fxtos(a2stg_fxtos), .a2stg_fxtod(a2stg_fxtod), .a3stg_exp_7ff(
        a3stg_exp_7ff), .a3stg_exp_ff(a3stg_exp_ff), .a3stg_exp_add(
        a3stg_exp_add), .a3stg_inc_exp_inv(a3stg_inc_exp_inv), 
        .a3stg_same_exp_inv(a3stg_same_exp_inv), .a3stg_dec_exp_inv(
        a3stg_dec_exp_inv), .a3stg_faddsubop(a3stg_faddsubop), 
        .a3stg_fdtos_inv(a3stg_fdtos_inv), .a4stg_fixtos_fxtod_inv(
        a4stg_fixtos_fxtod_inv), .a4stg_shl_cnt(a4stg_shl_cnt), 
        .a4stg_denorm_inv(a4stg_denorm_inv), .a4stg_rndadd_cout(
        a4stg_rndadd_cout), .add_exp_out_expinc(add_exp_out_expinc), 
        .add_exp_out_exp(add_exp_out_exp), .add_exp_out_exp1(add_exp_out_exp1), 
        .a4stg_in_of(a4stg_in_of), .add_exp_out_expadd(add_exp_out_expadd), 
        .a4stg_dblop(a4stg_dblop), .a4stg_to_0_inv(a4stg_to_0_inv), 
        .fadd_clken_l(fadd_clken_l), .rclk(rclk), .a1stg_expadd3_11(
        a1stg_expadd3_11), .a1stg_expadd1_11_0(a1stg_expadd1_11_0), 
        .a1stg_expadd4_inv(a1stg_expadd4_inv), .a1stg_expadd2_5_0(
        a1stg_expadd2_5_0), .a2stg_exp(a2stg_exp), .a2stg_expadd(a2stg_expadd), 
        .a3stg_exp_10_0(a3stg_exp_10_0), .a4stg_exp_11_0(a4stg_exp_11_0), 
        .add_exp_out(add_exp_out), .se(se_add_exp), .si(scan_out_fpu_add_ctl), 
        .so(scan_out_fpu_add_exp_dp) );
  fpu_add_frac_dp fpu_add_frac_dp ( .inq_in1(inq_in1[62:0]), .inq_in2(inq_in2), 
        .a1stg_step(a1stg_stepa), .a1stg_sngop(a1stg_sngop), 
        .a1stg_expadd3_11(a1stg_expadd3_11), .a1stg_norm_dbl_in1(
        a1stg_norm_dbl_in1), .a1stg_denorm_dbl_in1(a1stg_denorm_dbl_in1), 
        .a1stg_norm_sng_in1(a1stg_norm_sng_in1), .a1stg_denorm_sng_in1(
        a1stg_denorm_sng_in1), .a1stg_norm_dbl_in2(a1stg_norm_dbl_in2), 
        .a1stg_denorm_dbl_in2(a1stg_denorm_dbl_in2), .a1stg_norm_sng_in2(
        a1stg_norm_sng_in2), .a1stg_denorm_sng_in2(a1stg_denorm_sng_in2), 
        .a1stg_intlngop(a1stg_intlngop), .a2stg_frac1_in_frac1(
        a2stg_frac1_in_frac1), .a2stg_frac1_in_frac2(a2stg_frac1_in_frac2), 
        .a1stg_2nan_in_inv(a1stg_2nan_in_inv), .a1stg_faddsubop_inv(
        a1stg_faddsubop_inv), .a2stg_frac1_in_qnan(a2stg_frac1_in_qnan), 
        .a2stg_frac1_in_nv(a2stg_frac1_in_nv), .a2stg_frac1_in_nv_dbl(
        a2stg_frac1_in_nv_dbl), .a6stg_step(a6stg_step), 
        .a2stg_frac2_in_frac1(a2stg_frac2_in_frac1), .a2stg_frac2_in_qnan(
        a2stg_frac2_in_qnan), .a2stg_shr_cnt_in(a2stg_shr_cnt_in), 
        .a2stg_shr_cnt_5_inv_in(a2stg_shr_cnt_5_inv_in), 
        .a2stg_shr_frac2_shr_int(a2stg_shr_frac2_shr_int), 
        .a2stg_shr_frac2_shr_dbl(a2stg_shr_frac2_shr_dbl), 
        .a2stg_shr_frac2_shr_sng(a2stg_shr_frac2_shr_sng), 
        .a2stg_shr_frac2_max(a2stg_shr_frac2_max), .a2stg_expadd_11(
        a2stg_expadd[12]), .a2stg_sub_step(a2stg_sub_step), 
        .a2stg_fracadd_frac2_inv_in(a2stg_fracadd_frac2_inv_in), 
        .a2stg_fracadd_frac2_inv_shr1_in(a2stg_fracadd_frac2_inv_shr1_in), 
        .a2stg_fracadd_frac2(a2stg_fracadd_frac2), .a2stg_fracadd_cin_in(
        a2stg_fracadd_cin_in), .a2stg_exp(a2stg_exp[5:0]), 
        .a2stg_expdec_neq_0(a2stg_expdec_neq_0), .a3stg_faddsubopa(
        a3stg_faddsubopa), .a3stg_sub_in(a3stg_sub_in), .a3stg_exp10_0_eq0(
        a3stg_exp10_0_eq0), .a3stg_exp10_1_eq0(a3stg_exp10_1_eq0), 
        .a3stg_exp_0(a3stg_exp_10_0[0]), .a4stg_rnd_frac_add_inv(
        a4stg_rnd_frac_add_inv), .a3stg_fdtos_inv(a3stg_fdtos_inv), 
        .a4stg_fixtos_fxtod_inv(a4stg_fixtos_fxtod_inv), .a4stg_rnd_sng(
        a4stg_rnd_sng), .a4stg_rnd_dbl(a4stg_rnd_dbl), .a4stg_shl_cnt_in(
        a4stg_shl_cnt_in), .add_frac_out_rndadd(add_frac_out_rndadd), 
        .add_frac_out_rnd_frac(add_frac_out_rnd_frac), .a4stg_in_of(
        a4stg_in_of), .add_frac_out_shl(add_frac_out_shl), .a4stg_to_0(
        a4stg_to_0), .fadd_clken_l(fadd_clken_l), .rclk(rclk), 
        .a1stg_in2_neq_in1_frac(a1stg_in2_neq_in1_frac), 
        .a1stg_in2_gt_in1_frac(a1stg_in2_gt_in1_frac), .a1stg_in2_eq_in1_exp(
        a1stg_in2_eq_in1_exp), .a2stg_frac2_63(a2stg_frac2_63), 
        .a2stg_frac2hi_neq_0(a2stg_frac2hi_neq_0), .a2stg_frac2lo_neq_0(
        a2stg_frac2lo_neq_0), .a3stg_fsdtoix_nx(a3stg_fsdtoix_nx), 
        .a3stg_fsdtoi_nx(a3stg_fsdtoi_nx), .a3stg_denorm(a3stg_denorm), 
        .a3stg_denorm_inv(a3stg_denorm_inv), .a3stg_lead0(a3stg_lead0), 
        .a4stg_round(a4stg_round), .a4stg_shl_cnt(a4stg_shl_cnt), 
        .a4stg_denorm_inv(a4stg_denorm_inv), .a3stg_inc_exp_inv(
        a3stg_inc_exp_inv), .a3stg_same_exp_inv(a3stg_same_exp_inv), 
        .a3stg_dec_exp_inv(a3stg_dec_exp_inv), .a4stg_rnd_frac_40(
        a4stg_rnd_frac_40), .a4stg_rnd_frac_39(a4stg_rnd_frac_39), 
        .a4stg_rnd_frac_11(a4stg_rnd_frac_11), .a4stg_rnd_frac_10(
        a4stg_rnd_frac_10), .a4stg_rndadd_cout(a4stg_rndadd_cout), 
        .a4stg_frac_9_0_nx(a4stg_frac_9_0_nx), .a4stg_frac_dbl_nx(
        a4stg_frac_dbl_nx), .a4stg_frac_38_0_nx(a4stg_frac_38_0_nx), 
        .a4stg_frac_sng_nx(a4stg_frac_sng_nx), .a4stg_frac_neq_0(
        a4stg_frac_neq_0), .a4stg_shl_data_neq_0(a4stg_shl_data_neq_0), 
        .add_of_out_cout(add_of_out_cout), .add_frac_out(add_frac_out), .se(
        se_add_frac), .si(scan_out_fpu_add_exp_dp), .so(so) );
endmodule


module dffre_SIZE5 ( din, rst, en, clk, q, se, si, so );
  input [4:0] din;
  output [4:0] q;
  input [4:0] si;
  output [4:0] so;
  input rst, en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19;
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N19) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N19) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N19) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N19) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N19) );
  SELECT_OP C47 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(din), 
        .CONTROL1(N0), .CONTROL2(N17), .Z({N10, N9, N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  SELECT_OP C48 ( .DATA1(si), .DATA2({N10, N9, N8, N7, N6}), .CONTROL1(N1), 
        .CONTROL2(N2), .Z({N15, N14, N13, N12, N11}) );
  GTECH_BUF B_1 ( .A(se), .Z(N1) );
  GTECH_BUF B_2 ( .A(N3), .Z(N2) );
  GTECH_NOT I_0 ( .A(se), .Z(N3) );
  GTECH_OR2 C56 ( .A(en), .B(rst), .Z(N4) );
  GTECH_NOT I_1 ( .A(N4), .Z(N5) );
  GTECH_NOT I_2 ( .A(rst), .Z(N16) );
  GTECH_AND2 C59 ( .A(en), .B(N16), .Z(N17) );
  GTECH_AND2 C60 ( .A(N5), .B(N3), .Z(N18) );
  GTECH_NOT I_3 ( .A(N18), .Z(N19) );
endmodule


module dffe_SIZE6 ( din, en, clk, q, se, si, so );
  input [5:0] din;
  output [5:0] q;
  input [5:0] si;
  output [5:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11;
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N11) );
  SELECT_OP C39 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C47 ( .A(N3), .B(N2), .Z(N10) );
  GTECH_NOT I_2 ( .A(N10), .Z(N11) );
endmodule


module dffe_SIZE7 ( din, en, clk, q, se, si, so );
  input [6:0] din;
  output [6:0] q;
  input [6:0] si;
  output [6:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12;
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N12) );
  SELECT_OP C43 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C51 ( .A(N3), .B(N2), .Z(N11) );
  GTECH_NOT I_2 ( .A(N11), .Z(N12) );
endmodule


module fpu_mul_ctl ( inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, inq_op, inq_mul, inq_rnd_mode, inq_id, inq_in1_63, 
        inq_in2_63, mul_dest_rdy, mul_dest_rdya, m5stg_exp, m5stg_fracadd_cout, 
        m5stg_frac_neq_0, m5stg_frac_dbl_nx, m5stg_frac_sng_nx, m1stg_ld0_1, 
        m1stg_ld0_2, m3stg_exp, m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv, 
        m3stg_ld0_inv, m4stg_exp, m4stg_frac_105, m5stg_frac, arst_l, grst_l, 
        rclk, mul_pipe_active, m1stg_snan_sng_in1, m1stg_snan_dbl_in1, 
        m1stg_snan_sng_in2, m1stg_snan_dbl_in2, m1stg_step, m1stg_sngop, 
        m1stg_dblop, m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld, m2stg_fmuls, 
        m2stg_fmuld, m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda, 
        m6stg_fmul_in, m6stg_id_in, m6stg_fmul_dbl_dst, m6stg_fmuls, 
        m6stg_step, mul_sign_out, m5stg_in_of, mul_exc_out, 
        m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm, m2stg_frac1_sng_norm, 
        m2stg_frac1_sng_dnrm, m2stg_frac1_inf, m2stg_frac2_dbl_norm, 
        m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, m2stg_frac2_sng_dnrm, 
        m2stg_frac2_inf, m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, 
        m2stg_exp_expadd, m2stg_exp_0bff, m2stg_exp_017f, m2stg_exp_04ff, 
        m2stg_exp_zero, m3bstg_ld0_inv, m4stg_sh_cnt_in, m4stg_inc_exp_54, 
        m4stg_inc_exp_55, m4stg_inc_exp_105, m4stg_left_shift_step, 
        m4stg_right_shift_step, m5stg_to_0, m5stg_to_0_inv, 
        mul_frac_out_fracadd, mul_frac_out_frac, mul_exp_out_exp_plus1, 
        mul_exp_out_exp, mula_rst_l, se, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [12:0] m5stg_exp;
  input [5:0] m1stg_ld0_1;
  input [5:0] m1stg_ld0_2;
  input [12:0] m3stg_exp;
  input [5:0] m3stg_ld0_inv;
  input [12:0] m4stg_exp;
  input [32:0] m5stg_frac;
  output [9:0] m6stg_id_in;
  output [4:0] mul_exc_out;
  output [6:0] m3bstg_ld0_inv;
  output [5:0] m4stg_sh_cnt_in;
  input inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_mul,
         inq_in1_63, inq_in2_63, mul_dest_rdy, mul_dest_rdya,
         m5stg_fracadd_cout, m5stg_frac_neq_0, m5stg_frac_dbl_nx,
         m5stg_frac_sng_nx, m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv,
         m4stg_frac_105, arst_l, grst_l, rclk, se, si;
  output mul_pipe_active, m1stg_snan_sng_in1, m1stg_snan_dbl_in1,
         m1stg_snan_sng_in2, m1stg_snan_dbl_in2, m1stg_step, m1stg_sngop,
         m1stg_dblop, m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld, m2stg_fmuls,
         m2stg_fmuld, m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda,
         m6stg_fmul_in, m6stg_fmul_dbl_dst, m6stg_fmuls, m6stg_step,
         mul_sign_out, m5stg_in_of, m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm,
         m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, m2stg_frac1_inf,
         m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm,
         m2stg_frac2_sng_dnrm, m2stg_frac2_inf, m1stg_inf_zero_in,
         m1stg_inf_zero_in_dbl, m2stg_exp_expadd, m2stg_exp_0bff,
         m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero, m4stg_inc_exp_54,
         m4stg_inc_exp_55, m4stg_inc_exp_105, m4stg_left_shift_step,
         m4stg_right_shift_step, m5stg_to_0, m5stg_to_0_inv,
         mul_frac_out_fracadd, mul_frac_out_frac, mul_exp_out_exp_plus1,
         mul_exp_out_exp, mula_rst_l, so;
  wire   mul_exc_out_0, reset, mul_frac_in1_51, mul_frac_in1_54,
         mul_frac_in1_53_0_neq_0, mul_frac_in1_50_0_neq_0,
         mul_frac_in1_53_32_neq_0, mul_exp_in1_exp_eq_0,
         mul_exp_in1_exp_neq_ffs, mul_frac_in2_51, mul_frac_in2_54,
         mul_frac_in2_53_0_neq_0, mul_frac_in2_50_0_neq_0,
         mul_frac_in2_53_32_neq_0, mul_exp_in2_exp_eq_0,
         mul_exp_in2_exp_neq_ffs, m1stg_denorm_sng_in1, m1stg_denorm_dbl_in1,
         m1stg_denorm_sng_in2, m1stg_denorm_dbl_in2, m1stg_denorm_in1,
         m1stg_denorm_in2, m1stg_norm_sng_in1, m1stg_norm_dbl_in1,
         m1stg_norm_sng_in2, m1stg_norm_dbl_in2, m1stg_qnan_sng_in1,
         m1stg_qnan_dbl_in1, m1stg_qnan_sng_in2, m1stg_qnan_dbl_in2,
         m1stg_snan_in1, m1stg_snan_in2, m1stg_qnan_in1, m1stg_qnan_in2,
         m2stg_snan_in1, m2stg_snan_in2, m2stg_qnan_in1, m2stg_qnan_in2,
         m1stg_nan_sng_in1, m1stg_nan_dbl_in1, m1stg_nan_sng_in2,
         m1stg_nan_dbl_in2, m1stg_nan_in1, m1stg_nan_in2, m2stg_nan_in2,
         m1stg_inf_sng_in1, m1stg_inf_dbl_in1, m1stg_inf_sng_in2,
         m1stg_inf_dbl_in2, m1stg_inf_in1, m1stg_inf_in2, m1stg_inf_in,
         m2stg_inf_in1, m2stg_inf_in2, m2stg_inf_in, m1stg_infnan_sng_in1,
         m1stg_infnan_dbl_in1, m1stg_infnan_sng_in2, m1stg_infnan_dbl_in2,
         m1stg_infnan_in1, m1stg_infnan_in2, m1stg_infnan_in, m1stg_zero_in1,
         m1stg_zero_in2, m1stg_zero_in, m2stg_zero_in1, m2stg_zero_in2,
         m2stg_zero_in, m6stg_stepa, m1stg_mul, N0, N1, m1stg_mul_in,
         m1stg_dblop_inv_in, N2, m6stg_hold, m6stg_holda, mul_pipe_active_in,
         m1stg_sign1, m1stg_sign2, m2stg_sign1, m2stg_sign2, m1stg_of_mask,
         m2stg_of_mask, N3, m2stg_sign, m3astg_sign, m2stg_nv, m3astg_nv,
         m3astg_of_mask, m3bstg_sign, m3bstg_nv, m3bstg_of_mask, m3stg_sign,
         m3stg_nv, m3stg_of_mask, m4stg_sign, m4stg_nv, m4stg_of_mask,
         m5stg_sign, m5stg_nv, m5stg_of_mask, N4, m5stg_rndup,
         mul_of_out_tmp1_in, mul_of_out_tmp1, mul_of_out_tmp2, mul_of_out_cout,
         mul_uf_out_in, mul_nx_out_in, mul_nx_out, N5, m4stg_expadd_eq_0,
         m3stg_exp_lte_0, m4stg_right_shift_in, m4stg_right_shift,
         m3stg_exp_lt_neg57, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, net14450,
         net14451, net14452, net14453, net14454, net14455, net14456, net14457,
         net14458, net14459, net14460, net14461, net14462, net14463, net14464,
         net14465, net14466, net14467, net14468, net14469, net14470, net14471,
         net14472, net14473, net14474, net14475, net14476, net14477, net14478,
         net14479, net14480, net14481, net14482, net14483, net14484, net14485,
         net14486, net14487, net14488, net14489, net14490, net14491, net14492,
         net14493, net14494, net14495, net14496, net14497, net14498, net14499,
         net14500, net14501, net14502, net14503, net14504, net14505, net14506,
         net14507, net14508, net14509, net14510, net14511, net14512, net14513,
         net14514, net14515, net14516, net14517, net14518, net14519, net14520,
         net14521, net14522, net14523, net14524, net14525, net14526, net14527,
         net14528, net14529, net14530, net14531, net14532, net14533, net14534,
         net14535, net14536, net14537, net14538, net14539, net14540, net14541,
         net14542, net14543, net14544, net14545, net14546, net14547, net14548,
         net14549, net14550, net14551, net14552, net14553, net14554, net14555,
         net14556, net14557, net14558, net14559, net14560, net14561, net14562,
         net14563, net14564, net14565, net14566, net14567, net14568, net14569,
         net14570, net14571, net14572, net14573, net14574, net14575, net14576,
         net14577, net14578, net14579, net14580, net14581, net14582, net14583,
         net14584, net14585, net14586, net14587, net14588, net14589, net14590,
         net14591, net14592, net14593, net14594, net14595, net14596, net14597,
         net14598, net14599, net14600, net14601, net14602, net14603, net14604,
         net14605, net14606, net14607, net14608, net14609, net14610, net14611,
         net14612, net14613, net14614, net14615, net14616, net14617, net14618,
         net14619, net14620, net14621, net14622, net14623, net14624, net14625,
         net14626, net14627, net14628, net14629, net14630, net14631, net14632,
         net14633, net14634, net14635, net14636, net14637, net14638, net14639,
         net14640;
  wire   [3:0] m1stg_sngopa;
  wire   [3:0] m1stg_dblopa;
  wire   [7:0] m1stg_op;
  wire   [7:0] m1stg_op_in;
  wire   [1:0] m1stg_rnd_mode;
  wire   [4:0] m1stg_id;
  wire   [3:3] m1stg_opdec;
  wire   [4:3] m2stg_opdec;
  wire   [1:0] m2stg_rnd_mode;
  wire   [4:0] m2stg_id;
  wire   [4:1] m3astg_opdec;
  wire   [1:0] m3astg_rnd_mode;
  wire   [4:0] m3astg_id;
  wire   [4:1] m3bstg_opdec;
  wire   [1:0] m3bstg_rnd_mode;
  wire   [4:0] m3bstg_id;
  wire   [4:1] m3stg_opdec;
  wire   [1:0] m3stg_rnd_mode;
  wire   [4:0] m3stg_id;
  wire   [4:1] m4stg_opdec;
  wire   [1:0] m4stg_rnd_mode;
  wire   [4:0] m4stg_id;
  wire   [4:3] m5stg_opdec;
  wire   [1:0] m5stg_rnd_mode;
  wire   [4:0] m5stg_id;
  wire   [4:4] m6stg_opdec;
  wire   [9:0] m6stg_id;
  wire   [5:0] m2stg_ld0_1_in;
  wire   [5:0] m2stg_ld0_1;
  wire   [5:0] m2stg_ld0_2_in;
  wire   [5:0] m2stg_ld0_2;
  wire   [6:0] m2stg_ld0;
  wire   [6:0] m2stg_ld0_inv;
  wire   [6:0] m3astg_ld0_inv;
  wire   [5:0] m3stg_exp_minus1;
  wire   [5:0] m3stg_exp_inv_plus2;
  assign mul_exc_out[1] = 1'b0;
  assign mul_exc_out[0] = mul_exc_out_0;
  assign m1stg_fsmuld = N62;

  dffrl_async_SIZE1 dffrl_mul_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(mula_rst_l), .se(se), .si(net14640) );
  dffe_SIZE1 i_mul_frac_in1_51 ( .din(inq_in1_51), .en(m6stg_step), .clk(rclk), 
        .q(mul_frac_in1_51), .se(se), .si(net14639) );
  dffe_SIZE1 i_mul_frac_in1_54 ( .din(inq_in1_54), .en(m6stg_step), .clk(rclk), 
        .q(mul_frac_in1_54), .se(se), .si(net14638) );
  dffe_SIZE1 i_mul_frac_in1_53_0_neq_0 ( .din(inq_in1_53_0_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in1_53_0_neq_0), .se(se), .si(
        net14637) );
  dffe_SIZE1 i_mul_frac_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in1_50_0_neq_0), .se(se), .si(
        net14636) );
  dffe_SIZE1 i_mul_frac_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in1_53_32_neq_0), .se(se), .si(
        net14635) );
  dffe_SIZE1 i_mul_exp_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(m6stg_step), 
        .clk(rclk), .q(mul_exp_in1_exp_eq_0), .se(se), .si(net14634) );
  dffe_SIZE1 i_mul_exp_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        m6stg_step), .clk(rclk), .q(mul_exp_in1_exp_neq_ffs), .se(se), .si(
        net14633) );
  dffe_SIZE1 i_mul_frac_in2_51 ( .din(inq_in2_51), .en(m6stg_step), .clk(rclk), 
        .q(mul_frac_in2_51), .se(se), .si(net14632) );
  dffe_SIZE1 i_mul_frac_in2_54 ( .din(inq_in2_54), .en(m6stg_step), .clk(rclk), 
        .q(mul_frac_in2_54), .se(se), .si(net14631) );
  dffe_SIZE1 i_mul_frac_in2_53_0_neq_0 ( .din(inq_in2_53_0_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in2_53_0_neq_0), .se(se), .si(
        net14630) );
  dffe_SIZE1 i_mul_frac_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in2_50_0_neq_0), .se(se), .si(
        net14629) );
  dffe_SIZE1 i_mul_frac_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        m6stg_step), .clk(rclk), .q(mul_frac_in2_53_32_neq_0), .se(se), .si(
        net14628) );
  dffe_SIZE1 i_mul_exp_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(m6stg_step), 
        .clk(rclk), .q(mul_exp_in2_exp_eq_0), .se(se), .si(net14627) );
  dffe_SIZE1 i_mul_exp_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        m6stg_step), .clk(rclk), .q(mul_exp_in2_exp_neq_ffs), .se(se), .si(
        net14626) );
  dffe_SIZE1 i_m2stg_snan_in1 ( .din(m1stg_snan_in1), .en(m6stg_step), .clk(
        rclk), .q(m2stg_snan_in1), .se(se), .si(net14625) );
  dffe_SIZE1 i_m2stg_snan_in2 ( .din(m1stg_snan_in2), .en(m6stg_step), .clk(
        rclk), .q(m2stg_snan_in2), .se(se), .si(net14624) );
  dffe_SIZE1 i_m2stg_qnan_in1 ( .din(m1stg_qnan_in1), .en(m6stg_step), .clk(
        rclk), .q(m2stg_qnan_in1), .se(se), .si(net14623) );
  dffe_SIZE1 i_m2stg_qnan_in2 ( .din(m1stg_qnan_in2), .en(m6stg_step), .clk(
        rclk), .q(m2stg_qnan_in2), .se(se), .si(net14622) );
  dffe_SIZE1 i_m2stg_nan_in2 ( .din(m1stg_nan_in2), .en(m6stg_step), .clk(rclk), .q(m2stg_nan_in2), .se(se), .si(net14621) );
  dffe_SIZE1 i_m2stg_inf_in1 ( .din(m1stg_inf_in1), .en(m6stg_step), .clk(rclk), .q(m2stg_inf_in1), .se(se), .si(net14620) );
  dffe_SIZE1 i_m2stg_inf_in2 ( .din(m1stg_inf_in2), .en(m6stg_step), .clk(rclk), .q(m2stg_inf_in2), .se(se), .si(net14619) );
  dffe_SIZE1 i_m2stg_inf_in ( .din(m1stg_inf_in), .en(m6stg_step), .clk(rclk), 
        .q(m2stg_inf_in), .se(se), .si(net14618) );
  dffe_SIZE1 i_m2stg_zero_in1 ( .din(m1stg_zero_in1), .en(m6stg_step), .clk(
        rclk), .q(m2stg_zero_in1), .se(se), .si(net14617) );
  dffe_SIZE1 i_m2stg_zero_in2 ( .din(m1stg_zero_in2), .en(m6stg_step), .clk(
        rclk), .q(m2stg_zero_in2), .se(se), .si(net14616) );
  dffe_SIZE1 i_m2stg_zero_in ( .din(m1stg_zero_in), .en(m6stg_step), .clk(rclk), .q(m2stg_zero_in), .se(se), .si(net14615) );
  dff_SIZE8 i_m1stg_op ( .din(m1stg_op_in), .clk(rclk), .q(m1stg_op), .se(se), 
        .si({net14607, net14608, net14609, net14610, net14611, net14612, 
        net14613, net14614}) );
  dff_SIZE1 i_m1stg_mul ( .din(m1stg_mul_in), .clk(rclk), .q(m1stg_mul), .se(
        se), .si(net14606) );
  dffe_SIZE1 i_m1stg_sngop ( .din(inq_op[0]), .en(m6stg_step), .clk(rclk), .q(
        m1stg_sngop), .se(se), .si(net14605) );
  dffe_SIZE4 i_m1stg_sngopa ( .din({inq_op[0], inq_op[0], inq_op[0], inq_op[0]}), .en(m6stg_step), .clk(rclk), .q(m1stg_sngopa), .se(se), .si({net14601, 
        net14602, net14603, net14604}) );
  dffe_SIZE1 i_m1stg_dblop ( .din(inq_op[1]), .en(m6stg_step), .clk(rclk), .q(
        m1stg_dblop), .se(se), .si(net14600) );
  dffe_SIZE4 i_m1stg_dblopa ( .din({inq_op[1], inq_op[1], inq_op[1], inq_op[1]}), .en(m6stg_step), .clk(rclk), .q(m1stg_dblopa), .se(se), .si({net14596, 
        net14597, net14598, net14599}) );
  dffe_SIZE1 i_m1stg_dblop_inv ( .din(m1stg_dblop_inv_in), .en(m6stg_step), 
        .clk(rclk), .q(m1stg_dblop_inv), .se(se), .si(net14595) );
  dffe_SIZE2 i_m1stg_rnd_mode ( .din(inq_rnd_mode), .en(m6stg_step), .clk(rclk), .q(m1stg_rnd_mode), .se(se), .si({net14593, net14594}) );
  dffe_SIZE5 i_m1stg_id ( .din(inq_id), .en(m6stg_step), .clk(rclk), .q(
        m1stg_id), .se(se), .si({net14588, net14589, net14590, net14591, 
        net14592}) );
  dffre_SIZE5 i_m2stg_opdec ( .din({m1stg_fmul, m1stg_opdec[3], N53, N44, N62}), .rst(reset), .en(m6stg_step), .clk(rclk), .q({m2stg_opdec, m2stg_fmuls, 
        m2stg_fmuld, m2stg_fsmuld}), .se(se), .si({net14583, net14584, 
        net14585, net14586, net14587}) );
  dffe_SIZE2 i_m2stg_rnd_mode ( .din(m1stg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m2stg_rnd_mode), .se(se), .si({net14581, net14582}) );
  dffe_SIZE5 i_m2stg_id ( .din(m1stg_id), .en(m6stg_step), .clk(rclk), .q(
        m2stg_id), .se(se), .si({net14576, net14577, net14578, net14579, 
        net14580}) );
  dffre_SIZE4 i_m3astg_opdec ( .din({m2stg_opdec, m2stg_fmuls, m2stg_fmuld}), 
        .rst(reset), .en(m6stg_step), .clk(rclk), .q(m3astg_opdec), .se(se), 
        .si({net14572, net14573, net14574, net14575}) );
  dffe_SIZE2 i_m3astg_rnd_mode ( .din(m2stg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m3astg_rnd_mode), .se(se), .si({net14570, net14571}) );
  dffe_SIZE5 i_m3astg_id ( .din(m2stg_id), .en(m6stg_step), .clk(rclk), .q(
        m3astg_id), .se(se), .si({net14565, net14566, net14567, net14568, 
        net14569}) );
  dffre_SIZE4 i_m3bstg_opdec ( .din(m3astg_opdec), .rst(reset), .en(m6stg_step), .clk(rclk), .q(m3bstg_opdec), .se(se), .si({net14561, net14562, net14563, 
        net14564}) );
  dffe_SIZE2 i_m3bstg_rnd_mode ( .din(m3astg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m3bstg_rnd_mode), .se(se), .si({net14559, net14560}) );
  dffe_SIZE5 i_m3bstg_id ( .din(m3astg_id), .en(m6stg_step), .clk(rclk), .q(
        m3bstg_id), .se(se), .si({net14554, net14555, net14556, net14557, 
        net14558}) );
  dffre_SIZE4 i_m3stg_opdec ( .din(m3bstg_opdec), .rst(reset), .en(m6stg_step), 
        .clk(rclk), .q(m3stg_opdec), .se(se), .si({net14550, net14551, 
        net14552, net14553}) );
  dffe_SIZE2 i_m3stg_rnd_mode ( .din(m3bstg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m3stg_rnd_mode), .se(se), .si({net14548, net14549}) );
  dffe_SIZE5 i_m3stg_id ( .din(m3bstg_id), .en(m6stg_step), .clk(rclk), .q(
        m3stg_id), .se(se), .si({net14543, net14544, net14545, net14546, 
        net14547}) );
  dffre_SIZE4 i_m4stg_opdec ( .din(m3stg_opdec), .rst(reset), .en(m6stg_step), 
        .clk(rclk), .q(m4stg_opdec), .se(se), .si({net14539, net14540, 
        net14541, net14542}) );
  dffe_SIZE2 i_m4stg_rnd_mode ( .din(m3stg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m4stg_rnd_mode), .se(se), .si({net14537, net14538}) );
  dffe_SIZE5 i_m4stg_id ( .din(m3stg_id), .en(m6stg_step), .clk(rclk), .q(
        m4stg_id), .se(se), .si({net14532, net14533, net14534, net14535, 
        net14536}) );
  dffre_SIZE4 i_m5stg_opdec ( .din(m4stg_opdec), .rst(reset), .en(m6stg_step), 
        .clk(rclk), .q({m5stg_opdec, m5stg_fmuls, m5stg_fmuld}), .se(se), .si(
        {net14528, net14529, net14530, net14531}) );
  dffe_SIZE2 i_m5stg_rnd_mode ( .din(m4stg_rnd_mode), .en(m6stg_step), .clk(
        rclk), .q(m5stg_rnd_mode), .se(se), .si({net14526, net14527}) );
  dffe_SIZE5 i_m5stg_id ( .din(m4stg_id), .en(m6stg_step), .clk(rclk), .q(
        m5stg_id), .se(se), .si({net14521, net14522, net14523, net14524, 
        net14525}) );
  dffre_SIZE1 i_m5stg_fmulda ( .din(m4stg_opdec[1]), .rst(reset), .en(
        m6stg_step), .clk(rclk), .q(m5stg_fmulda), .se(se), .si(net14520) );
  dffre_SIZE3 i_m6stg_opdec ( .din({m5stg_opdec, m5stg_fmuls}), .rst(reset), 
        .en(m6stg_step), .clk(rclk), .q({m6stg_opdec[4], m6stg_fmul_dbl_dst, 
        m6stg_fmuls}), .se(se), .si({net14517, net14518, net14519}) );
  dffe_SIZE10 i_m6stg_id ( .din(m6stg_id_in), .en(m6stg_step), .clk(rclk), .q(
        m6stg_id), .se(se), .si({net14507, net14508, net14509, net14510, 
        net14511, net14512, net14513, net14514, net14515, net14516}) );
  dffre_SIZE1 i_mul_pipe_active ( .din(mul_pipe_active_in), .rst(reset), .en(
        1'b1), .clk(rclk), .q(mul_pipe_active), .se(se), .si(net14506) );
  dffe_SIZE1 i_m1stg_sign1 ( .din(inq_in1_63), .en(m6stg_step), .clk(rclk), 
        .q(m1stg_sign1), .se(se), .si(net14505) );
  dffe_SIZE1 i_m1stg_sign2 ( .din(inq_in2_63), .en(m6stg_step), .clk(rclk), 
        .q(m1stg_sign2), .se(se), .si(net14504) );
  dffe_SIZE1 i_m2stg_sign1 ( .din(m1stg_sign1), .en(m6stg_step), .clk(rclk), 
        .q(m2stg_sign1), .se(se), .si(net14503) );
  dffe_SIZE1 i_m2stg_sign2 ( .din(m1stg_sign2), .en(m6stg_step), .clk(rclk), 
        .q(m2stg_sign2), .se(se), .si(net14502) );
  dffe_SIZE1 i_m2stg_of_mask ( .din(m1stg_of_mask), .en(m6stg_step), .clk(rclk), .q(m2stg_of_mask), .se(se), .si(net14501) );
  dffe_SIZE1 i_m3astg_sign ( .din(m2stg_sign), .en(m6stg_step), .clk(rclk), 
        .q(m3astg_sign), .se(se), .si(net14500) );
  dffe_SIZE1 i_m3astg_nv ( .din(m2stg_nv), .en(m6stg_step), .clk(rclk), .q(
        m3astg_nv), .se(se), .si(net14499) );
  dffe_SIZE1 i_m3astg_of_mask ( .din(m2stg_of_mask), .en(m6stg_step), .clk(
        rclk), .q(m3astg_of_mask), .se(se), .si(net14498) );
  dffe_SIZE1 i_m3bstg_sign ( .din(m3astg_sign), .en(m6stg_step), .clk(rclk), 
        .q(m3bstg_sign), .se(se), .si(net14497) );
  dffe_SIZE1 i_m3bstg_nv ( .din(m3astg_nv), .en(m6stg_step), .clk(rclk), .q(
        m3bstg_nv), .se(se), .si(net14496) );
  dffe_SIZE1 i_m3bstg_of_mask ( .din(m3astg_of_mask), .en(m6stg_step), .clk(
        rclk), .q(m3bstg_of_mask), .se(se), .si(net14495) );
  dffe_SIZE1 i_m3stg_sign ( .din(m3bstg_sign), .en(m6stg_step), .clk(rclk), 
        .q(m3stg_sign), .se(se), .si(net14494) );
  dffe_SIZE1 i_m3stg_nv ( .din(m3bstg_nv), .en(m6stg_step), .clk(rclk), .q(
        m3stg_nv), .se(se), .si(net14493) );
  dffe_SIZE1 i_m3stg_of_mask ( .din(m3bstg_of_mask), .en(m6stg_step), .clk(
        rclk), .q(m3stg_of_mask), .se(se), .si(net14492) );
  dffe_SIZE1 i_m4stg_sign ( .din(m3stg_sign), .en(m6stg_step), .clk(rclk), .q(
        m4stg_sign), .se(se), .si(net14491) );
  dffe_SIZE1 i_m4stg_nv ( .din(m3stg_nv), .en(m6stg_step), .clk(rclk), .q(
        m4stg_nv), .se(se), .si(net14490) );
  dffe_SIZE1 i_m4stg_of_mask ( .din(m3stg_of_mask), .en(m6stg_step), .clk(rclk), .q(m4stg_of_mask), .se(se), .si(net14489) );
  dffe_SIZE1 i_m5stg_sign ( .din(m4stg_sign), .en(m6stg_step), .clk(rclk), .q(
        m5stg_sign), .se(se), .si(net14488) );
  dffe_SIZE1 i_m5stg_nv ( .din(m4stg_nv), .en(m6stg_step), .clk(rclk), .q(
        m5stg_nv), .se(se), .si(net14487) );
  dffe_SIZE1 i_m5stg_of_mask ( .din(m4stg_of_mask), .en(m6stg_step), .clk(rclk), .q(m5stg_of_mask), .se(se), .si(net14486) );
  dffe_SIZE1 i_mul_sign_out ( .din(m5stg_sign), .en(m6stg_step), .clk(rclk), 
        .q(mul_sign_out), .se(se), .si(net14485) );
  dffe_SIZE1 i_mul_nv_out ( .din(m5stg_nv), .en(m6stg_step), .clk(rclk), .q(
        mul_exc_out[4]), .se(se), .si(net14484) );
  dffe_SIZE1 i_mul_of_out_tmp1 ( .din(mul_of_out_tmp1_in), .en(m6stg_step), 
        .clk(rclk), .q(mul_of_out_tmp1), .se(se), .si(net14483) );
  dffe_SIZE1 i_mul_of_out_tmp2 ( .din(m5stg_in_of), .en(m6stg_step), .clk(rclk), .q(mul_of_out_tmp2), .se(se), .si(net14482) );
  dffe_SIZE1 i_mul_of_out_cout ( .din(m5stg_fracadd_cout), .en(m6stg_step), 
        .clk(rclk), .q(mul_of_out_cout), .se(se), .si(net14481) );
  dffe_SIZE1 i_mul_uf_out ( .din(mul_uf_out_in), .en(m6stg_step), .clk(rclk), 
        .q(mul_exc_out[2]), .se(se), .si(net14480) );
  dffe_SIZE1 i_mul_nx_out ( .din(mul_nx_out_in), .en(m6stg_step), .clk(rclk), 
        .q(mul_nx_out), .se(se), .si(net14479) );
  dffe_SIZE6 i_m2stg_ld0_1 ( .din(m2stg_ld0_1_in), .en(m6stg_step), .clk(rclk), 
        .q(m2stg_ld0_1), .se(se), .si({net14473, net14474, net14475, net14476, 
        net14477, net14478}) );
  dffe_SIZE6 i_m2stg_ld0_2 ( .din(m2stg_ld0_2_in), .en(m6stg_step), .clk(rclk), 
        .q(m2stg_ld0_2), .se(se), .si({net14467, net14468, net14469, net14470, 
        net14471, net14472}) );
  dffe_SIZE7 i_m3astg_ld0_inv ( .din(m2stg_ld0_inv), .en(m6stg_step), .clk(
        rclk), .q(m3astg_ld0_inv), .se(se), .si({net14460, net14461, net14462, 
        net14463, net14464, net14465, net14466}) );
  dffe_SIZE7 i_m3bstg_ld0_inv ( .din(m3astg_ld0_inv), .en(m6stg_step), .clk(
        rclk), .q(m3bstg_ld0_inv), .se(se), .si({net14453, net14454, net14455, 
        net14456, net14457, net14458, net14459}) );
  dffe_SIZE1 i_m4stg_expadd_eq_0 ( .din(m3stg_expadd_eq_0), .en(m6stg_step), 
        .clk(rclk), .q(m4stg_expadd_eq_0), .se(se), .si(net14452) );
  dffe_SIZE1 i_m4stg_right_shift ( .din(m4stg_right_shift_in), .en(m6stg_step), 
        .clk(rclk), .q(m4stg_right_shift), .se(se), .si(net14451) );
  GTECH_AND2 C162 ( .A(m5stg_id[3]), .B(m5stg_id[4]), .Z(N8) );
  GTECH_AND2 C163 ( .A(m5stg_id[2]), .B(N8), .Z(N9) );
  GTECH_NOT I_0 ( .A(m5stg_id[4]), .Z(N10) );
  GTECH_NOT I_1 ( .A(m5stg_id[3]), .Z(N11) );
  GTECH_OR2 C166 ( .A(N11), .B(N10), .Z(N12) );
  GTECH_OR2 C167 ( .A(m5stg_id[2]), .B(N12), .Z(N13) );
  GTECH_NOT I_2 ( .A(N13), .Z(N14) );
  GTECH_NOT I_3 ( .A(m5stg_id[2]), .Z(N15) );
  GTECH_OR2 C171 ( .A(m5stg_id[3]), .B(N10), .Z(N16) );
  GTECH_OR2 C172 ( .A(N15), .B(N16), .Z(N17) );
  GTECH_NOT I_4 ( .A(N17), .Z(N18) );
  GTECH_OR2 C175 ( .A(m5stg_id[3]), .B(N10), .Z(N19) );
  GTECH_OR2 C176 ( .A(m5stg_id[2]), .B(N19), .Z(N20) );
  GTECH_NOT I_5 ( .A(N20), .Z(N21) );
  GTECH_OR2 C180 ( .A(N11), .B(m5stg_id[4]), .Z(N22) );
  GTECH_OR2 C181 ( .A(N15), .B(N22), .Z(N23) );
  GTECH_NOT I_6 ( .A(N23), .Z(N24) );
  GTECH_OR2 C184 ( .A(N11), .B(m5stg_id[4]), .Z(N25) );
  GTECH_OR2 C185 ( .A(m5stg_id[2]), .B(N25), .Z(N26) );
  GTECH_NOT I_7 ( .A(N26), .Z(N27) );
  GTECH_OR2 C188 ( .A(m5stg_id[3]), .B(m5stg_id[4]), .Z(N28) );
  GTECH_OR2 C189 ( .A(N15), .B(N28), .Z(N29) );
  GTECH_NOT I_8 ( .A(N29), .Z(N30) );
  GTECH_OR2 C191 ( .A(m5stg_id[3]), .B(m5stg_id[4]), .Z(N31) );
  GTECH_OR2 C192 ( .A(m5stg_id[2]), .B(N31), .Z(N32) );
  GTECH_NOT I_9 ( .A(N32), .Z(N33) );
  GTECH_NOT I_10 ( .A(m1stg_op[6]), .Z(N34) );
  GTECH_NOT I_11 ( .A(m1stg_op[3]), .Z(N35) );
  GTECH_NOT I_12 ( .A(m1stg_op[1]), .Z(N36) );
  GTECH_OR2 C197 ( .A(N34), .B(m1stg_op[7]), .Z(N37) );
  GTECH_OR2 C198 ( .A(m1stg_op[5]), .B(N37), .Z(N38) );
  GTECH_OR2 C199 ( .A(m1stg_op[4]), .B(N38), .Z(N39) );
  GTECH_OR2 C200 ( .A(N35), .B(N39), .Z(N40) );
  GTECH_OR2 C201 ( .A(m1stg_op[2]), .B(N40), .Z(N41) );
  GTECH_OR2 C202 ( .A(N36), .B(N41), .Z(N42) );
  GTECH_OR2 C203 ( .A(m1stg_op[0]), .B(N42), .Z(N43) );
  GTECH_NOT I_13 ( .A(N43), .Z(N44) );
  GTECH_NOT I_14 ( .A(m1stg_op[0]), .Z(N45) );
  GTECH_OR2 C208 ( .A(N34), .B(m1stg_op[7]), .Z(N46) );
  GTECH_OR2 C209 ( .A(m1stg_op[5]), .B(N46), .Z(N47) );
  GTECH_OR2 C210 ( .A(m1stg_op[4]), .B(N47), .Z(N48) );
  GTECH_OR2 C211 ( .A(N35), .B(N48), .Z(N49) );
  GTECH_OR2 C212 ( .A(m1stg_op[2]), .B(N49), .Z(N50) );
  GTECH_OR2 C213 ( .A(m1stg_op[1]), .B(N50), .Z(N51) );
  GTECH_OR2 C214 ( .A(N45), .B(N51), .Z(N52) );
  GTECH_NOT I_15 ( .A(N52), .Z(N53) );
  GTECH_NOT I_16 ( .A(m1stg_op[5]), .Z(N54) );
  GTECH_OR2 C220 ( .A(N34), .B(m1stg_op[7]), .Z(N55) );
  GTECH_OR2 C221 ( .A(N54), .B(N55), .Z(N56) );
  GTECH_OR2 C222 ( .A(m1stg_op[4]), .B(N56), .Z(N57) );
  GTECH_OR2 C223 ( .A(N35), .B(N57), .Z(N58) );
  GTECH_OR2 C224 ( .A(m1stg_op[2]), .B(N58), .Z(N59) );
  GTECH_OR2 C225 ( .A(m1stg_op[1]), .B(N59), .Z(N60) );
  GTECH_OR2 C226 ( .A(N45), .B(N60), .Z(N61) );
  GTECH_NOT I_17 ( .A(N61), .Z(N62) );
  GTECH_OR2 C231 ( .A(N34), .B(m1stg_op[7]), .Z(N63) );
  GTECH_OR2 C232 ( .A(m1stg_op[5]), .B(N63), .Z(N64) );
  GTECH_OR2 C233 ( .A(m1stg_op[4]), .B(N64), .Z(N65) );
  GTECH_OR2 C234 ( .A(N35), .B(N65), .Z(N66) );
  GTECH_OR2 C235 ( .A(m1stg_op[2]), .B(N66), .Z(N67) );
  GTECH_OR2 C236 ( .A(N36), .B(N67), .Z(N68) );
  GTECH_OR2 C237 ( .A(m1stg_op[0]), .B(N68), .Z(N69) );
  GTECH_NOT I_18 ( .A(N69), .Z(N70) );
  GTECH_OR2 C243 ( .A(N34), .B(m1stg_op[7]), .Z(N71) );
  GTECH_OR2 C244 ( .A(N54), .B(N71), .Z(N72) );
  GTECH_OR2 C245 ( .A(m1stg_op[4]), .B(N72), .Z(N73) );
  GTECH_OR2 C246 ( .A(N35), .B(N73), .Z(N74) );
  GTECH_OR2 C247 ( .A(m1stg_op[2]), .B(N74), .Z(N75) );
  GTECH_OR2 C248 ( .A(m1stg_op[1]), .B(N75), .Z(N76) );
  GTECH_OR2 C249 ( .A(N45), .B(N76), .Z(N77) );
  GTECH_NOT I_19 ( .A(N77), .Z(N78) );
  GTECH_NOT I_20 ( .A(m5stg_rnd_mode[0]), .Z(N79) );
  GTECH_OR2 C252 ( .A(N79), .B(m5stg_rnd_mode[1]), .Z(N80) );
  GTECH_NOT I_21 ( .A(N80), .Z(N81) );
  GTECH_NOT I_22 ( .A(m5stg_rnd_mode[1]), .Z(N82) );
  GTECH_OR2 C255 ( .A(m5stg_rnd_mode[0]), .B(N82), .Z(N83) );
  GTECH_NOT I_23 ( .A(N83), .Z(N84) );
  GTECH_AND2 C257 ( .A(m5stg_rnd_mode[0]), .B(m5stg_rnd_mode[1]), .Z(N85) );
  GTECH_OR2 C261 ( .A(N34), .B(m1stg_op[7]), .Z(N86) );
  GTECH_OR2 C262 ( .A(m1stg_op[5]), .B(N86), .Z(N87) );
  GTECH_OR2 C263 ( .A(m1stg_op[4]), .B(N87), .Z(N88) );
  GTECH_OR2 C264 ( .A(N35), .B(N88), .Z(N89) );
  GTECH_OR2 C265 ( .A(m1stg_op[2]), .B(N89), .Z(N90) );
  GTECH_OR2 C266 ( .A(m1stg_op[1]), .B(N90), .Z(N91) );
  GTECH_OR2 C267 ( .A(N45), .B(N91), .Z(N92) );
  GTECH_NOT I_24 ( .A(N92), .Z(N93) );
  GTECH_OR2 C272 ( .A(N34), .B(m1stg_op[7]), .Z(N94) );
  GTECH_OR2 C273 ( .A(m1stg_op[5]), .B(N94), .Z(N95) );
  GTECH_OR2 C274 ( .A(m1stg_op[4]), .B(N95), .Z(N96) );
  GTECH_OR2 C275 ( .A(N35), .B(N96), .Z(N97) );
  GTECH_OR2 C276 ( .A(m1stg_op[2]), .B(N97), .Z(N98) );
  GTECH_OR2 C277 ( .A(N36), .B(N98), .Z(N99) );
  GTECH_OR2 C278 ( .A(m1stg_op[0]), .B(N99), .Z(N100) );
  GTECH_NOT I_25 ( .A(N100), .Z(N101) );
  GTECH_OR2 C284 ( .A(N34), .B(m1stg_op[7]), .Z(N102) );
  GTECH_OR2 C285 ( .A(N54), .B(N102), .Z(N103) );
  GTECH_OR2 C286 ( .A(m1stg_op[4]), .B(N103), .Z(N104) );
  GTECH_OR2 C287 ( .A(N35), .B(N104), .Z(N105) );
  GTECH_OR2 C288 ( .A(m1stg_op[2]), .B(N105), .Z(N106) );
  GTECH_OR2 C289 ( .A(m1stg_op[1]), .B(N106), .Z(N107) );
  GTECH_OR2 C290 ( .A(N45), .B(N107), .Z(N108) );
  GTECH_NOT I_26 ( .A(N108), .Z(N109) );
  GTECH_OR2 C293 ( .A(m5stg_rnd_mode[0]), .B(N82), .Z(N110) );
  GTECH_NOT I_27 ( .A(N110), .Z(N111) );
  GTECH_OR2 C295 ( .A(m5stg_frac[1]), .B(m5stg_frac[2]), .Z(N112) );
  GTECH_OR2 C296 ( .A(m5stg_frac[0]), .B(N112), .Z(N113) );
  GTECH_AND2 C299 ( .A(m5stg_rnd_mode[0]), .B(m5stg_rnd_mode[1]), .Z(N114) );
  GTECH_OR2 C304 ( .A(m5stg_rnd_mode[0]), .B(m5stg_rnd_mode[1]), .Z(N115) );
  GTECH_NOT I_28 ( .A(N115), .Z(N116) );
  GTECH_OR2 C306 ( .A(m5stg_frac[0]), .B(m5stg_frac[1]), .Z(N117) );
  GTECH_OR2 C310 ( .A(m5stg_rnd_mode[0]), .B(N82), .Z(N118) );
  GTECH_NOT I_29 ( .A(N118), .Z(N119) );
  GTECH_OR2 C312 ( .A(m5stg_frac[30]), .B(m5stg_frac[31]), .Z(N120) );
  GTECH_OR2 C313 ( .A(m5stg_frac[29]), .B(N120), .Z(N121) );
  GTECH_OR2 C314 ( .A(m5stg_frac[28]), .B(N121), .Z(N122) );
  GTECH_OR2 C315 ( .A(m5stg_frac[27]), .B(N122), .Z(N123) );
  GTECH_OR2 C316 ( .A(m5stg_frac[26]), .B(N123), .Z(N124) );
  GTECH_OR2 C317 ( .A(m5stg_frac[25]), .B(N124), .Z(N125) );
  GTECH_OR2 C318 ( .A(m5stg_frac[24]), .B(N125), .Z(N126) );
  GTECH_OR2 C319 ( .A(m5stg_frac[23]), .B(N126), .Z(N127) );
  GTECH_OR2 C320 ( .A(m5stg_frac[22]), .B(N127), .Z(N128) );
  GTECH_OR2 C321 ( .A(m5stg_frac[21]), .B(N128), .Z(N129) );
  GTECH_OR2 C322 ( .A(m5stg_frac[20]), .B(N129), .Z(N130) );
  GTECH_OR2 C323 ( .A(m5stg_frac[19]), .B(N130), .Z(N131) );
  GTECH_OR2 C324 ( .A(m5stg_frac[18]), .B(N131), .Z(N132) );
  GTECH_OR2 C325 ( .A(m5stg_frac[17]), .B(N132), .Z(N133) );
  GTECH_OR2 C326 ( .A(m5stg_frac[16]), .B(N133), .Z(N134) );
  GTECH_OR2 C327 ( .A(m5stg_frac[15]), .B(N134), .Z(N135) );
  GTECH_OR2 C328 ( .A(m5stg_frac[14]), .B(N135), .Z(N136) );
  GTECH_OR2 C329 ( .A(m5stg_frac[13]), .B(N136), .Z(N137) );
  GTECH_OR2 C330 ( .A(m5stg_frac[12]), .B(N137), .Z(N138) );
  GTECH_OR2 C331 ( .A(m5stg_frac[11]), .B(N138), .Z(N139) );
  GTECH_OR2 C332 ( .A(m5stg_frac[10]), .B(N139), .Z(N140) );
  GTECH_OR2 C333 ( .A(m5stg_frac[9]), .B(N140), .Z(N141) );
  GTECH_OR2 C334 ( .A(m5stg_frac[8]), .B(N141), .Z(N142) );
  GTECH_OR2 C335 ( .A(m5stg_frac[7]), .B(N142), .Z(N143) );
  GTECH_OR2 C336 ( .A(m5stg_frac[6]), .B(N143), .Z(N144) );
  GTECH_OR2 C337 ( .A(m5stg_frac[5]), .B(N144), .Z(N145) );
  GTECH_OR2 C338 ( .A(m5stg_frac[4]), .B(N145), .Z(N146) );
  GTECH_OR2 C339 ( .A(m5stg_frac[3]), .B(N146), .Z(N147) );
  GTECH_OR2 C340 ( .A(m5stg_frac[2]), .B(N147), .Z(N148) );
  GTECH_OR2 C341 ( .A(m5stg_frac[1]), .B(N148), .Z(N149) );
  GTECH_OR2 C342 ( .A(m5stg_frac[0]), .B(N149), .Z(N150) );
  GTECH_AND2 C345 ( .A(m5stg_rnd_mode[0]), .B(m5stg_rnd_mode[1]), .Z(N151) );
  GTECH_OR2 C379 ( .A(m5stg_rnd_mode[0]), .B(m5stg_rnd_mode[1]), .Z(N152) );
  GTECH_NOT I_30 ( .A(N152), .Z(N153) );
  GTECH_OR2 C381 ( .A(m5stg_frac[29]), .B(m5stg_frac[30]), .Z(N154) );
  GTECH_OR2 C382 ( .A(m5stg_frac[28]), .B(N154), .Z(N155) );
  GTECH_OR2 C383 ( .A(m5stg_frac[27]), .B(N155), .Z(N156) );
  GTECH_OR2 C384 ( .A(m5stg_frac[26]), .B(N156), .Z(N157) );
  GTECH_OR2 C385 ( .A(m5stg_frac[25]), .B(N157), .Z(N158) );
  GTECH_OR2 C386 ( .A(m5stg_frac[24]), .B(N158), .Z(N159) );
  GTECH_OR2 C387 ( .A(m5stg_frac[23]), .B(N159), .Z(N160) );
  GTECH_OR2 C388 ( .A(m5stg_frac[22]), .B(N160), .Z(N161) );
  GTECH_OR2 C389 ( .A(m5stg_frac[21]), .B(N161), .Z(N162) );
  GTECH_OR2 C390 ( .A(m5stg_frac[20]), .B(N162), .Z(N163) );
  GTECH_OR2 C391 ( .A(m5stg_frac[19]), .B(N163), .Z(N164) );
  GTECH_OR2 C392 ( .A(m5stg_frac[18]), .B(N164), .Z(N165) );
  GTECH_OR2 C393 ( .A(m5stg_frac[17]), .B(N165), .Z(N166) );
  GTECH_OR2 C394 ( .A(m5stg_frac[16]), .B(N166), .Z(N167) );
  GTECH_OR2 C395 ( .A(m5stg_frac[15]), .B(N167), .Z(N168) );
  GTECH_OR2 C396 ( .A(m5stg_frac[14]), .B(N168), .Z(N169) );
  GTECH_OR2 C397 ( .A(m5stg_frac[13]), .B(N169), .Z(N170) );
  GTECH_OR2 C398 ( .A(m5stg_frac[12]), .B(N170), .Z(N171) );
  GTECH_OR2 C399 ( .A(m5stg_frac[11]), .B(N171), .Z(N172) );
  GTECH_OR2 C400 ( .A(m5stg_frac[10]), .B(N172), .Z(N173) );
  GTECH_OR2 C401 ( .A(m5stg_frac[9]), .B(N173), .Z(N174) );
  GTECH_OR2 C402 ( .A(m5stg_frac[8]), .B(N174), .Z(N175) );
  GTECH_OR2 C403 ( .A(m5stg_frac[7]), .B(N175), .Z(N176) );
  GTECH_OR2 C404 ( .A(m5stg_frac[6]), .B(N176), .Z(N177) );
  GTECH_OR2 C405 ( .A(m5stg_frac[5]), .B(N177), .Z(N178) );
  GTECH_OR2 C406 ( .A(m5stg_frac[4]), .B(N178), .Z(N179) );
  GTECH_OR2 C407 ( .A(m5stg_frac[3]), .B(N179), .Z(N180) );
  GTECH_OR2 C408 ( .A(m5stg_frac[2]), .B(N180), .Z(N181) );
  GTECH_OR2 C409 ( .A(m5stg_frac[1]), .B(N181), .Z(N182) );
  GTECH_OR2 C410 ( .A(m5stg_frac[0]), .B(N182), .Z(N183) );
  ADD_UNS_OP add_2061 ( .A(m2stg_ld0_1), .B(m2stg_ld0_2), .Z(m2stg_ld0) );
  ADD_UNS_OP add_2136 ( .A(m3stg_exp[5:0]), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1}), .Z(m3stg_exp_minus1) );
  ADD_UNS_OP add_2139_ni_cf ( .A(1'b1), .B({N184, N185, N186, N187, N188, N189}), .Z(m3stg_exp_inv_plus2) );
  SUB_UNS_OP sub_add_2139_b0 ( .A(1'b0), .B(m3stg_exp[5:0]), .Z({N184, N185, 
        N186, N187, N188, N189}) );
  GTECH_NOT I_31 ( .A(mula_rst_l), .Z(reset) );
  GTECH_AND2 C416 ( .A(mul_exp_in1_exp_eq_0), .B(m1stg_sngopa[0]), .Z(
        m1stg_denorm_sng_in1) );
  GTECH_AND2 C417 ( .A(mul_exp_in1_exp_eq_0), .B(m1stg_dblopa[0]), .Z(
        m1stg_denorm_dbl_in1) );
  GTECH_AND2 C418 ( .A(mul_exp_in2_exp_eq_0), .B(m1stg_sngopa[0]), .Z(
        m1stg_denorm_sng_in2) );
  GTECH_AND2 C419 ( .A(mul_exp_in2_exp_eq_0), .B(m1stg_dblopa[0]), .Z(
        m1stg_denorm_dbl_in2) );
  GTECH_OR2 C420 ( .A(m1stg_denorm_sng_in1), .B(m1stg_denorm_dbl_in1), .Z(
        m1stg_denorm_in1) );
  GTECH_OR2 C421 ( .A(m1stg_denorm_sng_in2), .B(m1stg_denorm_dbl_in2), .Z(
        m1stg_denorm_in2) );
  GTECH_AND2 C422 ( .A(N190), .B(m1stg_sngopa[0]), .Z(m1stg_norm_sng_in1) );
  GTECH_NOT I_32 ( .A(mul_exp_in1_exp_eq_0), .Z(N190) );
  GTECH_AND2 C424 ( .A(N190), .B(m1stg_dblopa[0]), .Z(m1stg_norm_dbl_in1) );
  GTECH_AND2 C426 ( .A(N191), .B(m1stg_sngopa[0]), .Z(m1stg_norm_sng_in2) );
  GTECH_NOT I_33 ( .A(mul_exp_in2_exp_eq_0), .Z(N191) );
  GTECH_AND2 C428 ( .A(N191), .B(m1stg_dblopa[0]), .Z(m1stg_norm_dbl_in2) );
  GTECH_AND2 C430 ( .A(N195), .B(m1stg_sngopa[1]), .Z(m1stg_snan_sng_in1) );
  GTECH_AND2 C431 ( .A(N194), .B(mul_frac_in1_53_32_neq_0), .Z(N195) );
  GTECH_AND2 C432 ( .A(N192), .B(N193), .Z(N194) );
  GTECH_NOT I_34 ( .A(mul_exp_in1_exp_neq_ffs), .Z(N192) );
  GTECH_NOT I_35 ( .A(mul_frac_in1_54), .Z(N193) );
  GTECH_AND2 C435 ( .A(N198), .B(m1stg_dblopa[1]), .Z(m1stg_snan_dbl_in1) );
  GTECH_AND2 C436 ( .A(N197), .B(mul_frac_in1_50_0_neq_0), .Z(N198) );
  GTECH_AND2 C437 ( .A(N192), .B(N196), .Z(N197) );
  GTECH_NOT I_36 ( .A(mul_frac_in1_51), .Z(N196) );
  GTECH_AND2 C440 ( .A(N202), .B(m1stg_sngopa[1]), .Z(m1stg_snan_sng_in2) );
  GTECH_AND2 C441 ( .A(N201), .B(mul_frac_in2_53_32_neq_0), .Z(N202) );
  GTECH_AND2 C442 ( .A(N199), .B(N200), .Z(N201) );
  GTECH_NOT I_37 ( .A(mul_exp_in2_exp_neq_ffs), .Z(N199) );
  GTECH_NOT I_38 ( .A(mul_frac_in2_54), .Z(N200) );
  GTECH_AND2 C445 ( .A(N205), .B(m1stg_dblopa[1]), .Z(m1stg_snan_dbl_in2) );
  GTECH_AND2 C446 ( .A(N204), .B(mul_frac_in2_50_0_neq_0), .Z(N205) );
  GTECH_AND2 C447 ( .A(N199), .B(N203), .Z(N204) );
  GTECH_NOT I_39 ( .A(mul_frac_in2_51), .Z(N203) );
  GTECH_AND2 C450 ( .A(N206), .B(m1stg_sngopa[1]), .Z(m1stg_qnan_sng_in1) );
  GTECH_AND2 C451 ( .A(N192), .B(mul_frac_in1_54), .Z(N206) );
  GTECH_AND2 C453 ( .A(N207), .B(m1stg_dblopa[1]), .Z(m1stg_qnan_dbl_in1) );
  GTECH_AND2 C454 ( .A(N192), .B(mul_frac_in1_51), .Z(N207) );
  GTECH_AND2 C456 ( .A(N208), .B(m1stg_sngopa[1]), .Z(m1stg_qnan_sng_in2) );
  GTECH_AND2 C457 ( .A(N199), .B(mul_frac_in2_54), .Z(N208) );
  GTECH_AND2 C459 ( .A(N209), .B(m1stg_dblopa[1]), .Z(m1stg_qnan_dbl_in2) );
  GTECH_AND2 C460 ( .A(N199), .B(mul_frac_in2_51), .Z(N209) );
  GTECH_OR2 C462 ( .A(m1stg_snan_sng_in1), .B(m1stg_snan_dbl_in1), .Z(
        m1stg_snan_in1) );
  GTECH_OR2 C463 ( .A(m1stg_snan_sng_in2), .B(m1stg_snan_dbl_in2), .Z(
        m1stg_snan_in2) );
  GTECH_OR2 C464 ( .A(m1stg_qnan_sng_in1), .B(m1stg_qnan_dbl_in1), .Z(
        m1stg_qnan_in1) );
  GTECH_OR2 C465 ( .A(m1stg_qnan_sng_in2), .B(m1stg_qnan_dbl_in2), .Z(
        m1stg_qnan_in2) );
  GTECH_AND2 C466 ( .A(N211), .B(m1stg_sngopa[2]), .Z(m1stg_nan_sng_in1) );
  GTECH_AND2 C467 ( .A(N192), .B(N210), .Z(N211) );
  GTECH_OR2 C469 ( .A(mul_frac_in1_54), .B(mul_frac_in1_53_32_neq_0), .Z(N210)
         );
  GTECH_AND2 C470 ( .A(N213), .B(m1stg_dblopa[2]), .Z(m1stg_nan_dbl_in1) );
  GTECH_AND2 C471 ( .A(N192), .B(N212), .Z(N213) );
  GTECH_OR2 C473 ( .A(mul_frac_in1_51), .B(mul_frac_in1_50_0_neq_0), .Z(N212)
         );
  GTECH_AND2 C474 ( .A(N215), .B(m1stg_sngopa[2]), .Z(m1stg_nan_sng_in2) );
  GTECH_AND2 C475 ( .A(N199), .B(N214), .Z(N215) );
  GTECH_OR2 C477 ( .A(mul_frac_in2_54), .B(mul_frac_in2_53_32_neq_0), .Z(N214)
         );
  GTECH_AND2 C478 ( .A(N217), .B(m1stg_dblopa[2]), .Z(m1stg_nan_dbl_in2) );
  GTECH_AND2 C479 ( .A(N199), .B(N216), .Z(N217) );
  GTECH_OR2 C481 ( .A(mul_frac_in2_51), .B(mul_frac_in2_50_0_neq_0), .Z(N216)
         );
  GTECH_OR2 C482 ( .A(m1stg_nan_sng_in1), .B(m1stg_nan_dbl_in1), .Z(
        m1stg_nan_in1) );
  GTECH_OR2 C483 ( .A(m1stg_nan_sng_in2), .B(m1stg_nan_dbl_in2), .Z(
        m1stg_nan_in2) );
  GTECH_AND2 C484 ( .A(N220), .B(m1stg_sngopa[2]), .Z(m1stg_inf_sng_in1) );
  GTECH_AND2 C485 ( .A(N218), .B(N219), .Z(N220) );
  GTECH_AND2 C486 ( .A(N192), .B(N193), .Z(N218) );
  GTECH_NOT I_40 ( .A(mul_frac_in1_53_32_neq_0), .Z(N219) );
  GTECH_AND2 C490 ( .A(N223), .B(m1stg_dblopa[2]), .Z(m1stg_inf_dbl_in1) );
  GTECH_AND2 C491 ( .A(N221), .B(N222), .Z(N223) );
  GTECH_AND2 C492 ( .A(N192), .B(N196), .Z(N221) );
  GTECH_NOT I_41 ( .A(mul_frac_in1_50_0_neq_0), .Z(N222) );
  GTECH_AND2 C496 ( .A(N226), .B(m1stg_sngopa[2]), .Z(m1stg_inf_sng_in2) );
  GTECH_AND2 C497 ( .A(N224), .B(N225), .Z(N226) );
  GTECH_AND2 C498 ( .A(N199), .B(N200), .Z(N224) );
  GTECH_NOT I_42 ( .A(mul_frac_in2_53_32_neq_0), .Z(N225) );
  GTECH_AND2 C502 ( .A(N229), .B(m1stg_dblopa[2]), .Z(m1stg_inf_dbl_in2) );
  GTECH_AND2 C503 ( .A(N227), .B(N228), .Z(N229) );
  GTECH_AND2 C504 ( .A(N199), .B(N203), .Z(N227) );
  GTECH_NOT I_43 ( .A(mul_frac_in2_50_0_neq_0), .Z(N228) );
  GTECH_OR2 C508 ( .A(m1stg_inf_sng_in1), .B(m1stg_inf_dbl_in1), .Z(
        m1stg_inf_in1) );
  GTECH_OR2 C509 ( .A(m1stg_inf_sng_in2), .B(m1stg_inf_dbl_in2), .Z(
        m1stg_inf_in2) );
  GTECH_OR2 C510 ( .A(m1stg_inf_in1), .B(m1stg_inf_in2), .Z(m1stg_inf_in) );
  GTECH_AND2 C511 ( .A(N192), .B(m1stg_sngopa[3]), .Z(m1stg_infnan_sng_in1) );
  GTECH_AND2 C513 ( .A(N192), .B(m1stg_dblopa[3]), .Z(m1stg_infnan_dbl_in1) );
  GTECH_AND2 C515 ( .A(N199), .B(m1stg_sngopa[3]), .Z(m1stg_infnan_sng_in2) );
  GTECH_AND2 C517 ( .A(N199), .B(m1stg_dblopa[3]), .Z(m1stg_infnan_dbl_in2) );
  GTECH_OR2 C519 ( .A(m1stg_infnan_sng_in1), .B(m1stg_infnan_dbl_in1), .Z(
        m1stg_infnan_in1) );
  GTECH_OR2 C520 ( .A(m1stg_infnan_sng_in2), .B(m1stg_infnan_dbl_in2), .Z(
        m1stg_infnan_in2) );
  GTECH_OR2 C521 ( .A(m1stg_infnan_in1), .B(m1stg_infnan_in2), .Z(
        m1stg_infnan_in) );
  GTECH_AND2 C522 ( .A(N231), .B(N193), .Z(m1stg_zero_in1) );
  GTECH_AND2 C523 ( .A(mul_exp_in1_exp_eq_0), .B(N230), .Z(N231) );
  GTECH_NOT I_44 ( .A(mul_frac_in1_53_0_neq_0), .Z(N230) );
  GTECH_AND2 C526 ( .A(N233), .B(N200), .Z(m1stg_zero_in2) );
  GTECH_AND2 C527 ( .A(mul_exp_in2_exp_eq_0), .B(N232), .Z(N233) );
  GTECH_NOT I_45 ( .A(mul_frac_in2_53_0_neq_0), .Z(N232) );
  GTECH_OR2 C530 ( .A(m1stg_zero_in1), .B(m1stg_zero_in2), .Z(m1stg_zero_in)
         );
  GTECH_AND2 C531 ( .A(m6stg_stepa), .B(N234), .Z(m1stg_step) );
  GTECH_NOT I_46 ( .A(m1stg_mul), .Z(N234) );
  GTECH_NOT I_47 ( .A(reset), .Z(N0) );
  GTECH_OR2 C534 ( .A(N237), .B(N240), .Z(m1stg_op_in[7]) );
  GTECH_AND2 C535 ( .A(N235), .B(N236), .Z(N237) );
  GTECH_AND2 C536 ( .A(m1stg_step), .B(N0), .Z(N235) );
  GTECH_AND2 C537 ( .A(inq_op[7]), .B(inq_mul), .Z(N236) );
  GTECH_AND2 C538 ( .A(N239), .B(m1stg_op[7]), .Z(N240) );
  GTECH_AND2 C539 ( .A(N238), .B(N0), .Z(N239) );
  GTECH_NOT I_48 ( .A(m6stg_step), .Z(N238) );
  GTECH_OR2 C541 ( .A(N243), .B(N246), .Z(m1stg_op_in[6]) );
  GTECH_AND2 C542 ( .A(N241), .B(N242), .Z(N243) );
  GTECH_AND2 C543 ( .A(m1stg_step), .B(N0), .Z(N241) );
  GTECH_AND2 C544 ( .A(inq_op[6]), .B(inq_mul), .Z(N242) );
  GTECH_AND2 C545 ( .A(N245), .B(m1stg_op[6]), .Z(N246) );
  GTECH_AND2 C546 ( .A(N244), .B(N0), .Z(N245) );
  GTECH_NOT I_49 ( .A(m6stg_step), .Z(N244) );
  GTECH_OR2 C548 ( .A(N249), .B(N252), .Z(m1stg_op_in[5]) );
  GTECH_AND2 C549 ( .A(N247), .B(N248), .Z(N249) );
  GTECH_AND2 C550 ( .A(m1stg_step), .B(N0), .Z(N247) );
  GTECH_AND2 C551 ( .A(inq_op[5]), .B(inq_mul), .Z(N248) );
  GTECH_AND2 C552 ( .A(N251), .B(m1stg_op[5]), .Z(N252) );
  GTECH_AND2 C553 ( .A(N250), .B(N0), .Z(N251) );
  GTECH_NOT I_50 ( .A(m6stg_step), .Z(N250) );
  GTECH_OR2 C555 ( .A(N255), .B(N258), .Z(m1stg_op_in[4]) );
  GTECH_AND2 C556 ( .A(N253), .B(N254), .Z(N255) );
  GTECH_AND2 C557 ( .A(m1stg_step), .B(N0), .Z(N253) );
  GTECH_AND2 C558 ( .A(inq_op[4]), .B(inq_mul), .Z(N254) );
  GTECH_AND2 C559 ( .A(N257), .B(m1stg_op[4]), .Z(N258) );
  GTECH_AND2 C560 ( .A(N256), .B(N0), .Z(N257) );
  GTECH_NOT I_51 ( .A(m6stg_step), .Z(N256) );
  GTECH_OR2 C562 ( .A(N261), .B(N264), .Z(m1stg_op_in[3]) );
  GTECH_AND2 C563 ( .A(N259), .B(N260), .Z(N261) );
  GTECH_AND2 C564 ( .A(m1stg_step), .B(N0), .Z(N259) );
  GTECH_AND2 C565 ( .A(inq_op[3]), .B(inq_mul), .Z(N260) );
  GTECH_AND2 C566 ( .A(N263), .B(m1stg_op[3]), .Z(N264) );
  GTECH_AND2 C567 ( .A(N262), .B(N0), .Z(N263) );
  GTECH_NOT I_52 ( .A(m6stg_step), .Z(N262) );
  GTECH_OR2 C569 ( .A(N267), .B(N270), .Z(m1stg_op_in[2]) );
  GTECH_AND2 C570 ( .A(N265), .B(N266), .Z(N267) );
  GTECH_AND2 C571 ( .A(m1stg_step), .B(N0), .Z(N265) );
  GTECH_AND2 C572 ( .A(inq_op[2]), .B(inq_mul), .Z(N266) );
  GTECH_AND2 C573 ( .A(N269), .B(m1stg_op[2]), .Z(N270) );
  GTECH_AND2 C574 ( .A(N268), .B(N0), .Z(N269) );
  GTECH_NOT I_53 ( .A(m6stg_step), .Z(N268) );
  GTECH_OR2 C576 ( .A(N273), .B(N276), .Z(m1stg_op_in[1]) );
  GTECH_AND2 C577 ( .A(N271), .B(N272), .Z(N273) );
  GTECH_AND2 C578 ( .A(m1stg_step), .B(N0), .Z(N271) );
  GTECH_AND2 C579 ( .A(inq_op[1]), .B(inq_mul), .Z(N272) );
  GTECH_AND2 C580 ( .A(N275), .B(m1stg_op[1]), .Z(N276) );
  GTECH_AND2 C581 ( .A(N274), .B(N0), .Z(N275) );
  GTECH_NOT I_54 ( .A(m6stg_step), .Z(N274) );
  GTECH_OR2 C583 ( .A(N279), .B(N282), .Z(m1stg_op_in[0]) );
  GTECH_AND2 C584 ( .A(N277), .B(N278), .Z(N279) );
  GTECH_AND2 C585 ( .A(m1stg_step), .B(N0), .Z(N277) );
  GTECH_AND2 C586 ( .A(inq_op[0]), .B(inq_mul), .Z(N278) );
  GTECH_AND2 C587 ( .A(N281), .B(m1stg_op[0]), .Z(N282) );
  GTECH_AND2 C588 ( .A(N280), .B(N0), .Z(N281) );
  GTECH_NOT I_55 ( .A(m6stg_step), .Z(N280) );
  GTECH_NOT I_56 ( .A(reset), .Z(N1) );
  GTECH_OR2 C591 ( .A(N284), .B(N287), .Z(m1stg_mul_in) );
  GTECH_AND2 C592 ( .A(N283), .B(inq_mul), .Z(N284) );
  GTECH_AND2 C593 ( .A(m1stg_step), .B(N1), .Z(N283) );
  GTECH_AND2 C594 ( .A(N286), .B(m1stg_mul), .Z(N287) );
  GTECH_AND2 C595 ( .A(N285), .B(N1), .Z(N286) );
  GTECH_NOT I_57 ( .A(m6stg_step), .Z(N285) );
  GTECH_NOT I_58 ( .A(inq_op[1]), .Z(m1stg_dblop_inv_in) );
  GTECH_OR2 C598 ( .A(N288), .B(N109), .Z(m1stg_fmul) );
  GTECH_OR2 C599 ( .A(N93), .B(N101), .Z(N288) );
  GTECH_OR2 C600 ( .A(N70), .B(N78), .Z(m1stg_opdec[3]) );
  GTECH_NOT I_59 ( .A(reset), .Z(N2) );
  GTECH_OR2 C602 ( .A(N290), .B(N293), .Z(m6stg_fmul_in) );
  GTECH_AND2 C603 ( .A(N289), .B(m5stg_opdec[4]), .Z(N290) );
  GTECH_AND2 C604 ( .A(m6stg_stepa), .B(N2), .Z(N289) );
  GTECH_AND2 C605 ( .A(N292), .B(m6stg_opdec[4]), .Z(N293) );
  GTECH_AND2 C606 ( .A(N291), .B(N2), .Z(N292) );
  GTECH_NOT I_60 ( .A(m6stg_stepa), .Z(N291) );
  GTECH_OR2 C608 ( .A(N294), .B(N295), .Z(m6stg_id_in[9]) );
  GTECH_AND2 C609 ( .A(m6stg_stepa), .B(N9), .Z(N294) );
  GTECH_AND2 C610 ( .A(N291), .B(m6stg_id[9]), .Z(N295) );
  GTECH_OR2 C612 ( .A(N296), .B(N297), .Z(m6stg_id_in[8]) );
  GTECH_AND2 C613 ( .A(m6stg_stepa), .B(N14), .Z(N296) );
  GTECH_AND2 C614 ( .A(N291), .B(m6stg_id[8]), .Z(N297) );
  GTECH_OR2 C616 ( .A(N298), .B(N299), .Z(m6stg_id_in[7]) );
  GTECH_AND2 C617 ( .A(m6stg_stepa), .B(N18), .Z(N298) );
  GTECH_AND2 C618 ( .A(N291), .B(m6stg_id[7]), .Z(N299) );
  GTECH_OR2 C620 ( .A(N300), .B(N301), .Z(m6stg_id_in[6]) );
  GTECH_AND2 C621 ( .A(m6stg_stepa), .B(N21), .Z(N300) );
  GTECH_AND2 C622 ( .A(N291), .B(m6stg_id[6]), .Z(N301) );
  GTECH_OR2 C624 ( .A(N302), .B(N303), .Z(m6stg_id_in[5]) );
  GTECH_AND2 C625 ( .A(m6stg_stepa), .B(N24), .Z(N302) );
  GTECH_AND2 C626 ( .A(N291), .B(m6stg_id[5]), .Z(N303) );
  GTECH_OR2 C628 ( .A(N304), .B(N305), .Z(m6stg_id_in[4]) );
  GTECH_AND2 C629 ( .A(m6stg_stepa), .B(N27), .Z(N304) );
  GTECH_AND2 C630 ( .A(N291), .B(m6stg_id[4]), .Z(N305) );
  GTECH_OR2 C632 ( .A(N306), .B(N307), .Z(m6stg_id_in[3]) );
  GTECH_AND2 C633 ( .A(m6stg_stepa), .B(N30), .Z(N306) );
  GTECH_AND2 C634 ( .A(N291), .B(m6stg_id[3]), .Z(N307) );
  GTECH_OR2 C636 ( .A(N308), .B(N309), .Z(m6stg_id_in[2]) );
  GTECH_AND2 C637 ( .A(m6stg_stepa), .B(N33), .Z(N308) );
  GTECH_AND2 C638 ( .A(N291), .B(m6stg_id[2]), .Z(N309) );
  GTECH_OR2 C640 ( .A(N310), .B(N311), .Z(m6stg_id_in[1]) );
  GTECH_AND2 C641 ( .A(m6stg_stepa), .B(m5stg_id[1]), .Z(N310) );
  GTECH_AND2 C642 ( .A(N291), .B(m6stg_id[1]), .Z(N311) );
  GTECH_OR2 C644 ( .A(N312), .B(N313), .Z(m6stg_id_in[0]) );
  GTECH_AND2 C645 ( .A(m6stg_stepa), .B(m5stg_id[0]), .Z(N312) );
  GTECH_AND2 C646 ( .A(N291), .B(m6stg_id[0]), .Z(N313) );
  GTECH_AND2 C648 ( .A(m6stg_opdec[4]), .B(N314), .Z(m6stg_hold) );
  GTECH_NOT I_61 ( .A(mul_dest_rdy), .Z(N314) );
  GTECH_AND2 C650 ( .A(m6stg_opdec[4]), .B(N315), .Z(m6stg_holda) );
  GTECH_NOT I_62 ( .A(mul_dest_rdya), .Z(N315) );
  GTECH_NOT I_63 ( .A(m6stg_hold), .Z(m6stg_step) );
  GTECH_NOT I_64 ( .A(m6stg_holda), .Z(m6stg_stepa) );
  GTECH_OR2 C654 ( .A(N321), .B(m6stg_opdec[4]), .Z(mul_pipe_active_in) );
  GTECH_OR2 C655 ( .A(N320), .B(m5stg_opdec[4]), .Z(N321) );
  GTECH_OR2 C656 ( .A(N319), .B(m4stg_opdec[4]), .Z(N320) );
  GTECH_OR2 C657 ( .A(N318), .B(m3stg_opdec[4]), .Z(N319) );
  GTECH_OR2 C658 ( .A(N317), .B(m3bstg_opdec[4]), .Z(N318) );
  GTECH_OR2 C659 ( .A(N316), .B(m3astg_opdec[4]), .Z(N317) );
  GTECH_OR2 C660 ( .A(m1stg_fmul), .B(m2stg_opdec[4]), .Z(N316) );
  GTECH_NOT I_65 ( .A(m1stg_infnan_in), .Z(m1stg_of_mask) );
  GTECH_NOT I_66 ( .A(m2stg_snan_in2), .Z(N3) );
  GTECH_AND2 C663 ( .A(N334), .B(N336), .Z(m2stg_sign) );
  GTECH_XOR2 C664 ( .A(N326), .B(N333), .Z(N334) );
  GTECH_AND2 C665 ( .A(N322), .B(N325), .Z(N326) );
  GTECH_AND2 C666 ( .A(m2stg_sign1), .B(N3), .Z(N322) );
  GTECH_NOT I_67 ( .A(N324), .Z(N325) );
  GTECH_AND2 C668 ( .A(m2stg_qnan_in2), .B(N323), .Z(N324) );
  GTECH_NOT I_68 ( .A(m2stg_snan_in1), .Z(N323) );
  GTECH_AND2 C670 ( .A(N329), .B(N332), .Z(N333) );
  GTECH_AND2 C671 ( .A(m2stg_sign2), .B(N328), .Z(N329) );
  GTECH_NOT I_69 ( .A(N327), .Z(N328) );
  GTECH_AND2 C673 ( .A(m2stg_snan_in1), .B(N3), .Z(N327) );
  GTECH_NOT I_70 ( .A(N331), .Z(N332) );
  GTECH_AND2 C675 ( .A(m2stg_qnan_in1), .B(N330), .Z(N331) );
  GTECH_NOT I_71 ( .A(m2stg_nan_in2), .Z(N330) );
  GTECH_NOT I_72 ( .A(N335), .Z(N336) );
  GTECH_AND2 C678 ( .A(m2stg_inf_in), .B(m2stg_zero_in), .Z(N335) );
  GTECH_OR2 C679 ( .A(N339), .B(N340), .Z(m2stg_nv) );
  GTECH_OR2 C680 ( .A(N337), .B(N338), .Z(N339) );
  GTECH_OR2 C681 ( .A(m2stg_snan_in1), .B(m2stg_snan_in2), .Z(N337) );
  GTECH_AND2 C682 ( .A(m2stg_zero_in1), .B(m2stg_inf_in2), .Z(N338) );
  GTECH_AND2 C683 ( .A(m2stg_inf_in1), .B(m2stg_zero_in2), .Z(N340) );
  GTECH_NOT I_73 ( .A(m5stg_exp[12]), .Z(N4) );
  GTECH_OR2 C685 ( .A(N354), .B(N368), .Z(m5stg_in_of) );
  GTECH_AND2 C686 ( .A(N353), .B(m5stg_of_mask), .Z(N354) );
  GTECH_AND2 C687 ( .A(N341), .B(N352), .Z(N353) );
  GTECH_AND2 C688 ( .A(N4), .B(m5stg_fmuld), .Z(N341) );
  GTECH_OR2 C689 ( .A(m5stg_exp[11]), .B(N351), .Z(N352) );
  GTECH_AND2 C690 ( .A(N350), .B(m5stg_exp[0]), .Z(N351) );
  GTECH_AND2 C691 ( .A(N349), .B(m5stg_exp[1]), .Z(N350) );
  GTECH_AND2 C692 ( .A(N348), .B(m5stg_exp[2]), .Z(N349) );
  GTECH_AND2 C693 ( .A(N347), .B(m5stg_exp[3]), .Z(N348) );
  GTECH_AND2 C694 ( .A(N346), .B(m5stg_exp[4]), .Z(N347) );
  GTECH_AND2 C695 ( .A(N345), .B(m5stg_exp[5]), .Z(N346) );
  GTECH_AND2 C696 ( .A(N344), .B(m5stg_exp[6]), .Z(N345) );
  GTECH_AND2 C697 ( .A(N343), .B(m5stg_exp[7]), .Z(N344) );
  GTECH_AND2 C698 ( .A(N342), .B(m5stg_exp[8]), .Z(N343) );
  GTECH_AND2 C699 ( .A(m5stg_exp[10]), .B(m5stg_exp[9]), .Z(N342) );
  GTECH_AND2 C700 ( .A(N367), .B(m5stg_of_mask), .Z(N368) );
  GTECH_AND2 C701 ( .A(N355), .B(N366), .Z(N367) );
  GTECH_AND2 C702 ( .A(N4), .B(m5stg_fmuls), .Z(N355) );
  GTECH_OR2 C703 ( .A(N358), .B(N365), .Z(N366) );
  GTECH_OR2 C704 ( .A(N357), .B(m5stg_exp[8]), .Z(N358) );
  GTECH_OR2 C705 ( .A(N356), .B(m5stg_exp[9]), .Z(N357) );
  GTECH_OR2 C706 ( .A(m5stg_exp[11]), .B(m5stg_exp[10]), .Z(N356) );
  GTECH_AND2 C707 ( .A(N364), .B(m5stg_exp[0]), .Z(N365) );
  GTECH_AND2 C708 ( .A(N363), .B(m5stg_exp[1]), .Z(N364) );
  GTECH_AND2 C709 ( .A(N362), .B(m5stg_exp[2]), .Z(N363) );
  GTECH_AND2 C710 ( .A(N361), .B(m5stg_exp[3]), .Z(N362) );
  GTECH_AND2 C711 ( .A(N360), .B(m5stg_exp[4]), .Z(N361) );
  GTECH_AND2 C712 ( .A(N359), .B(m5stg_exp[5]), .Z(N360) );
  GTECH_AND2 C713 ( .A(m5stg_exp[7]), .B(m5stg_exp[6]), .Z(N359) );
  GTECH_OR2 C714 ( .A(N381), .B(N391), .Z(mul_of_out_tmp1_in) );
  GTECH_AND2 C715 ( .A(N380), .B(m5stg_of_mask), .Z(N381) );
  GTECH_AND2 C716 ( .A(N379), .B(m5stg_rndup), .Z(N380) );
  GTECH_AND2 C717 ( .A(N369), .B(N378), .Z(N379) );
  GTECH_AND2 C718 ( .A(N4), .B(m5stg_fmuld), .Z(N369) );
  GTECH_AND2 C719 ( .A(N377), .B(m5stg_exp[1]), .Z(N378) );
  GTECH_AND2 C720 ( .A(N376), .B(m5stg_exp[2]), .Z(N377) );
  GTECH_AND2 C721 ( .A(N375), .B(m5stg_exp[3]), .Z(N376) );
  GTECH_AND2 C722 ( .A(N374), .B(m5stg_exp[4]), .Z(N375) );
  GTECH_AND2 C723 ( .A(N373), .B(m5stg_exp[5]), .Z(N374) );
  GTECH_AND2 C724 ( .A(N372), .B(m5stg_exp[6]), .Z(N373) );
  GTECH_AND2 C725 ( .A(N371), .B(m5stg_exp[7]), .Z(N372) );
  GTECH_AND2 C726 ( .A(N370), .B(m5stg_exp[8]), .Z(N371) );
  GTECH_AND2 C727 ( .A(m5stg_exp[10]), .B(m5stg_exp[9]), .Z(N370) );
  GTECH_AND2 C728 ( .A(N390), .B(m5stg_of_mask), .Z(N391) );
  GTECH_AND2 C729 ( .A(N389), .B(m5stg_rndup), .Z(N390) );
  GTECH_AND2 C730 ( .A(N382), .B(N388), .Z(N389) );
  GTECH_AND2 C731 ( .A(N4), .B(m5stg_fmuls), .Z(N382) );
  GTECH_AND2 C732 ( .A(N387), .B(m5stg_exp[1]), .Z(N388) );
  GTECH_AND2 C733 ( .A(N386), .B(m5stg_exp[2]), .Z(N387) );
  GTECH_AND2 C734 ( .A(N385), .B(m5stg_exp[3]), .Z(N386) );
  GTECH_AND2 C735 ( .A(N384), .B(m5stg_exp[4]), .Z(N385) );
  GTECH_AND2 C736 ( .A(N383), .B(m5stg_exp[5]), .Z(N384) );
  GTECH_AND2 C737 ( .A(m5stg_exp[7]), .B(m5stg_exp[6]), .Z(N383) );
  GTECH_OR2 C738 ( .A(mul_of_out_tmp2), .B(N392), .Z(mul_exc_out[3]) );
  GTECH_AND2 C739 ( .A(mul_of_out_tmp1), .B(mul_of_out_cout), .Z(N392) );
  GTECH_AND2 C740 ( .A(N405), .B(m5stg_frac_neq_0), .Z(mul_uf_out_in) );
  GTECH_OR2 C741 ( .A(m5stg_exp[12]), .B(N404), .Z(N405) );
  GTECH_NOT I_74 ( .A(N403), .Z(N404) );
  GTECH_OR2 C743 ( .A(N402), .B(m5stg_exp[0]), .Z(N403) );
  GTECH_OR2 C744 ( .A(N401), .B(m5stg_exp[1]), .Z(N402) );
  GTECH_OR2 C745 ( .A(N400), .B(m5stg_exp[2]), .Z(N401) );
  GTECH_OR2 C746 ( .A(N399), .B(m5stg_exp[3]), .Z(N400) );
  GTECH_OR2 C747 ( .A(N398), .B(m5stg_exp[4]), .Z(N399) );
  GTECH_OR2 C748 ( .A(N397), .B(m5stg_exp[5]), .Z(N398) );
  GTECH_OR2 C749 ( .A(N396), .B(m5stg_exp[6]), .Z(N397) );
  GTECH_OR2 C750 ( .A(N395), .B(m5stg_exp[7]), .Z(N396) );
  GTECH_OR2 C751 ( .A(N394), .B(m5stg_exp[8]), .Z(N395) );
  GTECH_OR2 C752 ( .A(N393), .B(m5stg_exp[9]), .Z(N394) );
  GTECH_OR2 C753 ( .A(m5stg_exp[11]), .B(m5stg_exp[10]), .Z(N393) );
  GTECH_OR2 C754 ( .A(N406), .B(N407), .Z(mul_nx_out_in) );
  GTECH_AND2 C755 ( .A(m5stg_fmuld), .B(m5stg_frac_dbl_nx), .Z(N406) );
  GTECH_AND2 C756 ( .A(m5stg_fmuls), .B(m5stg_frac_sng_nx), .Z(N407) );
  GTECH_OR2 C757 ( .A(mul_nx_out), .B(mul_exc_out[3]), .Z(mul_exc_out_0) );
  GTECH_AND2 C758 ( .A(m1stg_norm_dbl_in1), .B(N415), .Z(m2stg_frac1_dbl_norm)
         );
  GTECH_OR2 C759 ( .A(N412), .B(N414), .Z(N415) );
  GTECH_OR2 C760 ( .A(N409), .B(N411), .Z(N412) );
  GTECH_NOT I_75 ( .A(N408), .Z(N409) );
  GTECH_OR2 C762 ( .A(m1stg_infnan_dbl_in1), .B(m1stg_infnan_dbl_in2), .Z(N408) );
  GTECH_AND2 C763 ( .A(m1stg_snan_dbl_in1), .B(N410), .Z(N411) );
  GTECH_NOT I_76 ( .A(m1stg_snan_dbl_in2), .Z(N410) );
  GTECH_AND2 C765 ( .A(m1stg_qnan_dbl_in1), .B(N413), .Z(N414) );
  GTECH_NOT I_77 ( .A(m1stg_nan_dbl_in2), .Z(N413) );
  GTECH_AND2 C767 ( .A(m1stg_denorm_dbl_in1), .B(N417), .Z(
        m2stg_frac1_dbl_dnrm) );
  GTECH_NOT I_78 ( .A(N416), .Z(N417) );
  GTECH_OR2 C769 ( .A(m1stg_infnan_dbl_in1), .B(m1stg_infnan_dbl_in2), .Z(N416) );
  GTECH_AND2 C770 ( .A(m1stg_norm_sng_in1), .B(N425), .Z(m2stg_frac1_sng_norm)
         );
  GTECH_OR2 C771 ( .A(N422), .B(N424), .Z(N425) );
  GTECH_OR2 C772 ( .A(N419), .B(N421), .Z(N422) );
  GTECH_NOT I_79 ( .A(N418), .Z(N419) );
  GTECH_OR2 C774 ( .A(m1stg_infnan_sng_in1), .B(m1stg_infnan_sng_in2), .Z(N418) );
  GTECH_AND2 C775 ( .A(m1stg_snan_sng_in1), .B(N420), .Z(N421) );
  GTECH_NOT I_80 ( .A(m1stg_snan_sng_in2), .Z(N420) );
  GTECH_AND2 C777 ( .A(m1stg_qnan_sng_in1), .B(N423), .Z(N424) );
  GTECH_NOT I_81 ( .A(m1stg_nan_sng_in2), .Z(N423) );
  GTECH_AND2 C779 ( .A(m1stg_denorm_sng_in1), .B(N427), .Z(
        m2stg_frac1_sng_dnrm) );
  GTECH_NOT I_82 ( .A(N426), .Z(N427) );
  GTECH_OR2 C781 ( .A(m1stg_infnan_sng_in1), .B(m1stg_infnan_sng_in2), .Z(N426) );
  GTECH_OR2 C782 ( .A(N432), .B(N434), .Z(m2stg_frac1_inf) );
  GTECH_OR2 C783 ( .A(N431), .B(m1stg_snan_in2), .Z(N432) );
  GTECH_AND2 C784 ( .A(N429), .B(N430), .Z(N431) );
  GTECH_AND2 C785 ( .A(m1stg_inf_in), .B(N428), .Z(N429) );
  GTECH_NOT I_83 ( .A(m1stg_nan_in1), .Z(N428) );
  GTECH_NOT I_84 ( .A(m1stg_nan_in2), .Z(N430) );
  GTECH_AND2 C788 ( .A(m1stg_qnan_in2), .B(N433), .Z(N434) );
  GTECH_NOT I_85 ( .A(m1stg_snan_in1), .Z(N433) );
  GTECH_AND2 C790 ( .A(m1stg_norm_dbl_in2), .B(N440), .Z(m2stg_frac2_dbl_norm)
         );
  GTECH_OR2 C791 ( .A(N437), .B(N439), .Z(N440) );
  GTECH_OR2 C792 ( .A(N436), .B(m1stg_snan_dbl_in2), .Z(N437) );
  GTECH_NOT I_86 ( .A(N435), .Z(N436) );
  GTECH_OR2 C794 ( .A(m1stg_infnan_dbl_in1), .B(m1stg_infnan_dbl_in2), .Z(N435) );
  GTECH_AND2 C795 ( .A(m1stg_qnan_dbl_in2), .B(N438), .Z(N439) );
  GTECH_NOT I_87 ( .A(m1stg_snan_dbl_in1), .Z(N438) );
  GTECH_AND2 C797 ( .A(m1stg_denorm_dbl_in2), .B(N442), .Z(
        m2stg_frac2_dbl_dnrm) );
  GTECH_NOT I_88 ( .A(N441), .Z(N442) );
  GTECH_OR2 C799 ( .A(m1stg_infnan_dbl_in1), .B(m1stg_infnan_dbl_in2), .Z(N441) );
  GTECH_AND2 C800 ( .A(m1stg_norm_sng_in2), .B(N448), .Z(m2stg_frac2_sng_norm)
         );
  GTECH_OR2 C801 ( .A(N445), .B(N447), .Z(N448) );
  GTECH_OR2 C802 ( .A(N444), .B(m1stg_snan_sng_in2), .Z(N445) );
  GTECH_NOT I_89 ( .A(N443), .Z(N444) );
  GTECH_OR2 C804 ( .A(m1stg_infnan_sng_in1), .B(m1stg_infnan_sng_in2), .Z(N443) );
  GTECH_AND2 C805 ( .A(m1stg_qnan_sng_in2), .B(N446), .Z(N447) );
  GTECH_NOT I_90 ( .A(m1stg_snan_sng_in1), .Z(N446) );
  GTECH_AND2 C807 ( .A(m1stg_denorm_sng_in2), .B(N450), .Z(
        m2stg_frac2_sng_dnrm) );
  GTECH_NOT I_91 ( .A(N449), .Z(N450) );
  GTECH_OR2 C809 ( .A(m1stg_infnan_sng_in1), .B(m1stg_infnan_sng_in2), .Z(N449) );
  GTECH_NOT I_92 ( .A(m1stg_nan_in2), .Z(N5) );
  GTECH_OR2 C811 ( .A(N455), .B(N456), .Z(m2stg_frac2_inf) );
  GTECH_OR2 C812 ( .A(N452), .B(N454), .Z(N455) );
  GTECH_AND2 C813 ( .A(N451), .B(N5), .Z(N452) );
  GTECH_AND2 C814 ( .A(m1stg_inf_in), .B(N428), .Z(N451) );
  GTECH_AND2 C816 ( .A(m1stg_snan_in1), .B(N453), .Z(N454) );
  GTECH_NOT I_93 ( .A(m1stg_snan_in2), .Z(N453) );
  GTECH_AND2 C818 ( .A(m1stg_qnan_in1), .B(N5), .Z(N456) );
  GTECH_OR2 C819 ( .A(N457), .B(N458), .Z(m1stg_inf_zero_in) );
  GTECH_AND2 C820 ( .A(m1stg_inf_in1), .B(m1stg_zero_in2), .Z(N457) );
  GTECH_AND2 C821 ( .A(m1stg_zero_in1), .B(m1stg_inf_in2), .Z(N458) );
  GTECH_AND2 C822 ( .A(N461), .B(m1stg_opdec[3]), .Z(m1stg_inf_zero_in_dbl) );
  GTECH_OR2 C823 ( .A(N459), .B(N460), .Z(N461) );
  GTECH_AND2 C824 ( .A(m1stg_inf_in1), .B(m1stg_zero_in2), .Z(N459) );
  GTECH_AND2 C825 ( .A(m1stg_zero_in1), .B(m1stg_inf_in2), .Z(N460) );
  GTECH_AND2 C826 ( .A(N463), .B(m1stg_ld0_1[5]), .Z(m2stg_ld0_1_in[5]) );
  GTECH_AND2 C827 ( .A(m1stg_denorm_in1), .B(N462), .Z(N463) );
  GTECH_NOT I_94 ( .A(m1stg_infnan_in), .Z(N462) );
  GTECH_AND2 C829 ( .A(N464), .B(m1stg_ld0_1[4]), .Z(m2stg_ld0_1_in[4]) );
  GTECH_AND2 C830 ( .A(m1stg_denorm_in1), .B(N462), .Z(N464) );
  GTECH_AND2 C832 ( .A(N465), .B(m1stg_ld0_1[3]), .Z(m2stg_ld0_1_in[3]) );
  GTECH_AND2 C833 ( .A(m1stg_denorm_in1), .B(N462), .Z(N465) );
  GTECH_AND2 C835 ( .A(N466), .B(m1stg_ld0_1[2]), .Z(m2stg_ld0_1_in[2]) );
  GTECH_AND2 C836 ( .A(m1stg_denorm_in1), .B(N462), .Z(N466) );
  GTECH_AND2 C838 ( .A(N467), .B(m1stg_ld0_1[1]), .Z(m2stg_ld0_1_in[1]) );
  GTECH_AND2 C839 ( .A(m1stg_denorm_in1), .B(N462), .Z(N467) );
  GTECH_AND2 C841 ( .A(N468), .B(m1stg_ld0_1[0]), .Z(m2stg_ld0_1_in[0]) );
  GTECH_AND2 C842 ( .A(m1stg_denorm_in1), .B(N462), .Z(N468) );
  GTECH_AND2 C844 ( .A(N469), .B(m1stg_ld0_2[5]), .Z(m2stg_ld0_2_in[5]) );
  GTECH_AND2 C845 ( .A(m1stg_denorm_in2), .B(N462), .Z(N469) );
  GTECH_AND2 C847 ( .A(N470), .B(m1stg_ld0_2[4]), .Z(m2stg_ld0_2_in[4]) );
  GTECH_AND2 C848 ( .A(m1stg_denorm_in2), .B(N462), .Z(N470) );
  GTECH_AND2 C850 ( .A(N471), .B(m1stg_ld0_2[3]), .Z(m2stg_ld0_2_in[3]) );
  GTECH_AND2 C851 ( .A(m1stg_denorm_in2), .B(N462), .Z(N471) );
  GTECH_AND2 C853 ( .A(N472), .B(m1stg_ld0_2[2]), .Z(m2stg_ld0_2_in[2]) );
  GTECH_AND2 C854 ( .A(m1stg_denorm_in2), .B(N462), .Z(N472) );
  GTECH_AND2 C856 ( .A(N473), .B(m1stg_ld0_2[1]), .Z(m2stg_ld0_2_in[1]) );
  GTECH_AND2 C857 ( .A(m1stg_denorm_in2), .B(N462), .Z(N473) );
  GTECH_AND2 C859 ( .A(N474), .B(m1stg_ld0_2[0]), .Z(m2stg_ld0_2_in[0]) );
  GTECH_AND2 C860 ( .A(m1stg_denorm_in2), .B(N462), .Z(N474) );
  GTECH_AND2 C862 ( .A(N462), .B(N475), .Z(m2stg_exp_expadd) );
  GTECH_NOT I_95 ( .A(m1stg_zero_in), .Z(N475) );
  GTECH_AND2 C865 ( .A(N44), .B(m1stg_infnan_in), .Z(m2stg_exp_0bff) );
  GTECH_AND2 C866 ( .A(N53), .B(m1stg_infnan_in), .Z(m2stg_exp_017f) );
  GTECH_AND2 C867 ( .A(N62), .B(m1stg_infnan_in), .Z(m2stg_exp_04ff) );
  GTECH_AND2 C868 ( .A(m1stg_zero_in), .B(N462), .Z(m2stg_exp_zero) );
  GTECH_NOT I_96 ( .A(m2stg_ld0[6]), .Z(m2stg_ld0_inv[6]) );
  GTECH_NOT I_97 ( .A(m2stg_ld0[5]), .Z(m2stg_ld0_inv[5]) );
  GTECH_NOT I_98 ( .A(m2stg_ld0[4]), .Z(m2stg_ld0_inv[4]) );
  GTECH_NOT I_99 ( .A(m2stg_ld0[3]), .Z(m2stg_ld0_inv[3]) );
  GTECH_NOT I_100 ( .A(m2stg_ld0[2]), .Z(m2stg_ld0_inv[2]) );
  GTECH_NOT I_101 ( .A(m2stg_ld0[1]), .Z(m2stg_ld0_inv[1]) );
  GTECH_NOT I_102 ( .A(m2stg_ld0[0]), .Z(m2stg_ld0_inv[0]) );
  GTECH_OR2 C877 ( .A(N487), .B(m3stg_exp[12]), .Z(m3stg_exp_lte_0) );
  GTECH_NOT I_103 ( .A(N486), .Z(N487) );
  GTECH_OR2 C879 ( .A(N485), .B(m3stg_exp[0]), .Z(N486) );
  GTECH_OR2 C880 ( .A(N484), .B(m3stg_exp[1]), .Z(N485) );
  GTECH_OR2 C881 ( .A(N483), .B(m3stg_exp[2]), .Z(N484) );
  GTECH_OR2 C882 ( .A(N482), .B(m3stg_exp[3]), .Z(N483) );
  GTECH_OR2 C883 ( .A(N481), .B(m3stg_exp[4]), .Z(N482) );
  GTECH_OR2 C884 ( .A(N480), .B(m3stg_exp[5]), .Z(N481) );
  GTECH_OR2 C885 ( .A(N479), .B(m3stg_exp[6]), .Z(N480) );
  GTECH_OR2 C886 ( .A(N478), .B(m3stg_exp[7]), .Z(N479) );
  GTECH_OR2 C887 ( .A(N477), .B(m3stg_exp[8]), .Z(N478) );
  GTECH_OR2 C888 ( .A(N476), .B(m3stg_exp[9]), .Z(N477) );
  GTECH_OR2 C889 ( .A(m3stg_exp[11]), .B(m3stg_exp[10]), .Z(N476) );
  GTECH_AND2 C890 ( .A(N488), .B(m3stg_exp_lte_0), .Z(m4stg_right_shift_in) );
  GTECH_NOT I_104 ( .A(m3stg_expadd_lte_0_inv), .Z(N488) );
  GTECH_AND2 C892 ( .A(N498), .B(m3stg_exp[12]), .Z(m3stg_exp_lt_neg57) );
  GTECH_OR2 C893 ( .A(N494), .B(N497), .Z(N498) );
  GTECH_NOT I_105 ( .A(N493), .Z(N494) );
  GTECH_AND2 C895 ( .A(N492), .B(m3stg_exp[6]), .Z(N493) );
  GTECH_AND2 C896 ( .A(N491), .B(m3stg_exp[7]), .Z(N492) );
  GTECH_AND2 C897 ( .A(N490), .B(m3stg_exp[8]), .Z(N491) );
  GTECH_AND2 C898 ( .A(N489), .B(m3stg_exp[9]), .Z(N490) );
  GTECH_AND2 C899 ( .A(m3stg_exp[11]), .B(m3stg_exp[10]), .Z(N489) );
  GTECH_NOT I_106 ( .A(N496), .Z(N497) );
  GTECH_OR2 C901 ( .A(N495), .B(m3stg_exp[3]), .Z(N496) );
  GTECH_OR2 C902 ( .A(m3stg_exp[5]), .B(m3stg_exp[4]), .Z(N495) );
  GTECH_AND2 C904 ( .A(N488), .B(m3stg_exp_lte_0), .Z(N6) );
  GTECH_OR2 C905 ( .A(N507), .B(N509), .Z(m4stg_sh_cnt_in[5]) );
  GTECH_OR2 C906 ( .A(N503), .B(N506), .Z(N507) );
  GTECH_OR2 C907 ( .A(N501), .B(N502), .Z(N503) );
  GTECH_AND2 C908 ( .A(N500), .B(m3stg_exp_minus1[5]), .Z(N501) );
  GTECH_AND2 C909 ( .A(N488), .B(N499), .Z(N500) );
  GTECH_NOT I_107 ( .A(m3stg_exp_lte_0), .Z(N499) );
  GTECH_AND2 C911 ( .A(N6), .B(m3stg_exp_lt_neg57), .Z(N502) );
  GTECH_AND2 C912 ( .A(N505), .B(m3stg_exp_inv_plus2[5]), .Z(N506) );
  GTECH_AND2 C913 ( .A(N6), .B(N504), .Z(N505) );
  GTECH_NOT I_108 ( .A(m3stg_exp_lt_neg57), .Z(N504) );
  GTECH_AND2 C915 ( .A(m3stg_expadd_lte_0_inv), .B(N508), .Z(N509) );
  GTECH_NOT I_109 ( .A(m3stg_ld0_inv[5]), .Z(N508) );
  GTECH_OR2 C917 ( .A(N516), .B(N518), .Z(m4stg_sh_cnt_in[4]) );
  GTECH_OR2 C918 ( .A(N513), .B(N515), .Z(N516) );
  GTECH_OR2 C919 ( .A(N511), .B(N512), .Z(N513) );
  GTECH_AND2 C920 ( .A(N510), .B(m3stg_exp_minus1[4]), .Z(N511) );
  GTECH_AND2 C921 ( .A(N488), .B(N499), .Z(N510) );
  GTECH_AND2 C923 ( .A(N6), .B(m3stg_exp_lt_neg57), .Z(N512) );
  GTECH_AND2 C924 ( .A(N514), .B(m3stg_exp_inv_plus2[4]), .Z(N515) );
  GTECH_AND2 C925 ( .A(N6), .B(N504), .Z(N514) );
  GTECH_AND2 C927 ( .A(m3stg_expadd_lte_0_inv), .B(N517), .Z(N518) );
  GTECH_NOT I_110 ( .A(m3stg_ld0_inv[4]), .Z(N517) );
  GTECH_OR2 C929 ( .A(N525), .B(N527), .Z(m4stg_sh_cnt_in[3]) );
  GTECH_OR2 C930 ( .A(N522), .B(N524), .Z(N525) );
  GTECH_OR2 C931 ( .A(N520), .B(N521), .Z(N522) );
  GTECH_AND2 C932 ( .A(N519), .B(m3stg_exp_minus1[3]), .Z(N520) );
  GTECH_AND2 C933 ( .A(N488), .B(N499), .Z(N519) );
  GTECH_AND2 C935 ( .A(N6), .B(m3stg_exp_lt_neg57), .Z(N521) );
  GTECH_AND2 C936 ( .A(N523), .B(m3stg_exp_inv_plus2[3]), .Z(N524) );
  GTECH_AND2 C937 ( .A(N6), .B(N504), .Z(N523) );
  GTECH_AND2 C939 ( .A(m3stg_expadd_lte_0_inv), .B(N526), .Z(N527) );
  GTECH_NOT I_111 ( .A(m3stg_ld0_inv[3]), .Z(N526) );
  GTECH_OR2 C941 ( .A(N532), .B(N534), .Z(m4stg_sh_cnt_in[2]) );
  GTECH_OR2 C942 ( .A(N529), .B(N531), .Z(N532) );
  GTECH_AND2 C943 ( .A(N528), .B(m3stg_exp_minus1[2]), .Z(N529) );
  GTECH_AND2 C944 ( .A(N488), .B(N499), .Z(N528) );
  GTECH_AND2 C946 ( .A(N530), .B(m3stg_exp_inv_plus2[2]), .Z(N531) );
  GTECH_AND2 C947 ( .A(N6), .B(N504), .Z(N530) );
  GTECH_AND2 C949 ( .A(m3stg_expadd_lte_0_inv), .B(N533), .Z(N534) );
  GTECH_NOT I_112 ( .A(m3stg_ld0_inv[2]), .Z(N533) );
  GTECH_OR2 C951 ( .A(N539), .B(N541), .Z(m4stg_sh_cnt_in[1]) );
  GTECH_OR2 C952 ( .A(N536), .B(N538), .Z(N539) );
  GTECH_AND2 C953 ( .A(N535), .B(m3stg_exp_minus1[1]), .Z(N536) );
  GTECH_AND2 C954 ( .A(N488), .B(N499), .Z(N535) );
  GTECH_AND2 C956 ( .A(N537), .B(m3stg_exp_inv_plus2[1]), .Z(N538) );
  GTECH_AND2 C957 ( .A(N6), .B(N504), .Z(N537) );
  GTECH_AND2 C959 ( .A(m3stg_expadd_lte_0_inv), .B(N540), .Z(N541) );
  GTECH_NOT I_113 ( .A(m3stg_ld0_inv[1]), .Z(N540) );
  GTECH_OR2 C961 ( .A(N548), .B(N550), .Z(m4stg_sh_cnt_in[0]) );
  GTECH_OR2 C962 ( .A(N545), .B(N547), .Z(N548) );
  GTECH_OR2 C963 ( .A(N543), .B(N544), .Z(N545) );
  GTECH_AND2 C964 ( .A(N542), .B(m3stg_exp_minus1[0]), .Z(N543) );
  GTECH_AND2 C965 ( .A(N488), .B(N499), .Z(N542) );
  GTECH_AND2 C967 ( .A(N6), .B(m3stg_exp_lt_neg57), .Z(N544) );
  GTECH_AND2 C968 ( .A(N546), .B(m3stg_exp_inv_plus2[0]), .Z(N547) );
  GTECH_AND2 C969 ( .A(N6), .B(N504), .Z(N546) );
  GTECH_AND2 C971 ( .A(m3stg_expadd_lte_0_inv), .B(N549), .Z(N550) );
  GTECH_NOT I_114 ( .A(m3stg_ld0_inv[0]), .Z(N549) );
  GTECH_AND2 C973 ( .A(N551), .B(m6stg_step), .Z(m4stg_left_shift_step) );
  GTECH_NOT I_115 ( .A(m4stg_right_shift), .Z(N551) );
  GTECH_AND2 C975 ( .A(m4stg_right_shift), .B(m6stg_step), .Z(
        m4stg_right_shift_step) );
  GTECH_AND2 C976 ( .A(N564), .B(N551), .Z(m4stg_inc_exp_54) );
  GTECH_NOT I_116 ( .A(N563), .Z(N564) );
  GTECH_OR2 C978 ( .A(N562), .B(m4stg_exp[0]), .Z(N563) );
  GTECH_OR2 C979 ( .A(N561), .B(m4stg_exp[1]), .Z(N562) );
  GTECH_OR2 C980 ( .A(N560), .B(m4stg_exp[2]), .Z(N561) );
  GTECH_OR2 C981 ( .A(N559), .B(m4stg_exp[3]), .Z(N560) );
  GTECH_OR2 C982 ( .A(N558), .B(m4stg_exp[4]), .Z(N559) );
  GTECH_OR2 C983 ( .A(N557), .B(m4stg_exp[5]), .Z(N558) );
  GTECH_OR2 C984 ( .A(N556), .B(m4stg_exp[6]), .Z(N557) );
  GTECH_OR2 C985 ( .A(N555), .B(m4stg_exp[7]), .Z(N556) );
  GTECH_OR2 C986 ( .A(N554), .B(m4stg_exp[8]), .Z(N555) );
  GTECH_OR2 C987 ( .A(N553), .B(m4stg_exp[9]), .Z(N554) );
  GTECH_OR2 C988 ( .A(N552), .B(m4stg_exp[10]), .Z(N553) );
  GTECH_OR2 C989 ( .A(m4stg_exp[12]), .B(m4stg_exp[11]), .Z(N552) );
  GTECH_NOT I_117 ( .A(m4stg_right_shift), .Z(m4stg_inc_exp_55) );
  GTECH_AND2 C992 ( .A(N565), .B(m4stg_frac_105), .Z(m4stg_inc_exp_105) );
  GTECH_AND2 C993 ( .A(m4stg_expadd_eq_0), .B(m4stg_right_shift), .Z(N565) );
  GTECH_NOT I_118 ( .A(m5stg_sign), .Z(N7) );
  GTECH_OR2 C995 ( .A(N575), .B(N585), .Z(m5stg_rndup) );
  GTECH_AND2 C996 ( .A(N574), .B(m5stg_fmuld), .Z(N575) );
  GTECH_OR2 C997 ( .A(N570), .B(N573), .Z(N574) );
  GTECH_OR2 C998 ( .A(N567), .B(N569), .Z(N570) );
  GTECH_AND2 C999 ( .A(N566), .B(N113), .Z(N567) );
  GTECH_AND2 C1000 ( .A(N111), .B(N7), .Z(N566) );
  GTECH_AND2 C1001 ( .A(N568), .B(N113), .Z(N569) );
  GTECH_AND2 C1002 ( .A(N114), .B(m5stg_sign), .Z(N568) );
  GTECH_AND2 C1003 ( .A(N571), .B(N572), .Z(N573) );
  GTECH_AND2 C1004 ( .A(N116), .B(m5stg_frac[2]), .Z(N571) );
  GTECH_OR2 C1005 ( .A(N117), .B(m5stg_frac[3]), .Z(N572) );
  GTECH_AND2 C1006 ( .A(N584), .B(m5stg_fmuls), .Z(N585) );
  GTECH_OR2 C1007 ( .A(N580), .B(N583), .Z(N584) );
  GTECH_OR2 C1008 ( .A(N577), .B(N579), .Z(N580) );
  GTECH_AND2 C1009 ( .A(N576), .B(N150), .Z(N577) );
  GTECH_AND2 C1010 ( .A(N119), .B(N7), .Z(N576) );
  GTECH_AND2 C1011 ( .A(N578), .B(N150), .Z(N579) );
  GTECH_AND2 C1012 ( .A(N151), .B(m5stg_sign), .Z(N578) );
  GTECH_AND2 C1013 ( .A(N581), .B(N582), .Z(N583) );
  GTECH_AND2 C1014 ( .A(N153), .B(m5stg_frac[31]), .Z(N581) );
  GTECH_OR2 C1015 ( .A(N183), .B(m5stg_frac[32]), .Z(N582) );
  GTECH_OR2 C1016 ( .A(N587), .B(N589), .Z(m5stg_to_0) );
  GTECH_OR2 C1017 ( .A(N81), .B(N586), .Z(N587) );
  GTECH_AND2 C1018 ( .A(N84), .B(m5stg_sign), .Z(N586) );
  GTECH_AND2 C1019 ( .A(N85), .B(N588), .Z(N589) );
  GTECH_NOT I_119 ( .A(m5stg_sign), .Z(N588) );
  GTECH_NOT I_120 ( .A(m5stg_to_0), .Z(m5stg_to_0_inv) );
  GTECH_AND2 C1022 ( .A(m5stg_rndup), .B(N590), .Z(mul_frac_out_fracadd) );
  GTECH_NOT I_121 ( .A(m5stg_in_of), .Z(N590) );
  GTECH_AND2 C1024 ( .A(N591), .B(N592), .Z(mul_frac_out_frac) );
  GTECH_NOT I_122 ( .A(m5stg_rndup), .Z(N591) );
  GTECH_NOT I_123 ( .A(m5stg_in_of), .Z(N592) );
  GTECH_AND2 C1027 ( .A(m5stg_rndup), .B(N593), .Z(mul_exp_out_exp_plus1) );
  GTECH_NOT I_124 ( .A(m5stg_in_of), .Z(N593) );
  GTECH_AND2 C1029 ( .A(N591), .B(N594), .Z(mul_exp_out_exp) );
  GTECH_NOT I_125 ( .A(m5stg_in_of), .Z(N594) );
endmodule


module fpu_mul_exp_dp ( inq_in1, inq_in2, m6stg_step, m1stg_dblop, m1stg_sngop, 
        m2stg_exp_expadd, m2stg_exp_0bff, m2stg_exp_017f, m2stg_exp_04ff, 
        m2stg_exp_zero, m1stg_fsmuld, m2stg_fmuld, m2stg_fmuls, m2stg_fsmuld, 
        m3stg_ld0_inv, m5stg_fracadd_cout, mul_exp_out_exp_plus1, 
        mul_exp_out_exp, m5stg_in_of, m5stg_fmuld, m5stg_to_0_inv, 
        m4stg_shl_54, m4stg_shl_55, m4stg_inc_exp_54, m4stg_inc_exp_55, 
        m4stg_inc_exp_105, fmul_clken_l, rclk, m3stg_exp, m3stg_expadd_eq_0, 
        m3stg_expadd_lte_0_inv, m4stg_exp, m5stg_exp, mul_exp_out, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [6:0] m3stg_ld0_inv;
  output [12:0] m3stg_exp;
  output [12:0] m4stg_exp;
  output [12:0] m5stg_exp;
  output [10:0] mul_exp_out;
  input m6stg_step, m1stg_dblop, m1stg_sngop, m2stg_exp_expadd, m2stg_exp_0bff,
         m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero, m1stg_fsmuld,
         m2stg_fmuld, m2stg_fmuls, m2stg_fsmuld, m5stg_fracadd_cout,
         mul_exp_out_exp_plus1, mul_exp_out_exp, m5stg_in_of, m5stg_fmuld,
         m5stg_to_0_inv, m4stg_shl_54, m4stg_shl_55, m4stg_inc_exp_54,
         m4stg_inc_exp_55, m4stg_inc_exp_105, fmul_clken_l, rclk, se, si;
  output m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv, so;
  wire   se_l, clk, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13,
         N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, m5stg_shl_55,
         m5stg_shl_54, m5stg_inc_exp_54, m5stg_inc_exp_55, m5stg_inc_exp_105,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         net14294, net14295, net14296, net14297, net14298, net14299, net14300,
         net14301, net14302, net14303, net14304, net14305, net14306, net14307,
         net14308, net14309, net14310, net14311, net14312, net14313, net14314,
         net14315, net14316, net14317, net14318, net14319, net14320, net14321,
         net14322, net14323, net14324, net14325, net14326, net14327, net14328,
         net14329, net14330, net14331, net14332, net14333, net14334, net14335,
         net14336, net14337, net14338, net14339, net14340, net14341, net14342,
         net14343, net14344, net14345, net14346, net14347, net14348, net14349,
         net14350, net14351, net14352, net14353, net14354, net14355, net14356,
         net14357, net14358, net14359, net14360, net14361, net14362, net14363,
         net14364, net14365, net14366, net14367, net14368, net14369, net14370,
         net14371, net14372, net14373, net14374, net14375, net14376, net14377,
         net14378, net14379, net14380, net14381, net14382, net14383, net14384,
         net14385, net14386, net14387, net14388, net14389, net14390, net14391,
         net14392, net14393, net14394, net14395, net14396, net14397, net14398,
         net14399, net14400, net14401, net14402, net14403, net14404, net14405,
         net14406, net14407, net14408, net14409, net14410, net14411, net14412,
         net14413, net14414, net14415, net14416, net14417, net14418, net14419,
         net14420, net14421, net14422, net14423, net14424, net14425, net14426,
         net14427, net14428, net14429, net14430, net14431, net14432, net14433,
         net14434, net14435, net14436, net14437, net14438, net14439, net14440,
         net14441, net14442, net14443, net14444, net14445, net14446, net14447,
         net14448, net14449;
  wire   [10:0] m1stg_exp_in1;
  wire   [10:0] m1stg_exp_in2;
  wire   [10:0] m1stg_expadd_in1;
  wire   [10:0] m1stg_expadd_in2;
  wire   [12:0] m1stg_expadd;
  wire   [12:0] m2stg_exp_in;
  wire   [12:0] m2stg_exp;
  wire   [12:8] m2stg_expadd_in2;
  wire   [12:0] m2stg_expadd;
  wire   [12:0] m3astg_exp;
  wire   [12:0] m3bstg_exp;
  wire   [12:0] m3stg_expa;
  wire   [12:0] m3stg_expadd;
  wire   [12:0] m4stg_exp_in;
  wire   [12:0] m4stg_exp_plus1;
  wire   [12:0] m5stg_exp_pre1_in;
  wire   [12:0] m5stg_exp_pre1;
  wire   [12:0] m5stg_exp_pre2_in;
  wire   [12:0] m5stg_exp_pre2;
  wire   [12:0] m5stg_exp_pre3_in;
  wire   [12:0] m5stg_exp_pre3;
  wire   [10:0] m5stg_exp_plus1;
  wire   [10:0] mul_exp_out_in;

  clken_buf ckbuf_mul_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fmul_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE11 i_m1stg_exp_in1 ( .din(inq_in1), .en(m6stg_step), .clk(clk), .q(
        m1stg_exp_in1), .se(se), .si({net14439, net14440, net14441, net14442, 
        net14443, net14444, net14445, net14446, net14447, net14448, net14449})
         );
  dffe_SIZE11 i_m1stg_exp_in2 ( .din(inq_in2), .en(m6stg_step), .clk(clk), .q(
        m1stg_exp_in2), .se(se), .si({net14428, net14429, net14430, net14431, 
        net14432, net14433, net14434, net14435, net14436, net14437, net14438})
         );
  dffe_SIZE13 i_m2stg_exp ( .din(m2stg_exp_in), .en(m6stg_step), .clk(clk), 
        .q(m2stg_exp), .se(se), .si({net14415, net14416, net14417, net14418, 
        net14419, net14420, net14421, net14422, net14423, net14424, net14425, 
        net14426, net14427}) );
  dffe_SIZE13 i_m3astg_exp ( .din(m2stg_expadd), .en(m6stg_step), .clk(clk), 
        .q(m3astg_exp), .se(se), .si({net14402, net14403, net14404, net14405, 
        net14406, net14407, net14408, net14409, net14410, net14411, net14412, 
        net14413, net14414}) );
  dffe_SIZE13 i_m3bstg_exp ( .din(m3astg_exp), .en(m6stg_step), .clk(clk), .q(
        m3bstg_exp), .se(se), .si({net14389, net14390, net14391, net14392, 
        net14393, net14394, net14395, net14396, net14397, net14398, net14399, 
        net14400, net14401}) );
  dffe_SIZE13 i_m3stg_exp ( .din(m3bstg_exp), .en(m6stg_step), .clk(clk), .q(
        m3stg_exp), .se(se), .si({net14376, net14377, net14378, net14379, 
        net14380, net14381, net14382, net14383, net14384, net14385, net14386, 
        net14387, net14388}) );
  dffe_SIZE13 i_m3stg_expa ( .din(m3bstg_exp), .en(m6stg_step), .clk(clk), .q(
        m3stg_expa), .se(se), .si({net14363, net14364, net14365, net14366, 
        net14367, net14368, net14369, net14370, net14371, net14372, net14373, 
        net14374, net14375}) );
  dffe_SIZE13 i_m4stg_exp ( .din(m4stg_exp_in), .en(m6stg_step), .clk(clk), 
        .q(m4stg_exp), .se(se), .si({net14350, net14351, net14352, net14353, 
        net14354, net14355, net14356, net14357, net14358, net14359, net14360, 
        net14361, net14362}) );
  dff_SIZE13 i_m5stg_exp_pre1 ( .din(m5stg_exp_pre1_in), .clk(clk), .q(
        m5stg_exp_pre1), .se(se), .si({net14337, net14338, net14339, net14340, 
        net14341, net14342, net14343, net14344, net14345, net14346, net14347, 
        net14348, net14349}) );
  dff_SIZE13 i_m5stg_exp_pre2 ( .din(m5stg_exp_pre2_in), .clk(clk), .q(
        m5stg_exp_pre2), .se(se), .si({net14324, net14325, net14326, net14327, 
        net14328, net14329, net14330, net14331, net14332, net14333, net14334, 
        net14335, net14336}) );
  dff_SIZE13 i_m5stg_exp_pre3 ( .din(m5stg_exp_pre3_in), .clk(clk), .q(
        m5stg_exp_pre3), .se(se), .si({net14311, net14312, net14313, net14314, 
        net14315, net14316, net14317, net14318, net14319, net14320, net14321, 
        net14322, net14323}) );
  dff_SIZE5 i_m5stg_inc_exp ( .din({m4stg_shl_55, m4stg_shl_54, 
        m4stg_inc_exp_54, m4stg_inc_exp_55, m4stg_inc_exp_105}), .clk(clk), 
        .q({m5stg_shl_55, m5stg_shl_54, m5stg_inc_exp_54, m5stg_inc_exp_55, 
        m5stg_inc_exp_105}), .se(se), .si({net14306, net14307, net14308, 
        net14309, net14310}) );
  dffe_SIZE11 i_mul_exp_out ( .din(mul_exp_out_in), .en(m6stg_step), .clk(clk), 
        .q(mul_exp_out), .se(se), .si({net14295, net14296, net14297, net14298, 
        net14299, net14300, net14301, net14302, net14303, net14304, net14305})
         );
  ADD_UNS_OP add_247 ( .A(m2stg_exp), .B({m2stg_expadd_in2, m2stg_fmuls, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Z(m2stg_expadd) );
  ADD_UNS_OP add_204 ( .A(m1stg_expadd_in1), .B(m1stg_expadd_in2), .Z({N11, 
        N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  ADD_UNS_OP add_325 ( .A(m3stg_expa), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        m3stg_ld0_inv}), .Z({N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12}) );
  ADD_UNS_OP add_356 ( .A(m4stg_exp), .B(1'b1), .Z(m4stg_exp_plus1) );
  ADD_UNS_OP add_204_2 ( .A({N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), .B(1'b1), .Z(m1stg_expadd) );
  ADD_UNS_OP add_325_2 ( .A({N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12}), .B(1'b1), .Z(m3stg_expadd) );
  ADD_UNS_OP add_462 ( .A(m5stg_exp[10:0]), .B(1'b1), .Z(m5stg_exp_plus1) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_AND2 C128 ( .A(m1stg_dblop), .B(m1stg_exp_in1[10]), .Z(
        m1stg_expadd_in1[10]) );
  GTECH_AND2 C129 ( .A(m1stg_dblop), .B(m1stg_exp_in1[9]), .Z(
        m1stg_expadd_in1[9]) );
  GTECH_AND2 C130 ( .A(m1stg_dblop), .B(m1stg_exp_in1[8]), .Z(
        m1stg_expadd_in1[8]) );
  GTECH_OR2 C131 ( .A(N26), .B(N27), .Z(m1stg_expadd_in1[7]) );
  GTECH_AND2 C132 ( .A(m1stg_dblop), .B(m1stg_exp_in1[7]), .Z(N26) );
  GTECH_AND2 C133 ( .A(m1stg_sngop), .B(m1stg_exp_in1[10]), .Z(N27) );
  GTECH_OR2 C134 ( .A(N28), .B(N29), .Z(m1stg_expadd_in1[6]) );
  GTECH_AND2 C135 ( .A(m1stg_dblop), .B(m1stg_exp_in1[6]), .Z(N28) );
  GTECH_AND2 C136 ( .A(m1stg_sngop), .B(m1stg_exp_in1[9]), .Z(N29) );
  GTECH_OR2 C137 ( .A(N30), .B(N31), .Z(m1stg_expadd_in1[5]) );
  GTECH_AND2 C138 ( .A(m1stg_dblop), .B(m1stg_exp_in1[5]), .Z(N30) );
  GTECH_AND2 C139 ( .A(m1stg_sngop), .B(m1stg_exp_in1[8]), .Z(N31) );
  GTECH_OR2 C140 ( .A(N32), .B(N33), .Z(m1stg_expadd_in1[4]) );
  GTECH_AND2 C141 ( .A(m1stg_dblop), .B(m1stg_exp_in1[4]), .Z(N32) );
  GTECH_AND2 C142 ( .A(m1stg_sngop), .B(m1stg_exp_in1[7]), .Z(N33) );
  GTECH_OR2 C143 ( .A(N34), .B(N35), .Z(m1stg_expadd_in1[3]) );
  GTECH_AND2 C144 ( .A(m1stg_dblop), .B(m1stg_exp_in1[3]), .Z(N34) );
  GTECH_AND2 C145 ( .A(m1stg_sngop), .B(m1stg_exp_in1[6]), .Z(N35) );
  GTECH_OR2 C146 ( .A(N36), .B(N37), .Z(m1stg_expadd_in1[2]) );
  GTECH_AND2 C147 ( .A(m1stg_dblop), .B(m1stg_exp_in1[2]), .Z(N36) );
  GTECH_AND2 C148 ( .A(m1stg_sngop), .B(m1stg_exp_in1[5]), .Z(N37) );
  GTECH_OR2 C149 ( .A(N38), .B(N39), .Z(m1stg_expadd_in1[1]) );
  GTECH_AND2 C150 ( .A(m1stg_dblop), .B(m1stg_exp_in1[1]), .Z(N38) );
  GTECH_AND2 C151 ( .A(m1stg_sngop), .B(m1stg_exp_in1[4]), .Z(N39) );
  GTECH_OR2 C152 ( .A(N40), .B(N41), .Z(m1stg_expadd_in1[0]) );
  GTECH_AND2 C153 ( .A(m1stg_dblop), .B(m1stg_exp_in1[0]), .Z(N40) );
  GTECH_AND2 C154 ( .A(m1stg_sngop), .B(m1stg_exp_in1[3]), .Z(N41) );
  GTECH_AND2 C155 ( .A(m1stg_dblop), .B(m1stg_exp_in2[10]), .Z(
        m1stg_expadd_in2[10]) );
  GTECH_AND2 C156 ( .A(m1stg_dblop), .B(m1stg_exp_in2[9]), .Z(
        m1stg_expadd_in2[9]) );
  GTECH_AND2 C157 ( .A(m1stg_dblop), .B(m1stg_exp_in2[8]), .Z(
        m1stg_expadd_in2[8]) );
  GTECH_OR2 C158 ( .A(N42), .B(N43), .Z(m1stg_expadd_in2[7]) );
  GTECH_AND2 C159 ( .A(m1stg_dblop), .B(m1stg_exp_in2[7]), .Z(N42) );
  GTECH_AND2 C160 ( .A(m1stg_sngop), .B(m1stg_exp_in2[10]), .Z(N43) );
  GTECH_OR2 C161 ( .A(N44), .B(N45), .Z(m1stg_expadd_in2[6]) );
  GTECH_AND2 C162 ( .A(m1stg_dblop), .B(m1stg_exp_in2[6]), .Z(N44) );
  GTECH_AND2 C163 ( .A(m1stg_sngop), .B(m1stg_exp_in2[9]), .Z(N45) );
  GTECH_OR2 C164 ( .A(N46), .B(N47), .Z(m1stg_expadd_in2[5]) );
  GTECH_AND2 C165 ( .A(m1stg_dblop), .B(m1stg_exp_in2[5]), .Z(N46) );
  GTECH_AND2 C166 ( .A(m1stg_sngop), .B(m1stg_exp_in2[8]), .Z(N47) );
  GTECH_OR2 C167 ( .A(N48), .B(N49), .Z(m1stg_expadd_in2[4]) );
  GTECH_AND2 C168 ( .A(m1stg_dblop), .B(m1stg_exp_in2[4]), .Z(N48) );
  GTECH_AND2 C169 ( .A(m1stg_sngop), .B(m1stg_exp_in2[7]), .Z(N49) );
  GTECH_OR2 C170 ( .A(N50), .B(N51), .Z(m1stg_expadd_in2[3]) );
  GTECH_AND2 C171 ( .A(m1stg_dblop), .B(m1stg_exp_in2[3]), .Z(N50) );
  GTECH_AND2 C172 ( .A(m1stg_sngop), .B(m1stg_exp_in2[6]), .Z(N51) );
  GTECH_OR2 C173 ( .A(N52), .B(N53), .Z(m1stg_expadd_in2[2]) );
  GTECH_AND2 C174 ( .A(m1stg_dblop), .B(m1stg_exp_in2[2]), .Z(N52) );
  GTECH_AND2 C175 ( .A(m1stg_sngop), .B(m1stg_exp_in2[5]), .Z(N53) );
  GTECH_OR2 C176 ( .A(N54), .B(N55), .Z(m1stg_expadd_in2[1]) );
  GTECH_AND2 C177 ( .A(m1stg_dblop), .B(m1stg_exp_in2[1]), .Z(N54) );
  GTECH_AND2 C178 ( .A(m1stg_sngop), .B(m1stg_exp_in2[4]), .Z(N55) );
  GTECH_OR2 C179 ( .A(N56), .B(N57), .Z(m1stg_expadd_in2[0]) );
  GTECH_AND2 C180 ( .A(m1stg_dblop), .B(m1stg_exp_in2[0]), .Z(N56) );
  GTECH_AND2 C181 ( .A(m1stg_sngop), .B(m1stg_exp_in2[3]), .Z(N57) );
  GTECH_OR2 C182 ( .A(N58), .B(N59), .Z(m2stg_exp_in[12]) );
  GTECH_AND2 C183 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[12]), .Z(N58) );
  GTECH_AND2 C184 ( .A(m2stg_exp_zero), .B(m1stg_fsmuld), .Z(N59) );
  GTECH_OR2 C185 ( .A(N61), .B(N62), .Z(m2stg_exp_in[11]) );
  GTECH_OR2 C186 ( .A(N60), .B(m2stg_exp_0bff), .Z(N61) );
  GTECH_AND2 C187 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[11]), .Z(N60) );
  GTECH_AND2 C188 ( .A(m2stg_exp_zero), .B(m1stg_fsmuld), .Z(N62) );
  GTECH_OR2 C189 ( .A(N64), .B(N65), .Z(m2stg_exp_in[10]) );
  GTECH_OR2 C190 ( .A(N63), .B(m2stg_exp_04ff), .Z(N64) );
  GTECH_AND2 C191 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[10]), .Z(N63) );
  GTECH_AND2 C192 ( .A(m2stg_exp_zero), .B(m1stg_fsmuld), .Z(N65) );
  GTECH_OR2 C193 ( .A(N66), .B(m2stg_exp_0bff), .Z(m2stg_exp_in[9]) );
  GTECH_AND2 C194 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[9]), .Z(N66) );
  GTECH_OR2 C195 ( .A(N68), .B(m2stg_exp_017f), .Z(m2stg_exp_in[8]) );
  GTECH_OR2 C196 ( .A(N67), .B(m2stg_exp_0bff), .Z(N68) );
  GTECH_AND2 C197 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[8]), .Z(N67) );
  GTECH_OR2 C198 ( .A(N70), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[7]) );
  GTECH_OR2 C199 ( .A(N69), .B(m2stg_exp_0bff), .Z(N70) );
  GTECH_AND2 C200 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[7]), .Z(N69) );
  GTECH_OR2 C201 ( .A(N73), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[6]) );
  GTECH_OR2 C202 ( .A(N72), .B(m2stg_exp_017f), .Z(N73) );
  GTECH_OR2 C203 ( .A(N71), .B(m2stg_exp_0bff), .Z(N72) );
  GTECH_AND2 C204 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[6]), .Z(N71) );
  GTECH_OR2 C205 ( .A(N76), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[5]) );
  GTECH_OR2 C206 ( .A(N75), .B(m2stg_exp_017f), .Z(N76) );
  GTECH_OR2 C207 ( .A(N74), .B(m2stg_exp_0bff), .Z(N75) );
  GTECH_AND2 C208 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[5]), .Z(N74) );
  GTECH_OR2 C209 ( .A(N79), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[4]) );
  GTECH_OR2 C210 ( .A(N78), .B(m2stg_exp_017f), .Z(N79) );
  GTECH_OR2 C211 ( .A(N77), .B(m2stg_exp_0bff), .Z(N78) );
  GTECH_AND2 C212 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[4]), .Z(N77) );
  GTECH_OR2 C213 ( .A(N82), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[3]) );
  GTECH_OR2 C214 ( .A(N81), .B(m2stg_exp_017f), .Z(N82) );
  GTECH_OR2 C215 ( .A(N80), .B(m2stg_exp_0bff), .Z(N81) );
  GTECH_AND2 C216 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[3]), .Z(N80) );
  GTECH_OR2 C217 ( .A(N85), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[2]) );
  GTECH_OR2 C218 ( .A(N84), .B(m2stg_exp_017f), .Z(N85) );
  GTECH_OR2 C219 ( .A(N83), .B(m2stg_exp_0bff), .Z(N84) );
  GTECH_AND2 C220 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[2]), .Z(N83) );
  GTECH_OR2 C221 ( .A(N88), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[1]) );
  GTECH_OR2 C222 ( .A(N87), .B(m2stg_exp_017f), .Z(N88) );
  GTECH_OR2 C223 ( .A(N86), .B(m2stg_exp_0bff), .Z(N87) );
  GTECH_AND2 C224 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[1]), .Z(N86) );
  GTECH_OR2 C225 ( .A(N91), .B(m2stg_exp_04ff), .Z(m2stg_exp_in[0]) );
  GTECH_OR2 C226 ( .A(N90), .B(m2stg_exp_017f), .Z(N91) );
  GTECH_OR2 C227 ( .A(N89), .B(m2stg_exp_0bff), .Z(N90) );
  GTECH_AND2 C228 ( .A(m2stg_exp_expadd), .B(m1stg_expadd[0]), .Z(N89) );
  GTECH_OR2 C229 ( .A(m2stg_fmuld), .B(m2stg_fmuls), .Z(m2stg_expadd_in2[12])
         );
  GTECH_OR2 C230 ( .A(m2stg_fmuld), .B(m2stg_fmuls), .Z(m2stg_expadd_in2[11])
         );
  GTECH_OR2 C231 ( .A(m2stg_fmuld), .B(m2stg_fmuls), .Z(m2stg_expadd_in2[10])
         );
  GTECH_OR2 C232 ( .A(m2stg_fmuls), .B(m2stg_fsmuld), .Z(m2stg_expadd_in2[9])
         );
  GTECH_OR2 C233 ( .A(m2stg_fmuls), .B(m2stg_fsmuld), .Z(m2stg_expadd_in2[8])
         );
  GTECH_AND2 C234 ( .A(N114), .B(N115), .Z(m3stg_expadd_eq_0) );
  GTECH_AND2 C235 ( .A(N112), .B(N113), .Z(N114) );
  GTECH_AND2 C236 ( .A(N110), .B(N111), .Z(N112) );
  GTECH_AND2 C237 ( .A(N108), .B(N109), .Z(N110) );
  GTECH_AND2 C238 ( .A(N106), .B(N107), .Z(N108) );
  GTECH_AND2 C239 ( .A(N104), .B(N105), .Z(N106) );
  GTECH_AND2 C240 ( .A(N102), .B(N103), .Z(N104) );
  GTECH_AND2 C241 ( .A(N100), .B(N101), .Z(N102) );
  GTECH_AND2 C242 ( .A(N98), .B(N99), .Z(N100) );
  GTECH_AND2 C243 ( .A(N96), .B(N97), .Z(N98) );
  GTECH_AND2 C244 ( .A(N94), .B(N95), .Z(N96) );
  GTECH_AND2 C245 ( .A(N92), .B(N93), .Z(N94) );
  GTECH_NOT I_1 ( .A(m3stg_exp[12]), .Z(N92) );
  GTECH_NOT I_2 ( .A(m3stg_exp[11]), .Z(N93) );
  GTECH_NOT I_3 ( .A(m3stg_exp[10]), .Z(N95) );
  GTECH_NOT I_4 ( .A(m3stg_exp[9]), .Z(N97) );
  GTECH_NOT I_5 ( .A(m3stg_exp[8]), .Z(N99) );
  GTECH_NOT I_6 ( .A(m3stg_exp[7]), .Z(N101) );
  GTECH_XOR2 C252 ( .A(m3stg_exp[6]), .B(m3stg_ld0_inv[6]), .Z(N103) );
  GTECH_XOR2 C253 ( .A(m3stg_exp[5]), .B(m3stg_ld0_inv[5]), .Z(N105) );
  GTECH_XOR2 C254 ( .A(m3stg_exp[4]), .B(m3stg_ld0_inv[4]), .Z(N107) );
  GTECH_XOR2 C255 ( .A(m3stg_exp[3]), .B(m3stg_ld0_inv[3]), .Z(N109) );
  GTECH_XOR2 C256 ( .A(m3stg_exp[2]), .B(m3stg_ld0_inv[2]), .Z(N111) );
  GTECH_XOR2 C257 ( .A(m3stg_exp[1]), .B(m3stg_ld0_inv[1]), .Z(N113) );
  GTECH_XOR2 C258 ( .A(m3stg_exp[0]), .B(m3stg_ld0_inv[0]), .Z(N115) );
  GTECH_NOT I_7 ( .A(N116), .Z(m3stg_expadd_lte_0_inv) );
  GTECH_OR2 C260 ( .A(m3stg_expadd[12]), .B(m3stg_expadd_eq_0), .Z(N116) );
  GTECH_AND2 C261 ( .A(m3stg_expadd[12]), .B(N117), .Z(m4stg_exp_in[12]) );
  GTECH_NOT I_8 ( .A(m3stg_expadd[12]), .Z(N117) );
  GTECH_AND2 C263 ( .A(m3stg_expadd[11]), .B(N117), .Z(m4stg_exp_in[11]) );
  GTECH_AND2 C265 ( .A(m3stg_expadd[10]), .B(N117), .Z(m4stg_exp_in[10]) );
  GTECH_AND2 C267 ( .A(m3stg_expadd[9]), .B(N117), .Z(m4stg_exp_in[9]) );
  GTECH_AND2 C269 ( .A(m3stg_expadd[8]), .B(N117), .Z(m4stg_exp_in[8]) );
  GTECH_AND2 C271 ( .A(m3stg_expadd[7]), .B(N117), .Z(m4stg_exp_in[7]) );
  GTECH_AND2 C273 ( .A(m3stg_expadd[6]), .B(N117), .Z(m4stg_exp_in[6]) );
  GTECH_AND2 C275 ( .A(m3stg_expadd[5]), .B(N117), .Z(m4stg_exp_in[5]) );
  GTECH_AND2 C277 ( .A(m3stg_expadd[4]), .B(N117), .Z(m4stg_exp_in[4]) );
  GTECH_AND2 C279 ( .A(m3stg_expadd[3]), .B(N117), .Z(m4stg_exp_in[3]) );
  GTECH_AND2 C281 ( .A(m3stg_expadd[2]), .B(N117), .Z(m4stg_exp_in[2]) );
  GTECH_AND2 C283 ( .A(m3stg_expadd[1]), .B(N117), .Z(m4stg_exp_in[1]) );
  GTECH_AND2 C285 ( .A(m3stg_expadd[0]), .B(N117), .Z(m4stg_exp_in[0]) );
  GTECH_AND2 C287 ( .A(m6stg_step), .B(m4stg_exp_plus1[12]), .Z(
        m5stg_exp_pre1_in[12]) );
  GTECH_AND2 C288 ( .A(m6stg_step), .B(m4stg_exp_plus1[11]), .Z(
        m5stg_exp_pre1_in[11]) );
  GTECH_AND2 C289 ( .A(m6stg_step), .B(m4stg_exp_plus1[10]), .Z(
        m5stg_exp_pre1_in[10]) );
  GTECH_AND2 C290 ( .A(m6stg_step), .B(m4stg_exp_plus1[9]), .Z(
        m5stg_exp_pre1_in[9]) );
  GTECH_AND2 C291 ( .A(m6stg_step), .B(m4stg_exp_plus1[8]), .Z(
        m5stg_exp_pre1_in[8]) );
  GTECH_AND2 C292 ( .A(m6stg_step), .B(m4stg_exp_plus1[7]), .Z(
        m5stg_exp_pre1_in[7]) );
  GTECH_AND2 C293 ( .A(m6stg_step), .B(m4stg_exp_plus1[6]), .Z(
        m5stg_exp_pre1_in[6]) );
  GTECH_AND2 C294 ( .A(m6stg_step), .B(m4stg_exp_plus1[5]), .Z(
        m5stg_exp_pre1_in[5]) );
  GTECH_AND2 C295 ( .A(m6stg_step), .B(m4stg_exp_plus1[4]), .Z(
        m5stg_exp_pre1_in[4]) );
  GTECH_AND2 C296 ( .A(m6stg_step), .B(m4stg_exp_plus1[3]), .Z(
        m5stg_exp_pre1_in[3]) );
  GTECH_AND2 C297 ( .A(m6stg_step), .B(m4stg_exp_plus1[2]), .Z(
        m5stg_exp_pre1_in[2]) );
  GTECH_AND2 C298 ( .A(m6stg_step), .B(m4stg_exp_plus1[1]), .Z(
        m5stg_exp_pre1_in[1]) );
  GTECH_AND2 C299 ( .A(m6stg_step), .B(m4stg_exp_plus1[0]), .Z(
        m5stg_exp_pre1_in[0]) );
  GTECH_AND2 C300 ( .A(m6stg_step), .B(m4stg_exp[12]), .Z(
        m5stg_exp_pre2_in[12]) );
  GTECH_AND2 C301 ( .A(m6stg_step), .B(m4stg_exp[11]), .Z(
        m5stg_exp_pre2_in[11]) );
  GTECH_AND2 C302 ( .A(m6stg_step), .B(m4stg_exp[10]), .Z(
        m5stg_exp_pre2_in[10]) );
  GTECH_AND2 C303 ( .A(m6stg_step), .B(m4stg_exp[9]), .Z(m5stg_exp_pre2_in[9])
         );
  GTECH_AND2 C304 ( .A(m6stg_step), .B(m4stg_exp[8]), .Z(m5stg_exp_pre2_in[8])
         );
  GTECH_AND2 C305 ( .A(m6stg_step), .B(m4stg_exp[7]), .Z(m5stg_exp_pre2_in[7])
         );
  GTECH_AND2 C306 ( .A(m6stg_step), .B(m4stg_exp[6]), .Z(m5stg_exp_pre2_in[6])
         );
  GTECH_AND2 C307 ( .A(m6stg_step), .B(m4stg_exp[5]), .Z(m5stg_exp_pre2_in[5])
         );
  GTECH_AND2 C308 ( .A(m6stg_step), .B(m4stg_exp[4]), .Z(m5stg_exp_pre2_in[4])
         );
  GTECH_AND2 C309 ( .A(m6stg_step), .B(m4stg_exp[3]), .Z(m5stg_exp_pre2_in[3])
         );
  GTECH_AND2 C310 ( .A(m6stg_step), .B(m4stg_exp[2]), .Z(m5stg_exp_pre2_in[2])
         );
  GTECH_AND2 C311 ( .A(m6stg_step), .B(m4stg_exp[1]), .Z(m5stg_exp_pre2_in[1])
         );
  GTECH_AND2 C312 ( .A(m6stg_step), .B(m4stg_exp[0]), .Z(m5stg_exp_pre2_in[0])
         );
  GTECH_NOT I_9 ( .A(N119), .Z(m5stg_exp_pre3_in[12]) );
  GTECH_AND2 C314 ( .A(N118), .B(m5stg_exp[12]), .Z(N119) );
  GTECH_NOT I_10 ( .A(m6stg_step), .Z(N118) );
  GTECH_NOT I_11 ( .A(N121), .Z(m5stg_exp_pre3_in[11]) );
  GTECH_AND2 C317 ( .A(N120), .B(m5stg_exp[11]), .Z(N121) );
  GTECH_NOT I_12 ( .A(m6stg_step), .Z(N120) );
  GTECH_NOT I_13 ( .A(N123), .Z(m5stg_exp_pre3_in[10]) );
  GTECH_AND2 C320 ( .A(N122), .B(m5stg_exp[10]), .Z(N123) );
  GTECH_NOT I_14 ( .A(m6stg_step), .Z(N122) );
  GTECH_NOT I_15 ( .A(N125), .Z(m5stg_exp_pre3_in[9]) );
  GTECH_AND2 C323 ( .A(N124), .B(m5stg_exp[9]), .Z(N125) );
  GTECH_NOT I_16 ( .A(m6stg_step), .Z(N124) );
  GTECH_NOT I_17 ( .A(N127), .Z(m5stg_exp_pre3_in[8]) );
  GTECH_AND2 C326 ( .A(N126), .B(m5stg_exp[8]), .Z(N127) );
  GTECH_NOT I_18 ( .A(m6stg_step), .Z(N126) );
  GTECH_NOT I_19 ( .A(N129), .Z(m5stg_exp_pre3_in[7]) );
  GTECH_AND2 C329 ( .A(N128), .B(m5stg_exp[7]), .Z(N129) );
  GTECH_NOT I_20 ( .A(m6stg_step), .Z(N128) );
  GTECH_NOT I_21 ( .A(N131), .Z(m5stg_exp_pre3_in[6]) );
  GTECH_AND2 C332 ( .A(N130), .B(m5stg_exp[6]), .Z(N131) );
  GTECH_NOT I_22 ( .A(m6stg_step), .Z(N130) );
  GTECH_NOT I_23 ( .A(N133), .Z(m5stg_exp_pre3_in[5]) );
  GTECH_AND2 C335 ( .A(N132), .B(m5stg_exp[5]), .Z(N133) );
  GTECH_NOT I_24 ( .A(m6stg_step), .Z(N132) );
  GTECH_NOT I_25 ( .A(N135), .Z(m5stg_exp_pre3_in[4]) );
  GTECH_AND2 C338 ( .A(N134), .B(m5stg_exp[4]), .Z(N135) );
  GTECH_NOT I_26 ( .A(m6stg_step), .Z(N134) );
  GTECH_NOT I_27 ( .A(N137), .Z(m5stg_exp_pre3_in[3]) );
  GTECH_AND2 C341 ( .A(N136), .B(m5stg_exp[3]), .Z(N137) );
  GTECH_NOT I_28 ( .A(m6stg_step), .Z(N136) );
  GTECH_NOT I_29 ( .A(N139), .Z(m5stg_exp_pre3_in[2]) );
  GTECH_AND2 C344 ( .A(N138), .B(m5stg_exp[2]), .Z(N139) );
  GTECH_NOT I_30 ( .A(m6stg_step), .Z(N138) );
  GTECH_NOT I_31 ( .A(N141), .Z(m5stg_exp_pre3_in[1]) );
  GTECH_AND2 C347 ( .A(N140), .B(m5stg_exp[1]), .Z(N141) );
  GTECH_NOT I_32 ( .A(m6stg_step), .Z(N140) );
  GTECH_NOT I_33 ( .A(N143), .Z(m5stg_exp_pre3_in[0]) );
  GTECH_AND2 C350 ( .A(N142), .B(m5stg_exp[0]), .Z(N143) );
  GTECH_NOT I_34 ( .A(m6stg_step), .Z(N142) );
  GTECH_OR2 C352 ( .A(N146), .B(m5stg_inc_exp_105), .Z(N25) );
  GTECH_OR2 C353 ( .A(N144), .B(N145), .Z(N146) );
  GTECH_AND2 C354 ( .A(m5stg_shl_54), .B(m5stg_inc_exp_54), .Z(N144) );
  GTECH_AND2 C355 ( .A(m5stg_shl_55), .B(m5stg_inc_exp_55), .Z(N145) );
  GTECH_OR2 C356 ( .A(N150), .B(N151), .Z(m5stg_exp[12]) );
  GTECH_OR2 C357 ( .A(N147), .B(N149), .Z(N150) );
  GTECH_AND2 C358 ( .A(N25), .B(m5stg_exp_pre1[12]), .Z(N147) );
  GTECH_AND2 C359 ( .A(N148), .B(m5stg_exp_pre2[12]), .Z(N149) );
  GTECH_NOT I_35 ( .A(N25), .Z(N148) );
  GTECH_NOT I_36 ( .A(m5stg_exp_pre3[12]), .Z(N151) );
  GTECH_OR2 C362 ( .A(N154), .B(N155), .Z(m5stg_exp[11]) );
  GTECH_OR2 C363 ( .A(N152), .B(N153), .Z(N154) );
  GTECH_AND2 C364 ( .A(N25), .B(m5stg_exp_pre1[11]), .Z(N152) );
  GTECH_AND2 C365 ( .A(N148), .B(m5stg_exp_pre2[11]), .Z(N153) );
  GTECH_NOT I_37 ( .A(m5stg_exp_pre3[11]), .Z(N155) );
  GTECH_OR2 C368 ( .A(N158), .B(N159), .Z(m5stg_exp[10]) );
  GTECH_OR2 C369 ( .A(N156), .B(N157), .Z(N158) );
  GTECH_AND2 C370 ( .A(N25), .B(m5stg_exp_pre1[10]), .Z(N156) );
  GTECH_AND2 C371 ( .A(N148), .B(m5stg_exp_pre2[10]), .Z(N157) );
  GTECH_NOT I_38 ( .A(m5stg_exp_pre3[10]), .Z(N159) );
  GTECH_OR2 C374 ( .A(N162), .B(N163), .Z(m5stg_exp[9]) );
  GTECH_OR2 C375 ( .A(N160), .B(N161), .Z(N162) );
  GTECH_AND2 C376 ( .A(N25), .B(m5stg_exp_pre1[9]), .Z(N160) );
  GTECH_AND2 C377 ( .A(N148), .B(m5stg_exp_pre2[9]), .Z(N161) );
  GTECH_NOT I_39 ( .A(m5stg_exp_pre3[9]), .Z(N163) );
  GTECH_OR2 C380 ( .A(N166), .B(N167), .Z(m5stg_exp[8]) );
  GTECH_OR2 C381 ( .A(N164), .B(N165), .Z(N166) );
  GTECH_AND2 C382 ( .A(N25), .B(m5stg_exp_pre1[8]), .Z(N164) );
  GTECH_AND2 C383 ( .A(N148), .B(m5stg_exp_pre2[8]), .Z(N165) );
  GTECH_NOT I_40 ( .A(m5stg_exp_pre3[8]), .Z(N167) );
  GTECH_OR2 C386 ( .A(N170), .B(N171), .Z(m5stg_exp[7]) );
  GTECH_OR2 C387 ( .A(N168), .B(N169), .Z(N170) );
  GTECH_AND2 C388 ( .A(N25), .B(m5stg_exp_pre1[7]), .Z(N168) );
  GTECH_AND2 C389 ( .A(N148), .B(m5stg_exp_pre2[7]), .Z(N169) );
  GTECH_NOT I_41 ( .A(m5stg_exp_pre3[7]), .Z(N171) );
  GTECH_OR2 C392 ( .A(N174), .B(N175), .Z(m5stg_exp[6]) );
  GTECH_OR2 C393 ( .A(N172), .B(N173), .Z(N174) );
  GTECH_AND2 C394 ( .A(N25), .B(m5stg_exp_pre1[6]), .Z(N172) );
  GTECH_AND2 C395 ( .A(N148), .B(m5stg_exp_pre2[6]), .Z(N173) );
  GTECH_NOT I_42 ( .A(m5stg_exp_pre3[6]), .Z(N175) );
  GTECH_OR2 C398 ( .A(N178), .B(N179), .Z(m5stg_exp[5]) );
  GTECH_OR2 C399 ( .A(N176), .B(N177), .Z(N178) );
  GTECH_AND2 C400 ( .A(N25), .B(m5stg_exp_pre1[5]), .Z(N176) );
  GTECH_AND2 C401 ( .A(N148), .B(m5stg_exp_pre2[5]), .Z(N177) );
  GTECH_NOT I_43 ( .A(m5stg_exp_pre3[5]), .Z(N179) );
  GTECH_OR2 C404 ( .A(N182), .B(N183), .Z(m5stg_exp[4]) );
  GTECH_OR2 C405 ( .A(N180), .B(N181), .Z(N182) );
  GTECH_AND2 C406 ( .A(N25), .B(m5stg_exp_pre1[4]), .Z(N180) );
  GTECH_AND2 C407 ( .A(N148), .B(m5stg_exp_pre2[4]), .Z(N181) );
  GTECH_NOT I_44 ( .A(m5stg_exp_pre3[4]), .Z(N183) );
  GTECH_OR2 C410 ( .A(N186), .B(N187), .Z(m5stg_exp[3]) );
  GTECH_OR2 C411 ( .A(N184), .B(N185), .Z(N186) );
  GTECH_AND2 C412 ( .A(N25), .B(m5stg_exp_pre1[3]), .Z(N184) );
  GTECH_AND2 C413 ( .A(N148), .B(m5stg_exp_pre2[3]), .Z(N185) );
  GTECH_NOT I_45 ( .A(m5stg_exp_pre3[3]), .Z(N187) );
  GTECH_OR2 C416 ( .A(N190), .B(N191), .Z(m5stg_exp[2]) );
  GTECH_OR2 C417 ( .A(N188), .B(N189), .Z(N190) );
  GTECH_AND2 C418 ( .A(N25), .B(m5stg_exp_pre1[2]), .Z(N188) );
  GTECH_AND2 C419 ( .A(N148), .B(m5stg_exp_pre2[2]), .Z(N189) );
  GTECH_NOT I_46 ( .A(m5stg_exp_pre3[2]), .Z(N191) );
  GTECH_OR2 C422 ( .A(N194), .B(N195), .Z(m5stg_exp[1]) );
  GTECH_OR2 C423 ( .A(N192), .B(N193), .Z(N194) );
  GTECH_AND2 C424 ( .A(N25), .B(m5stg_exp_pre1[1]), .Z(N192) );
  GTECH_AND2 C425 ( .A(N148), .B(m5stg_exp_pre2[1]), .Z(N193) );
  GTECH_NOT I_47 ( .A(m5stg_exp_pre3[1]), .Z(N195) );
  GTECH_OR2 C428 ( .A(N198), .B(N199), .Z(m5stg_exp[0]) );
  GTECH_OR2 C429 ( .A(N196), .B(N197), .Z(N198) );
  GTECH_AND2 C430 ( .A(N25), .B(m5stg_exp_pre1[0]), .Z(N196) );
  GTECH_AND2 C431 ( .A(N148), .B(m5stg_exp_pre2[0]), .Z(N197) );
  GTECH_NOT I_48 ( .A(m5stg_exp_pre3[0]), .Z(N199) );
  GTECH_OR2 C434 ( .A(N208), .B(N209), .Z(mul_exp_out_in[10]) );
  GTECH_OR2 C435 ( .A(N203), .B(N207), .Z(N208) );
  GTECH_OR2 C436 ( .A(N201), .B(N202), .Z(N203) );
  GTECH_AND2 C437 ( .A(N200), .B(m5stg_exp_plus1[10]), .Z(N201) );
  GTECH_AND2 C438 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N200) );
  GTECH_AND2 C439 ( .A(mul_exp_out_exp), .B(m5stg_exp[10]), .Z(N202) );
  GTECH_AND2 C440 ( .A(N206), .B(m5stg_exp[10]), .Z(N207) );
  GTECH_AND2 C441 ( .A(N204), .B(N205), .Z(N206) );
  GTECH_NOT I_49 ( .A(m5stg_fracadd_cout), .Z(N204) );
  GTECH_NOT I_50 ( .A(m5stg_in_of), .Z(N205) );
  GTECH_AND2 C444 ( .A(m5stg_in_of), .B(m5stg_fmuld), .Z(N209) );
  GTECH_OR2 C445 ( .A(N216), .B(N217), .Z(mul_exp_out_in[9]) );
  GTECH_OR2 C446 ( .A(N213), .B(N215), .Z(N216) );
  GTECH_OR2 C447 ( .A(N211), .B(N212), .Z(N213) );
  GTECH_AND2 C448 ( .A(N210), .B(m5stg_exp_plus1[9]), .Z(N211) );
  GTECH_AND2 C449 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N210) );
  GTECH_AND2 C450 ( .A(mul_exp_out_exp), .B(m5stg_exp[9]), .Z(N212) );
  GTECH_AND2 C451 ( .A(N214), .B(m5stg_exp[9]), .Z(N215) );
  GTECH_AND2 C452 ( .A(N204), .B(N205), .Z(N214) );
  GTECH_AND2 C455 ( .A(m5stg_in_of), .B(m5stg_fmuld), .Z(N217) );
  GTECH_OR2 C456 ( .A(N224), .B(N225), .Z(mul_exp_out_in[8]) );
  GTECH_OR2 C457 ( .A(N221), .B(N223), .Z(N224) );
  GTECH_OR2 C458 ( .A(N219), .B(N220), .Z(N221) );
  GTECH_AND2 C459 ( .A(N218), .B(m5stg_exp_plus1[8]), .Z(N219) );
  GTECH_AND2 C460 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N218) );
  GTECH_AND2 C461 ( .A(mul_exp_out_exp), .B(m5stg_exp[8]), .Z(N220) );
  GTECH_AND2 C462 ( .A(N222), .B(m5stg_exp[8]), .Z(N223) );
  GTECH_AND2 C463 ( .A(N204), .B(N205), .Z(N222) );
  GTECH_AND2 C466 ( .A(m5stg_in_of), .B(m5stg_fmuld), .Z(N225) );
  GTECH_OR2 C467 ( .A(N232), .B(m5stg_in_of), .Z(mul_exp_out_in[7]) );
  GTECH_OR2 C468 ( .A(N229), .B(N231), .Z(N232) );
  GTECH_OR2 C469 ( .A(N227), .B(N228), .Z(N229) );
  GTECH_AND2 C470 ( .A(N226), .B(m5stg_exp_plus1[7]), .Z(N227) );
  GTECH_AND2 C471 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N226) );
  GTECH_AND2 C472 ( .A(mul_exp_out_exp), .B(m5stg_exp[7]), .Z(N228) );
  GTECH_AND2 C473 ( .A(N230), .B(m5stg_exp[7]), .Z(N231) );
  GTECH_AND2 C474 ( .A(N204), .B(N205), .Z(N230) );
  GTECH_OR2 C477 ( .A(N239), .B(m5stg_in_of), .Z(mul_exp_out_in[6]) );
  GTECH_OR2 C478 ( .A(N236), .B(N238), .Z(N239) );
  GTECH_OR2 C479 ( .A(N234), .B(N235), .Z(N236) );
  GTECH_AND2 C480 ( .A(N233), .B(m5stg_exp_plus1[6]), .Z(N234) );
  GTECH_AND2 C481 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N233) );
  GTECH_AND2 C482 ( .A(mul_exp_out_exp), .B(m5stg_exp[6]), .Z(N235) );
  GTECH_AND2 C483 ( .A(N237), .B(m5stg_exp[6]), .Z(N238) );
  GTECH_AND2 C484 ( .A(N204), .B(N205), .Z(N237) );
  GTECH_OR2 C487 ( .A(N246), .B(m5stg_in_of), .Z(mul_exp_out_in[5]) );
  GTECH_OR2 C488 ( .A(N243), .B(N245), .Z(N246) );
  GTECH_OR2 C489 ( .A(N241), .B(N242), .Z(N243) );
  GTECH_AND2 C490 ( .A(N240), .B(m5stg_exp_plus1[5]), .Z(N241) );
  GTECH_AND2 C491 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N240) );
  GTECH_AND2 C492 ( .A(mul_exp_out_exp), .B(m5stg_exp[5]), .Z(N242) );
  GTECH_AND2 C493 ( .A(N244), .B(m5stg_exp[5]), .Z(N245) );
  GTECH_AND2 C494 ( .A(N204), .B(N205), .Z(N244) );
  GTECH_OR2 C497 ( .A(N253), .B(m5stg_in_of), .Z(mul_exp_out_in[4]) );
  GTECH_OR2 C498 ( .A(N250), .B(N252), .Z(N253) );
  GTECH_OR2 C499 ( .A(N248), .B(N249), .Z(N250) );
  GTECH_AND2 C500 ( .A(N247), .B(m5stg_exp_plus1[4]), .Z(N248) );
  GTECH_AND2 C501 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N247) );
  GTECH_AND2 C502 ( .A(mul_exp_out_exp), .B(m5stg_exp[4]), .Z(N249) );
  GTECH_AND2 C503 ( .A(N251), .B(m5stg_exp[4]), .Z(N252) );
  GTECH_AND2 C504 ( .A(N204), .B(N205), .Z(N251) );
  GTECH_OR2 C507 ( .A(N260), .B(m5stg_in_of), .Z(mul_exp_out_in[3]) );
  GTECH_OR2 C508 ( .A(N257), .B(N259), .Z(N260) );
  GTECH_OR2 C509 ( .A(N255), .B(N256), .Z(N257) );
  GTECH_AND2 C510 ( .A(N254), .B(m5stg_exp_plus1[3]), .Z(N255) );
  GTECH_AND2 C511 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N254) );
  GTECH_AND2 C512 ( .A(mul_exp_out_exp), .B(m5stg_exp[3]), .Z(N256) );
  GTECH_AND2 C513 ( .A(N258), .B(m5stg_exp[3]), .Z(N259) );
  GTECH_AND2 C514 ( .A(N204), .B(N205), .Z(N258) );
  GTECH_OR2 C517 ( .A(N267), .B(m5stg_in_of), .Z(mul_exp_out_in[2]) );
  GTECH_OR2 C518 ( .A(N264), .B(N266), .Z(N267) );
  GTECH_OR2 C519 ( .A(N262), .B(N263), .Z(N264) );
  GTECH_AND2 C520 ( .A(N261), .B(m5stg_exp_plus1[2]), .Z(N262) );
  GTECH_AND2 C521 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N261) );
  GTECH_AND2 C522 ( .A(mul_exp_out_exp), .B(m5stg_exp[2]), .Z(N263) );
  GTECH_AND2 C523 ( .A(N265), .B(m5stg_exp[2]), .Z(N266) );
  GTECH_AND2 C524 ( .A(N204), .B(N205), .Z(N265) );
  GTECH_OR2 C527 ( .A(N274), .B(m5stg_in_of), .Z(mul_exp_out_in[1]) );
  GTECH_OR2 C528 ( .A(N271), .B(N273), .Z(N274) );
  GTECH_OR2 C529 ( .A(N269), .B(N270), .Z(N271) );
  GTECH_AND2 C530 ( .A(N268), .B(m5stg_exp_plus1[1]), .Z(N269) );
  GTECH_AND2 C531 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N268) );
  GTECH_AND2 C532 ( .A(mul_exp_out_exp), .B(m5stg_exp[1]), .Z(N270) );
  GTECH_AND2 C533 ( .A(N272), .B(m5stg_exp[1]), .Z(N273) );
  GTECH_AND2 C534 ( .A(N204), .B(N205), .Z(N272) );
  GTECH_OR2 C537 ( .A(N281), .B(N282), .Z(mul_exp_out_in[0]) );
  GTECH_OR2 C538 ( .A(N278), .B(N280), .Z(N281) );
  GTECH_OR2 C539 ( .A(N276), .B(N277), .Z(N278) );
  GTECH_AND2 C540 ( .A(N275), .B(m5stg_exp_plus1[0]), .Z(N276) );
  GTECH_AND2 C541 ( .A(mul_exp_out_exp_plus1), .B(m5stg_fracadd_cout), .Z(N275) );
  GTECH_AND2 C542 ( .A(mul_exp_out_exp), .B(m5stg_exp[0]), .Z(N277) );
  GTECH_AND2 C543 ( .A(N279), .B(m5stg_exp[0]), .Z(N280) );
  GTECH_AND2 C544 ( .A(N204), .B(N205), .Z(N279) );
  GTECH_AND2 C547 ( .A(m5stg_in_of), .B(m5stg_to_0_inv), .Z(N282) );
endmodule


module fpu_cnt_lead0_53b ( din, lead0 );
  input [52:0] din;
  output [5:0] lead0;
  wire   din_52_49_eq_0, din_52_51_eq_0, lead0_52_49_0, din_48_45_eq_0,
         din_48_47_eq_0, lead0_48_45_0, din_44_41_eq_0, din_44_43_eq_0,
         lead0_44_41_0, din_40_37_eq_0, din_40_39_eq_0, lead0_40_37_0,
         din_36_33_eq_0, din_36_35_eq_0, lead0_36_33_0, din_32_29_eq_0,
         din_32_31_eq_0, lead0_32_29_0, din_28_25_eq_0, din_28_27_eq_0,
         lead0_28_25_0, din_24_21_eq_0, din_24_23_eq_0, lead0_24_21_0,
         din_20_17_eq_0, din_20_19_eq_0, lead0_20_17_0, din_16_13_eq_0,
         din_16_15_eq_0, lead0_16_13_0, din_12_9_eq_0, din_12_11_eq_0,
         lead0_12_9_0, din_8_5_eq_0, din_8_7_eq_0, lead0_8_5_0, din_4_1_eq_0,
         din_4_3_eq_0, lead0_4_1_0, lead0_0_0, din_52_45_eq_0, lead0_52_45_1,
         lead0_52_45_0, din_44_37_eq_0, lead0_44_37_1, lead0_44_37_0,
         din_36_29_eq_0, lead0_36_29_1, lead0_36_29_0, din_28_21_eq_0,
         lead0_28_21_1, lead0_28_21_0, din_20_13_eq_0, lead0_20_13_1,
         lead0_20_13_0, din_12_5_eq_0, lead0_12_5_1, lead0_12_5_0, lead0_4_0_1,
         lead0_4_0_0, din_52_37_eq_0, lead0_52_37_2, lead0_52_37_1,
         lead0_52_37_0, din_36_21_eq_0, lead0_36_21_2, lead0_36_21_1,
         lead0_36_21_0, din_20_5_eq_0, lead0_20_5_2, lead0_20_5_1,
         lead0_20_5_0, lead0_52_21_3, lead0_52_21_2, lead0_52_21_1,
         lead0_52_21_0, lead0_20_0_3, lead0_20_0_2, lead0_20_0_1, lead0_20_0_0,
         N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14;

  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_52_49 ( .din(din[52:49]), 
        .din_3_0_eq_0(din_52_49_eq_0), .din_3_2_eq_0(din_52_51_eq_0), 
        .lead0_4b_0(lead0_52_49_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_48_45 ( .din(din[48:45]), 
        .din_3_0_eq_0(din_48_45_eq_0), .din_3_2_eq_0(din_48_47_eq_0), 
        .lead0_4b_0(lead0_48_45_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_44_41 ( .din(din[44:41]), 
        .din_3_0_eq_0(din_44_41_eq_0), .din_3_2_eq_0(din_44_43_eq_0), 
        .lead0_4b_0(lead0_44_41_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_40_37 ( .din(din[40:37]), 
        .din_3_0_eq_0(din_40_37_eq_0), .din_3_2_eq_0(din_40_39_eq_0), 
        .lead0_4b_0(lead0_40_37_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_36_33 ( .din(din[36:33]), 
        .din_3_0_eq_0(din_36_33_eq_0), .din_3_2_eq_0(din_36_35_eq_0), 
        .lead0_4b_0(lead0_36_33_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_32_29 ( .din(din[32:29]), 
        .din_3_0_eq_0(din_32_29_eq_0), .din_3_2_eq_0(din_32_31_eq_0), 
        .lead0_4b_0(lead0_32_29_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_28_25 ( .din(din[28:25]), 
        .din_3_0_eq_0(din_28_25_eq_0), .din_3_2_eq_0(din_28_27_eq_0), 
        .lead0_4b_0(lead0_28_25_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_24_21 ( .din(din[24:21]), 
        .din_3_0_eq_0(din_24_21_eq_0), .din_3_2_eq_0(din_24_23_eq_0), 
        .lead0_4b_0(lead0_24_21_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_20_17 ( .din(din[20:17]), 
        .din_3_0_eq_0(din_20_17_eq_0), .din_3_2_eq_0(din_20_19_eq_0), 
        .lead0_4b_0(lead0_20_17_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_16_13 ( .din(din[16:13]), 
        .din_3_0_eq_0(din_16_13_eq_0), .din_3_2_eq_0(din_16_15_eq_0), 
        .lead0_4b_0(lead0_16_13_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_12_9 ( .din(din[12:9]), 
        .din_3_0_eq_0(din_12_9_eq_0), .din_3_2_eq_0(din_12_11_eq_0), 
        .lead0_4b_0(lead0_12_9_0) );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_8_5 ( .din(din[8:5]), .din_3_0_eq_0(
        din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), .lead0_4b_0(lead0_8_5_0)
         );
  fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_4_1 ( .din(din[4:1]), .din_3_0_eq_0(
        din_4_1_eq_0), .din_3_2_eq_0(din_4_3_eq_0), .lead0_4b_0(lead0_4_1_0)
         );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_52_45 ( .din_7_4_eq_0(din_52_49_eq_0), .din_7_6_eq_0(din_52_51_eq_0), .lead0_4b_0_hi(lead0_52_49_0), .din_3_0_eq_0(
        din_48_45_eq_0), .din_3_2_eq_0(din_48_47_eq_0), .lead0_4b_0_lo(
        lead0_48_45_0), .din_7_0_eq_0(din_52_45_eq_0), .lead0_8b_1(
        lead0_52_45_1), .lead0_8b_0(lead0_52_45_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_44_37 ( .din_7_4_eq_0(din_44_41_eq_0), .din_7_6_eq_0(din_44_43_eq_0), .lead0_4b_0_hi(lead0_44_41_0), .din_3_0_eq_0(
        din_40_37_eq_0), .din_3_2_eq_0(din_40_39_eq_0), .lead0_4b_0_lo(
        lead0_40_37_0), .din_7_0_eq_0(din_44_37_eq_0), .lead0_8b_1(
        lead0_44_37_1), .lead0_8b_0(lead0_44_37_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_36_29 ( .din_7_4_eq_0(din_36_33_eq_0), .din_7_6_eq_0(din_36_35_eq_0), .lead0_4b_0_hi(lead0_36_33_0), .din_3_0_eq_0(
        din_32_29_eq_0), .din_3_2_eq_0(din_32_31_eq_0), .lead0_4b_0_lo(
        lead0_32_29_0), .din_7_0_eq_0(din_36_29_eq_0), .lead0_8b_1(
        lead0_36_29_1), .lead0_8b_0(lead0_36_29_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_28_21 ( .din_7_4_eq_0(din_28_25_eq_0), .din_7_6_eq_0(din_28_27_eq_0), .lead0_4b_0_hi(lead0_28_25_0), .din_3_0_eq_0(
        din_24_21_eq_0), .din_3_2_eq_0(din_24_23_eq_0), .lead0_4b_0_lo(
        lead0_24_21_0), .din_7_0_eq_0(din_28_21_eq_0), .lead0_8b_1(
        lead0_28_21_1), .lead0_8b_0(lead0_28_21_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_20_13 ( .din_7_4_eq_0(din_20_17_eq_0), .din_7_6_eq_0(din_20_19_eq_0), .lead0_4b_0_hi(lead0_20_17_0), .din_3_0_eq_0(
        din_16_13_eq_0), .din_3_2_eq_0(din_16_15_eq_0), .lead0_4b_0_lo(
        lead0_16_13_0), .din_7_0_eq_0(din_20_13_eq_0), .lead0_8b_1(
        lead0_20_13_1), .lead0_8b_0(lead0_20_13_0) );
  fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_12_5 ( .din_7_4_eq_0(din_12_9_eq_0), 
        .din_7_6_eq_0(din_12_11_eq_0), .lead0_4b_0_hi(lead0_12_9_0), 
        .din_3_0_eq_0(din_8_5_eq_0), .din_3_2_eq_0(din_8_7_eq_0), 
        .lead0_4b_0_lo(lead0_8_5_0), .din_7_0_eq_0(din_12_5_eq_0), 
        .lead0_8b_1(lead0_12_5_1), .lead0_8b_0(lead0_12_5_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_52_37 ( .din_15_8_eq_0(
        din_52_45_eq_0), .din_15_12_eq_0(din_52_49_eq_0), .lead0_8b_1_hi(
        lead0_52_45_1), .lead0_8b_0_hi(lead0_52_45_0), .din_7_0_eq_0(
        din_44_37_eq_0), .din_7_4_eq_0(din_44_41_eq_0), .lead0_8b_1_lo(
        lead0_44_37_1), .lead0_8b_0_lo(lead0_44_37_0), .din_15_0_eq_0(
        din_52_37_eq_0), .lead0_16b_2(lead0_52_37_2), .lead0_16b_1(
        lead0_52_37_1), .lead0_16b_0(lead0_52_37_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_36_21 ( .din_15_8_eq_0(
        din_36_29_eq_0), .din_15_12_eq_0(din_36_33_eq_0), .lead0_8b_1_hi(
        lead0_36_29_1), .lead0_8b_0_hi(lead0_36_29_0), .din_7_0_eq_0(
        din_28_21_eq_0), .din_7_4_eq_0(din_28_25_eq_0), .lead0_8b_1_lo(
        lead0_28_21_1), .lead0_8b_0_lo(lead0_28_21_0), .din_15_0_eq_0(
        din_36_21_eq_0), .lead0_16b_2(lead0_36_21_2), .lead0_16b_1(
        lead0_36_21_1), .lead0_16b_0(lead0_36_21_0) );
  fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_20_5 ( .din_15_8_eq_0(din_20_13_eq_0), .din_15_12_eq_0(din_20_17_eq_0), .lead0_8b_1_hi(lead0_20_13_1), 
        .lead0_8b_0_hi(lead0_20_13_0), .din_7_0_eq_0(din_12_5_eq_0), 
        .din_7_4_eq_0(din_12_9_eq_0), .lead0_8b_1_lo(lead0_12_5_1), 
        .lead0_8b_0_lo(lead0_12_5_0), .din_15_0_eq_0(din_20_5_eq_0), 
        .lead0_16b_2(lead0_20_5_2), .lead0_16b_1(lead0_20_5_1), .lead0_16b_0(
        lead0_20_5_0) );
  fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_52_21 ( .din_31_16_eq_0(
        din_52_37_eq_0), .din_31_24_eq_0(din_52_45_eq_0), .lead0_16b_2_hi(
        lead0_52_37_2), .lead0_16b_1_hi(lead0_52_37_1), .lead0_16b_0_hi(
        lead0_52_37_0), .din_15_0_eq_0(din_36_21_eq_0), .din_15_8_eq_0(
        din_36_29_eq_0), .lead0_16b_2_lo(lead0_36_21_2), .lead0_16b_1_lo(
        lead0_36_21_1), .lead0_16b_0_lo(lead0_36_21_0), .din_31_0_eq_0(
        lead0[5]), .lead0_32b_3(lead0_52_21_3), .lead0_32b_2(lead0_52_21_2), 
        .lead0_32b_1(lead0_52_21_1), .lead0_32b_0(lead0_52_21_0) );
  fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_20_0 ( .din_31_16_eq_0(din_20_5_eq_0), .din_31_24_eq_0(din_20_13_eq_0), .lead0_16b_2_hi(lead0_20_5_2), 
        .lead0_16b_1_hi(lead0_20_5_1), .lead0_16b_0_hi(lead0_20_5_0), 
        .din_15_0_eq_0(1'b0), .din_15_8_eq_0(1'b0), .lead0_16b_2_lo(
        din_4_1_eq_0), .lead0_16b_1_lo(lead0_4_0_1), .lead0_16b_0_lo(
        lead0_4_0_0), .lead0_32b_3(lead0_20_0_3), .lead0_32b_2(lead0_20_0_2), 
        .lead0_32b_1(lead0_20_0_1), .lead0_32b_0(lead0_20_0_0) );
  GTECH_NOT I_0 ( .A(din[0]), .Z(lead0_0_0) );
  GTECH_AND2 C16 ( .A(N0), .B(din_4_3_eq_0), .Z(lead0_4_0_1) );
  GTECH_NOT I_1 ( .A(din_4_1_eq_0), .Z(N0) );
  GTECH_OR2 C18 ( .A(N2), .B(N3), .Z(lead0_4_0_0) );
  GTECH_AND2 C19 ( .A(N1), .B(lead0_4_1_0), .Z(N2) );
  GTECH_NOT I_2 ( .A(din_4_1_eq_0), .Z(N1) );
  GTECH_AND2 C21 ( .A(din_4_1_eq_0), .B(lead0_0_0), .Z(N3) );
  GTECH_OR2 C22 ( .A(N5), .B(N6), .Z(lead0[4]) );
  GTECH_AND2 C23 ( .A(N4), .B(din_52_37_eq_0), .Z(N5) );
  GTECH_NOT I_3 ( .A(lead0[5]), .Z(N4) );
  GTECH_AND2 C25 ( .A(lead0[5]), .B(din_20_5_eq_0), .Z(N6) );
  GTECH_OR2 C26 ( .A(N7), .B(N8), .Z(lead0[3]) );
  GTECH_AND2 C27 ( .A(N4), .B(lead0_52_21_3), .Z(N7) );
  GTECH_AND2 C29 ( .A(lead0[5]), .B(lead0_20_0_3), .Z(N8) );
  GTECH_OR2 C30 ( .A(N9), .B(N10), .Z(lead0[2]) );
  GTECH_AND2 C31 ( .A(N4), .B(lead0_52_21_2), .Z(N9) );
  GTECH_AND2 C33 ( .A(lead0[5]), .B(lead0_20_0_2), .Z(N10) );
  GTECH_OR2 C34 ( .A(N11), .B(N12), .Z(lead0[1]) );
  GTECH_AND2 C35 ( .A(N4), .B(lead0_52_21_1), .Z(N11) );
  GTECH_AND2 C37 ( .A(lead0[5]), .B(lead0_20_0_1), .Z(N12) );
  GTECH_OR2 C38 ( .A(N13), .B(N14), .Z(lead0[0]) );
  GTECH_AND2 C39 ( .A(N4), .B(lead0_52_21_0), .Z(N13) );
  GTECH_AND2 C41 ( .A(lead0[5]), .B(lead0_20_0_0), .Z(N14) );
endmodule


module dffe_SIZE56 ( din, en, clk, q, se, si, so );
  input [55:0] din;
  output [55:0] q;
  input [55:0] si;
  output [55:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61;
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N61) );
  SELECT_OP C239 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C247 ( .A(N3), .B(N2), .Z(N60) );
  GTECH_NOT I_2 ( .A(N60), .Z(N61) );
endmodule


module dff_SIZE55 ( din, clk, q, se, si, so );
  input [54:0] din;
  output [54:0] q;
  input [54:0] si;
  output [54:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57;
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C65 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dffe_SIZE52 ( din, en, clk, q, se, si, so );
  input [51:0] din;
  output [51:0] q;
  input [51:0] si;
  output [51:0] so;
  input en, clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57;
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N57) );
  SELECT_OP C223 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
  GTECH_NOT I_1 ( .A(en), .Z(N3) );
  GTECH_AND2 C231 ( .A(N3), .B(N2), .Z(N56) );
  GTECH_NOT I_2 ( .A(N56), .Z(N57) );
endmodule


module fpu_mul_frac_dp ( inq_in1, inq_in2, m6stg_step, m2stg_frac1_dbl_norm, 
        m2stg_frac1_dbl_dnrm, m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, 
        m2stg_frac1_inf, m1stg_snan_dbl_in1, m1stg_snan_sng_in1, 
        m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, 
        m2stg_frac2_sng_dnrm, m2stg_frac2_inf, m1stg_snan_dbl_in2, 
        m1stg_snan_sng_in2, m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, 
        m1stg_dblop, m1stg_dblop_inv, m4stg_frac, m4stg_sh_cnt_in, 
        m3bstg_ld0_inv, m4stg_left_shift_step, m4stg_right_shift_step, 
        m5stg_fmuls, m5stg_fmulda, mul_frac_out_fracadd, mul_frac_out_frac, 
        m5stg_in_of, m5stg_to_0, fmul_clken_l, rclk, m2stg_frac1_array_in, 
        m2stg_frac2_array_in, m1stg_ld0_1, m1stg_ld0_2, m4stg_frac_105, 
        m3stg_ld0_inv, m4stg_shl_54, m4stg_shl_55, m5stg_frac_32_0, 
        m5stg_frac_dbl_nx, m5stg_frac_sng_nx, m5stg_frac_neq_0, 
        m5stg_fracadd_cout, mul_frac_out, se, si, so );
  input [54:0] inq_in1;
  input [54:0] inq_in2;
  input [105:0] m4stg_frac;
  input [5:0] m4stg_sh_cnt_in;
  input [6:0] m3bstg_ld0_inv;
  output [52:0] m2stg_frac1_array_in;
  output [52:0] m2stg_frac2_array_in;
  output [5:0] m1stg_ld0_1;
  output [5:0] m1stg_ld0_2;
  output [6:0] m3stg_ld0_inv;
  output [32:0] m5stg_frac_32_0;
  output [51:0] mul_frac_out;
  input m6stg_step, m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm,
         m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, m2stg_frac1_inf,
         m1stg_snan_dbl_in1, m1stg_snan_sng_in1, m2stg_frac2_dbl_norm,
         m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm, m2stg_frac2_sng_dnrm,
         m2stg_frac2_inf, m1stg_snan_dbl_in2, m1stg_snan_sng_in2,
         m1stg_inf_zero_in, m1stg_inf_zero_in_dbl, m1stg_dblop,
         m1stg_dblop_inv, m4stg_left_shift_step, m4stg_right_shift_step,
         m5stg_fmuls, m5stg_fmulda, mul_frac_out_fracadd, mul_frac_out_frac,
         m5stg_in_of, m5stg_to_0, fmul_clken_l, rclk, se, si;
  output m4stg_frac_105, m4stg_shl_54, m4stg_shl_55, m5stg_frac_dbl_nx,
         m5stg_frac_sng_nx, m5stg_frac_neq_0, m5stg_fracadd_cout, so;
  wire   se_l, clk, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13,
         N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285,
         N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296,
         N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307,
         N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318,
         N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329,
         N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340,
         N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351,
         N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362,
         N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384,
         N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417,
         N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450,
         N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483,
         N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516,
         N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
         N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538,
         N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604,
         N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648,
         N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714,
         N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725,
         N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901,
         N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020,
         N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030,
         N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040,
         N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050,
         N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060,
         N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070,
         N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080,
         N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090,
         N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100,
         N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110,
         N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120,
         N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130,
         N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140,
         N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150,
         N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160,
         N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170,
         N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180,
         N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190,
         N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200,
         N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210,
         N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220,
         N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230,
         N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240,
         N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250,
         N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260,
         N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270,
         N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280,
         N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290,
         N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300,
         N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310,
         N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320,
         N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330,
         N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340,
         N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350,
         N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370,
         N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380,
         N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390,
         N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400,
         N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410,
         N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420,
         N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430,
         N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440,
         N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470,
         N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480,
         N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490,
         N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500,
         N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510,
         N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, N1519, N1520,
         N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530,
         N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540,
         N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550,
         N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560,
         N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570,
         N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580,
         N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590,
         N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600,
         N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610,
         N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620,
         N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630,
         N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640,
         N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650,
         N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660,
         N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670,
         N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680,
         N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690,
         N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700,
         N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710,
         N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720,
         N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730,
         N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740,
         N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750,
         N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760,
         N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770,
         N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780,
         N1781, net13855, net13856, net13857, net13858, net13859, net13860,
         net13861, net13862, net13863, net13864, net13865, net13866, net13867,
         net13868, net13869, net13870, net13871, net13872, net13873, net13874,
         net13875, net13876, net13877, net13878, net13879, net13880, net13881,
         net13882, net13883, net13884, net13885, net13886, net13887, net13888,
         net13889, net13890, net13891, net13892, net13893, net13894, net13895,
         net13896, net13897, net13898, net13899, net13900, net13901, net13902,
         net13903, net13904, net13905, net13906, net13907, net13908, net13909,
         net13910, net13911, net13912, net13913, net13914, net13915, net13916,
         net13917, net13918, net13919, net13920, net13921, net13922, net13923,
         net13924, net13925, net13926, net13927, net13928, net13929, net13930,
         net13931, net13932, net13933, net13934, net13935, net13936, net13937,
         net13938, net13939, net13940, net13941, net13942, net13943, net13944,
         net13945, net13946, net13947, net13948, net13949, net13950, net13951,
         net13952, net13953, net13954, net13955, net13956, net13957, net13958,
         net13959, net13960, net13961, net13962, net13963, net13964, net13965,
         net13966, net13967, net13968, net13969, net13970, net13971, net13972,
         net13973, net13974, net13975, net13976, net13977, net13978, net13979,
         net13980, net13981, net13982, net13983, net13984, net13985, net13986,
         net13987, net13988, net13989, net13990, net13991, net13992, net13993,
         net13994, net13995, net13996, net13997, net13998, net13999, net14000,
         net14001, net14002, net14003, net14004, net14005, net14006, net14007,
         net14008, net14009, net14010, net14011, net14012, net14013, net14014,
         net14015, net14016, net14017, net14018, net14019, net14020, net14021,
         net14022, net14023, net14024, net14025, net14026, net14027, net14028,
         net14029, net14030, net14031, net14032, net14033, net14034, net14035,
         net14036, net14037, net14038, net14039, net14040, net14041, net14042,
         net14043, net14044, net14045, net14046, net14047, net14048, net14049,
         net14050, net14051, net14052, net14053, net14054, net14055, net14056,
         net14057, net14058, net14059, net14060, net14061, net14062, net14063,
         net14064, net14065, net14066, net14067, net14068, net14069, net14070,
         net14071, net14072, net14073, net14074, net14075, net14076, net14077,
         net14078, net14079, net14080, net14081, net14082, net14083, net14084,
         net14085, net14086, net14087, net14088, net14089, net14090, net14091,
         net14092, net14093, net14094, net14095, net14096, net14097, net14098,
         net14099, net14100, net14101, net14102, net14103, net14104, net14105,
         net14106, net14107, net14108, net14109, net14110, net14111, net14112,
         net14113, net14114, net14115, net14116, net14117, net14118, net14119,
         net14120, net14121, net14122, net14123, net14124, net14125, net14126,
         net14127, net14128, net14129, net14130, net14131, net14132, net14133,
         net14134, net14135, net14136, net14137, net14138, net14139, net14140,
         net14141, net14142, net14143, net14144, net14145, net14146, net14147,
         net14148, net14149, net14150, net14151, net14152, net14153, net14154,
         net14155, net14156, net14157, net14158, net14159, net14160, net14161,
         net14162, net14163, net14164, net14165, net14166, net14167, net14168,
         net14169, net14170, net14171, net14172, net14173, net14174, net14175,
         net14176, net14177, net14178, net14179, net14180, net14181, net14182,
         net14183, net14184, net14185, net14186, net14187, net14188, net14189,
         net14190, net14191, net14192, net14193, net14194, net14195, net14196,
         net14197, net14198, net14199, net14200, net14201, net14202, net14203,
         net14204, net14205, net14206, net14207, net14208, net14209, net14210,
         net14211, net14212, net14213, net14214, net14215, net14216, net14217,
         net14218, net14219, net14220, net14221, net14222, net14223, net14224,
         net14225, net14226, net14227, net14228, net14229, net14230, net14231,
         net14232, net14233, net14234, net14235, net14236, net14237, net14238,
         net14239, net14240, net14241, net14242, net14243, net14244, net14245,
         net14246, net14247, net14248, net14249, net14250, net14251, net14252,
         net14253, net14254, net14255, net14256, net14257, net14258, net14259,
         net14260, net14261, net14262, net14263, net14264, net14265, net14266,
         net14267, net14268, net14269, net14270, net14271, net14272, net14273,
         net14274, net14275, net14276, net14277, net14278, net14279, net14280,
         net14281, net14282, net14283, net14284, net14285, net14286, net14287,
         net14288, net14289, net14290, net14291, net14292, net14293;
  wire   [54:0] mul_frac_in1;
  wire   [54:0] mul_frac_in2;
  wire   [52:0] m2stg_frac1_in;
  wire   [52:1] m1stg_ld0_1_din;
  wire   [52:1] m1stg_ld0_2_din;
  wire   [5:0] m4stg_sh_cnt_5;
  wire   [5:0] m4stg_sh_cnt_4;
  wire   [5:0] m4stg_sh_cnt;
  wire   [30:0] mstg_xtra_regs;
  wire   [166:63] m4stg_shl_tmp;
  wire   [0:0] m4stg_shl;
  wire   [168:0] m4stg_shr_tmp;
  wire   [0:0] m4stg_shr;
  wire   [54:0] m5stg_frac_pre1_in;
  wire   [54:0] m5stg_frac_pre1;
  wire   [54:1] m5stg_frac_pre2_in;
  wire   [54:0] m5stg_frac_pre2;
  wire   [54:0] m5stg_frac_pre3_in;
  wire   [54:0] m5stg_frac_pre3;
  wire   [54:1] m5stg_frac_pre4_in;
  wire   [54:0] m5stg_frac_pre4;
  wire   [54:33] m5stg_frac_54_33;
  wire   [51:0] m5stg_fracadd_tmp;
  wire   [51:0] mul_frac_out_in;
  assign m4stg_frac_105 = m4stg_frac[105];

  clken_buf ckbuf_mul_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fmul_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE55 i_mul_frac_in1 ( .din(inq_in1), .en(m6stg_step), .clk(clk), .q(
        mul_frac_in1), .se(se), .si({net14239, net14240, net14241, net14242, 
        net14243, net14244, net14245, net14246, net14247, net14248, net14249, 
        net14250, net14251, net14252, net14253, net14254, net14255, net14256, 
        net14257, net14258, net14259, net14260, net14261, net14262, net14263, 
        net14264, net14265, net14266, net14267, net14268, net14269, net14270, 
        net14271, net14272, net14273, net14274, net14275, net14276, net14277, 
        net14278, net14279, net14280, net14281, net14282, net14283, net14284, 
        net14285, net14286, net14287, net14288, net14289, net14290, net14291, 
        net14292, net14293}) );
  dffe_SIZE55 i_mul_frac_in2 ( .din(inq_in2), .en(m6stg_step), .clk(clk), .q(
        mul_frac_in2), .se(se), .si({net14184, net14185, net14186, net14187, 
        net14188, net14189, net14190, net14191, net14192, net14193, net14194, 
        net14195, net14196, net14197, net14198, net14199, net14200, net14201, 
        net14202, net14203, net14204, net14205, net14206, net14207, net14208, 
        net14209, net14210, net14211, net14212, net14213, net14214, net14215, 
        net14216, net14217, net14218, net14219, net14220, net14221, net14222, 
        net14223, net14224, net14225, net14226, net14227, net14228, net14229, 
        net14230, net14231, net14232, net14233, net14234, net14235, net14236, 
        net14237, net14238}) );
  fpu_cnt_lead0_53b i_m1stg_ld0_1 ( .din({m1stg_ld0_1_din, 1'b0}), .lead0(
        m1stg_ld0_1) );
  fpu_cnt_lead0_53b i_m1stg_ld0_2 ( .din({m1stg_ld0_2_din, 1'b0}), .lead0(
        m1stg_ld0_2) );
  dffe_SIZE56 i_mstg_xtra_regs ( .din({m4stg_sh_cnt_in[5], m4stg_sh_cnt_in[5], 
        m4stg_sh_cnt_in[5], m4stg_sh_cnt_in[5], m4stg_sh_cnt_in[5], 
        m4stg_sh_cnt_in[5:4], m4stg_sh_cnt_in[4], m4stg_sh_cnt_in[4], 
        m4stg_sh_cnt_in[4], m4stg_sh_cnt_in[4], m4stg_sh_cnt_in[4], 
        m4stg_sh_cnt_in[5], m4stg_sh_cnt_in[4:0], m3bstg_ld0_inv, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .en(m6stg_step), .clk(clk), .q({
        m4stg_sh_cnt_5, m4stg_sh_cnt_4, m4stg_sh_cnt, m3stg_ld0_inv, 
        mstg_xtra_regs}), .se(se), .si({net14128, net14129, net14130, net14131, 
        net14132, net14133, net14134, net14135, net14136, net14137, net14138, 
        net14139, net14140, net14141, net14142, net14143, net14144, net14145, 
        net14146, net14147, net14148, net14149, net14150, net14151, net14152, 
        net14153, net14154, net14155, net14156, net14157, net14158, net14159, 
        net14160, net14161, net14162, net14163, net14164, net14165, net14166, 
        net14167, net14168, net14169, net14170, net14171, net14172, net14173, 
        net14174, net14175, net14176, net14177, net14178, net14179, net14180, 
        net14181, net14182, net14183}) );
  ASH_UNS_UNS_OP sll_334 ( .A(m4stg_frac), .SH({m4stg_sh_cnt_5[0], 
        m4stg_sh_cnt[4:0]}), .Z({m4stg_shl_55, m4stg_shl_54, m4stg_shl_tmp})
         );
  ASHR_UNS_UNS_OP srl_348 ( .A({m4stg_frac, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SH(
        m4stg_sh_cnt), .Z(m4stg_shr_tmp) );
  dff_SIZE55 i_m5stg_frac_pre1 ( .din(m5stg_frac_pre1_in), .clk(clk), .q(
        m5stg_frac_pre1), .se(se), .si({net14073, net14074, net14075, net14076, 
        net14077, net14078, net14079, net14080, net14081, net14082, net14083, 
        net14084, net14085, net14086, net14087, net14088, net14089, net14090, 
        net14091, net14092, net14093, net14094, net14095, net14096, net14097, 
        net14098, net14099, net14100, net14101, net14102, net14103, net14104, 
        net14105, net14106, net14107, net14108, net14109, net14110, net14111, 
        net14112, net14113, net14114, net14115, net14116, net14117, net14118, 
        net14119, net14120, net14121, net14122, net14123, net14124, net14125, 
        net14126, net14127}) );
  dff_SIZE55 i_m5stg_frac_pre2 ( .din({m5stg_frac_pre2_in, 1'b1}), .clk(clk), 
        .q(m5stg_frac_pre2), .se(se), .si({net14018, net14019, net14020, 
        net14021, net14022, net14023, net14024, net14025, net14026, net14027, 
        net14028, net14029, net14030, net14031, net14032, net14033, net14034, 
        net14035, net14036, net14037, net14038, net14039, net14040, net14041, 
        net14042, net14043, net14044, net14045, net14046, net14047, net14048, 
        net14049, net14050, net14051, net14052, net14053, net14054, net14055, 
        net14056, net14057, net14058, net14059, net14060, net14061, net14062, 
        net14063, net14064, net14065, net14066, net14067, net14068, net14069, 
        net14070, net14071, net14072}) );
  dff_SIZE55 i_m5stg_frac_pre3 ( .din(m5stg_frac_pre3_in), .clk(clk), .q(
        m5stg_frac_pre3), .se(se), .si({net13963, net13964, net13965, net13966, 
        net13967, net13968, net13969, net13970, net13971, net13972, net13973, 
        net13974, net13975, net13976, net13977, net13978, net13979, net13980, 
        net13981, net13982, net13983, net13984, net13985, net13986, net13987, 
        net13988, net13989, net13990, net13991, net13992, net13993, net13994, 
        net13995, net13996, net13997, net13998, net13999, net14000, net14001, 
        net14002, net14003, net14004, net14005, net14006, net14007, net14008, 
        net14009, net14010, net14011, net14012, net14013, net14014, net14015, 
        net14016, net14017}) );
  dff_SIZE55 i_m5stg_frac_pre4 ( .din({m5stg_frac_pre4_in, 1'b1}), .clk(clk), 
        .q(m5stg_frac_pre4), .se(se), .si({net13908, net13909, net13910, 
        net13911, net13912, net13913, net13914, net13915, net13916, net13917, 
        net13918, net13919, net13920, net13921, net13922, net13923, net13924, 
        net13925, net13926, net13927, net13928, net13929, net13930, net13931, 
        net13932, net13933, net13934, net13935, net13936, net13937, net13938, 
        net13939, net13940, net13941, net13942, net13943, net13944, net13945, 
        net13946, net13947, net13948, net13949, net13950, net13951, net13952, 
        net13953, net13954, net13955, net13956, net13957, net13958, net13959, 
        net13960, net13961, net13962}) );
  dffe_SIZE52 i_mul_frac_out ( .din(mul_frac_out_in), .en(m6stg_step), .clk(
        clk), .q(mul_frac_out), .se(se), .si({net13856, net13857, net13858, 
        net13859, net13860, net13861, net13862, net13863, net13864, net13865, 
        net13866, net13867, net13868, net13869, net13870, net13871, net13872, 
        net13873, net13874, net13875, net13876, net13877, net13878, net13879, 
        net13880, net13881, net13882, net13883, net13884, net13885, net13886, 
        net13887, net13888, net13889, net13890, net13891, net13892, net13893, 
        net13894, net13895, net13896, net13897, net13898, net13899, net13900, 
        net13901, net13902, net13903, net13904, net13905, net13906, net13907})
         );
  ADD_UNS_OP add_476 ( .A({m5stg_frac_54_33, m5stg_frac_32_0[32:3]}), .B({
        m5stg_fmuls, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m5stg_fmulda}), .Z({
        m5stg_fracadd_cout, m5stg_fracadd_tmp}) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_OR2 C602 ( .A(N4), .B(m2stg_frac1_inf), .Z(m2stg_frac1_in[52]) );
  GTECH_OR2 C603 ( .A(N2), .B(N3), .Z(N4) );
  GTECH_OR2 C604 ( .A(N1), .B(m2stg_frac1_sng_norm), .Z(N2) );
  GTECH_OR2 C605 ( .A(m2stg_frac1_dbl_norm), .B(N0), .Z(N1) );
  GTECH_AND2 C606 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[51]), .Z(N0) );
  GTECH_AND2 C607 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[54]), .Z(N3) );
  GTECH_OR2 C608 ( .A(N11), .B(N12), .Z(m2stg_frac1_in[51]) );
  GTECH_OR2 C609 ( .A(N8), .B(N10), .Z(N11) );
  GTECH_OR2 C610 ( .A(N6), .B(N7), .Z(N8) );
  GTECH_AND2 C611 ( .A(m2stg_frac1_dbl_norm), .B(N5), .Z(N6) );
  GTECH_OR2 C612 ( .A(mul_frac_in1[51]), .B(m1stg_snan_dbl_in1), .Z(N5) );
  GTECH_AND2 C613 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[50]), .Z(N7) );
  GTECH_AND2 C614 ( .A(m2stg_frac1_sng_norm), .B(N9), .Z(N10) );
  GTECH_OR2 C615 ( .A(mul_frac_in1[54]), .B(m1stg_snan_sng_in1), .Z(N9) );
  GTECH_AND2 C616 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[53]), .Z(N12) );
  GTECH_OR2 C617 ( .A(N17), .B(N18), .Z(m2stg_frac1_in[50]) );
  GTECH_OR2 C618 ( .A(N15), .B(N16), .Z(N17) );
  GTECH_OR2 C619 ( .A(N13), .B(N14), .Z(N15) );
  GTECH_AND2 C620 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[50]), .Z(N13) );
  GTECH_AND2 C621 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[49]), .Z(N14) );
  GTECH_AND2 C622 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[53]), .Z(N16) );
  GTECH_AND2 C623 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[52]), .Z(N18) );
  GTECH_OR2 C624 ( .A(N23), .B(N24), .Z(m2stg_frac1_in[49]) );
  GTECH_OR2 C625 ( .A(N21), .B(N22), .Z(N23) );
  GTECH_OR2 C626 ( .A(N19), .B(N20), .Z(N21) );
  GTECH_AND2 C627 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[49]), .Z(N19) );
  GTECH_AND2 C628 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[48]), .Z(N20) );
  GTECH_AND2 C629 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[52]), .Z(N22) );
  GTECH_AND2 C630 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[51]), .Z(N24) );
  GTECH_OR2 C631 ( .A(N29), .B(N30), .Z(m2stg_frac1_in[48]) );
  GTECH_OR2 C632 ( .A(N27), .B(N28), .Z(N29) );
  GTECH_OR2 C633 ( .A(N25), .B(N26), .Z(N27) );
  GTECH_AND2 C634 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[48]), .Z(N25) );
  GTECH_AND2 C635 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[47]), .Z(N26) );
  GTECH_AND2 C636 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[51]), .Z(N28) );
  GTECH_AND2 C637 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[50]), .Z(N30) );
  GTECH_OR2 C638 ( .A(N35), .B(N36), .Z(m2stg_frac1_in[47]) );
  GTECH_OR2 C639 ( .A(N33), .B(N34), .Z(N35) );
  GTECH_OR2 C640 ( .A(N31), .B(N32), .Z(N33) );
  GTECH_AND2 C641 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[47]), .Z(N31) );
  GTECH_AND2 C642 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[46]), .Z(N32) );
  GTECH_AND2 C643 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[50]), .Z(N34) );
  GTECH_AND2 C644 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[49]), .Z(N36) );
  GTECH_OR2 C645 ( .A(N41), .B(N42), .Z(m2stg_frac1_in[46]) );
  GTECH_OR2 C646 ( .A(N39), .B(N40), .Z(N41) );
  GTECH_OR2 C647 ( .A(N37), .B(N38), .Z(N39) );
  GTECH_AND2 C648 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[46]), .Z(N37) );
  GTECH_AND2 C649 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[45]), .Z(N38) );
  GTECH_AND2 C650 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[49]), .Z(N40) );
  GTECH_AND2 C651 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[48]), .Z(N42) );
  GTECH_OR2 C652 ( .A(N47), .B(N48), .Z(m2stg_frac1_in[45]) );
  GTECH_OR2 C653 ( .A(N45), .B(N46), .Z(N47) );
  GTECH_OR2 C654 ( .A(N43), .B(N44), .Z(N45) );
  GTECH_AND2 C655 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[45]), .Z(N43) );
  GTECH_AND2 C656 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[44]), .Z(N44) );
  GTECH_AND2 C657 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[48]), .Z(N46) );
  GTECH_AND2 C658 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[47]), .Z(N48) );
  GTECH_OR2 C659 ( .A(N53), .B(N54), .Z(m2stg_frac1_in[44]) );
  GTECH_OR2 C660 ( .A(N51), .B(N52), .Z(N53) );
  GTECH_OR2 C661 ( .A(N49), .B(N50), .Z(N51) );
  GTECH_AND2 C662 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[44]), .Z(N49) );
  GTECH_AND2 C663 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[43]), .Z(N50) );
  GTECH_AND2 C664 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[47]), .Z(N52) );
  GTECH_AND2 C665 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[46]), .Z(N54) );
  GTECH_OR2 C666 ( .A(N59), .B(N60), .Z(m2stg_frac1_in[43]) );
  GTECH_OR2 C667 ( .A(N57), .B(N58), .Z(N59) );
  GTECH_OR2 C668 ( .A(N55), .B(N56), .Z(N57) );
  GTECH_AND2 C669 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[43]), .Z(N55) );
  GTECH_AND2 C670 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[42]), .Z(N56) );
  GTECH_AND2 C671 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[46]), .Z(N58) );
  GTECH_AND2 C672 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[45]), .Z(N60) );
  GTECH_OR2 C673 ( .A(N65), .B(N66), .Z(m2stg_frac1_in[42]) );
  GTECH_OR2 C674 ( .A(N63), .B(N64), .Z(N65) );
  GTECH_OR2 C675 ( .A(N61), .B(N62), .Z(N63) );
  GTECH_AND2 C676 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[42]), .Z(N61) );
  GTECH_AND2 C677 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[41]), .Z(N62) );
  GTECH_AND2 C678 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[45]), .Z(N64) );
  GTECH_AND2 C679 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[44]), .Z(N66) );
  GTECH_OR2 C680 ( .A(N71), .B(N72), .Z(m2stg_frac1_in[41]) );
  GTECH_OR2 C681 ( .A(N69), .B(N70), .Z(N71) );
  GTECH_OR2 C682 ( .A(N67), .B(N68), .Z(N69) );
  GTECH_AND2 C683 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[41]), .Z(N67) );
  GTECH_AND2 C684 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[40]), .Z(N68) );
  GTECH_AND2 C685 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[44]), .Z(N70) );
  GTECH_AND2 C686 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[43]), .Z(N72) );
  GTECH_OR2 C687 ( .A(N77), .B(N78), .Z(m2stg_frac1_in[40]) );
  GTECH_OR2 C688 ( .A(N75), .B(N76), .Z(N77) );
  GTECH_OR2 C689 ( .A(N73), .B(N74), .Z(N75) );
  GTECH_AND2 C690 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[40]), .Z(N73) );
  GTECH_AND2 C691 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[39]), .Z(N74) );
  GTECH_AND2 C692 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[43]), .Z(N76) );
  GTECH_AND2 C693 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[42]), .Z(N78) );
  GTECH_OR2 C694 ( .A(N83), .B(N84), .Z(m2stg_frac1_in[39]) );
  GTECH_OR2 C695 ( .A(N81), .B(N82), .Z(N83) );
  GTECH_OR2 C696 ( .A(N79), .B(N80), .Z(N81) );
  GTECH_AND2 C697 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[39]), .Z(N79) );
  GTECH_AND2 C698 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[38]), .Z(N80) );
  GTECH_AND2 C699 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[42]), .Z(N82) );
  GTECH_AND2 C700 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[41]), .Z(N84) );
  GTECH_OR2 C701 ( .A(N89), .B(N90), .Z(m2stg_frac1_in[38]) );
  GTECH_OR2 C702 ( .A(N87), .B(N88), .Z(N89) );
  GTECH_OR2 C703 ( .A(N85), .B(N86), .Z(N87) );
  GTECH_AND2 C704 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[38]), .Z(N85) );
  GTECH_AND2 C705 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[37]), .Z(N86) );
  GTECH_AND2 C706 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[41]), .Z(N88) );
  GTECH_AND2 C707 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[40]), .Z(N90) );
  GTECH_OR2 C708 ( .A(N95), .B(N96), .Z(m2stg_frac1_in[37]) );
  GTECH_OR2 C709 ( .A(N93), .B(N94), .Z(N95) );
  GTECH_OR2 C710 ( .A(N91), .B(N92), .Z(N93) );
  GTECH_AND2 C711 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[37]), .Z(N91) );
  GTECH_AND2 C712 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[36]), .Z(N92) );
  GTECH_AND2 C713 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[40]), .Z(N94) );
  GTECH_AND2 C714 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[39]), .Z(N96) );
  GTECH_OR2 C715 ( .A(N101), .B(N102), .Z(m2stg_frac1_in[36]) );
  GTECH_OR2 C716 ( .A(N99), .B(N100), .Z(N101) );
  GTECH_OR2 C717 ( .A(N97), .B(N98), .Z(N99) );
  GTECH_AND2 C718 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[36]), .Z(N97) );
  GTECH_AND2 C719 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[35]), .Z(N98) );
  GTECH_AND2 C720 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[39]), .Z(N100)
         );
  GTECH_AND2 C721 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[38]), .Z(N102)
         );
  GTECH_OR2 C722 ( .A(N107), .B(N108), .Z(m2stg_frac1_in[35]) );
  GTECH_OR2 C723 ( .A(N105), .B(N106), .Z(N107) );
  GTECH_OR2 C724 ( .A(N103), .B(N104), .Z(N105) );
  GTECH_AND2 C725 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[35]), .Z(N103)
         );
  GTECH_AND2 C726 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[34]), .Z(N104)
         );
  GTECH_AND2 C727 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[38]), .Z(N106)
         );
  GTECH_AND2 C728 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[37]), .Z(N108)
         );
  GTECH_OR2 C729 ( .A(N113), .B(N114), .Z(m2stg_frac1_in[34]) );
  GTECH_OR2 C730 ( .A(N111), .B(N112), .Z(N113) );
  GTECH_OR2 C731 ( .A(N109), .B(N110), .Z(N111) );
  GTECH_AND2 C732 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[34]), .Z(N109)
         );
  GTECH_AND2 C733 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[33]), .Z(N110)
         );
  GTECH_AND2 C734 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[37]), .Z(N112)
         );
  GTECH_AND2 C735 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[36]), .Z(N114)
         );
  GTECH_OR2 C736 ( .A(N119), .B(N120), .Z(m2stg_frac1_in[33]) );
  GTECH_OR2 C737 ( .A(N117), .B(N118), .Z(N119) );
  GTECH_OR2 C738 ( .A(N115), .B(N116), .Z(N117) );
  GTECH_AND2 C739 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[33]), .Z(N115)
         );
  GTECH_AND2 C740 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[32]), .Z(N116)
         );
  GTECH_AND2 C741 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[36]), .Z(N118)
         );
  GTECH_AND2 C742 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[35]), .Z(N120)
         );
  GTECH_OR2 C743 ( .A(N125), .B(N126), .Z(m2stg_frac1_in[32]) );
  GTECH_OR2 C744 ( .A(N123), .B(N124), .Z(N125) );
  GTECH_OR2 C745 ( .A(N121), .B(N122), .Z(N123) );
  GTECH_AND2 C746 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[32]), .Z(N121)
         );
  GTECH_AND2 C747 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[31]), .Z(N122)
         );
  GTECH_AND2 C748 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[35]), .Z(N124)
         );
  GTECH_AND2 C749 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[34]), .Z(N126)
         );
  GTECH_OR2 C750 ( .A(N131), .B(N132), .Z(m2stg_frac1_in[31]) );
  GTECH_OR2 C751 ( .A(N129), .B(N130), .Z(N131) );
  GTECH_OR2 C752 ( .A(N127), .B(N128), .Z(N129) );
  GTECH_AND2 C753 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[31]), .Z(N127)
         );
  GTECH_AND2 C754 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[30]), .Z(N128)
         );
  GTECH_AND2 C755 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[34]), .Z(N130)
         );
  GTECH_AND2 C756 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[33]), .Z(N132)
         );
  GTECH_OR2 C757 ( .A(N137), .B(N138), .Z(m2stg_frac1_in[30]) );
  GTECH_OR2 C758 ( .A(N135), .B(N136), .Z(N137) );
  GTECH_OR2 C759 ( .A(N133), .B(N134), .Z(N135) );
  GTECH_AND2 C760 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[30]), .Z(N133)
         );
  GTECH_AND2 C761 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[29]), .Z(N134)
         );
  GTECH_AND2 C762 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[33]), .Z(N136)
         );
  GTECH_AND2 C763 ( .A(m2stg_frac1_sng_dnrm), .B(mul_frac_in1[32]), .Z(N138)
         );
  GTECH_OR2 C764 ( .A(N141), .B(N142), .Z(m2stg_frac1_in[29]) );
  GTECH_OR2 C765 ( .A(N139), .B(N140), .Z(N141) );
  GTECH_AND2 C766 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[29]), .Z(N139)
         );
  GTECH_AND2 C767 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[28]), .Z(N140)
         );
  GTECH_AND2 C768 ( .A(m2stg_frac1_sng_norm), .B(mul_frac_in1[32]), .Z(N142)
         );
  GTECH_OR2 C769 ( .A(N143), .B(N144), .Z(m2stg_frac1_in[28]) );
  GTECH_AND2 C770 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[28]), .Z(N143)
         );
  GTECH_AND2 C771 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[27]), .Z(N144)
         );
  GTECH_OR2 C772 ( .A(N145), .B(N146), .Z(m2stg_frac1_in[27]) );
  GTECH_AND2 C773 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[27]), .Z(N145)
         );
  GTECH_AND2 C774 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[26]), .Z(N146)
         );
  GTECH_OR2 C775 ( .A(N147), .B(N148), .Z(m2stg_frac1_in[26]) );
  GTECH_AND2 C776 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[26]), .Z(N147)
         );
  GTECH_AND2 C777 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[25]), .Z(N148)
         );
  GTECH_OR2 C778 ( .A(N149), .B(N150), .Z(m2stg_frac1_in[25]) );
  GTECH_AND2 C779 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[25]), .Z(N149)
         );
  GTECH_AND2 C780 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[24]), .Z(N150)
         );
  GTECH_OR2 C781 ( .A(N151), .B(N152), .Z(m2stg_frac1_in[24]) );
  GTECH_AND2 C782 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[24]), .Z(N151)
         );
  GTECH_AND2 C783 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[23]), .Z(N152)
         );
  GTECH_OR2 C784 ( .A(N153), .B(N154), .Z(m2stg_frac1_in[23]) );
  GTECH_AND2 C785 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[23]), .Z(N153)
         );
  GTECH_AND2 C786 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[22]), .Z(N154)
         );
  GTECH_OR2 C787 ( .A(N155), .B(N156), .Z(m2stg_frac1_in[22]) );
  GTECH_AND2 C788 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[22]), .Z(N155)
         );
  GTECH_AND2 C789 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[21]), .Z(N156)
         );
  GTECH_OR2 C790 ( .A(N157), .B(N158), .Z(m2stg_frac1_in[21]) );
  GTECH_AND2 C791 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[21]), .Z(N157)
         );
  GTECH_AND2 C792 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[20]), .Z(N158)
         );
  GTECH_OR2 C793 ( .A(N159), .B(N160), .Z(m2stg_frac1_in[20]) );
  GTECH_AND2 C794 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[20]), .Z(N159)
         );
  GTECH_AND2 C795 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[19]), .Z(N160)
         );
  GTECH_OR2 C796 ( .A(N161), .B(N162), .Z(m2stg_frac1_in[19]) );
  GTECH_AND2 C797 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[19]), .Z(N161)
         );
  GTECH_AND2 C798 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[18]), .Z(N162)
         );
  GTECH_OR2 C799 ( .A(N163), .B(N164), .Z(m2stg_frac1_in[18]) );
  GTECH_AND2 C800 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[18]), .Z(N163)
         );
  GTECH_AND2 C801 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[17]), .Z(N164)
         );
  GTECH_OR2 C802 ( .A(N165), .B(N166), .Z(m2stg_frac1_in[17]) );
  GTECH_AND2 C803 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[17]), .Z(N165)
         );
  GTECH_AND2 C804 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[16]), .Z(N166)
         );
  GTECH_OR2 C805 ( .A(N167), .B(N168), .Z(m2stg_frac1_in[16]) );
  GTECH_AND2 C806 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[16]), .Z(N167)
         );
  GTECH_AND2 C807 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[15]), .Z(N168)
         );
  GTECH_OR2 C808 ( .A(N169), .B(N170), .Z(m2stg_frac1_in[15]) );
  GTECH_AND2 C809 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[15]), .Z(N169)
         );
  GTECH_AND2 C810 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[14]), .Z(N170)
         );
  GTECH_OR2 C811 ( .A(N171), .B(N172), .Z(m2stg_frac1_in[14]) );
  GTECH_AND2 C812 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[14]), .Z(N171)
         );
  GTECH_AND2 C813 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[13]), .Z(N172)
         );
  GTECH_OR2 C814 ( .A(N173), .B(N174), .Z(m2stg_frac1_in[13]) );
  GTECH_AND2 C815 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[13]), .Z(N173)
         );
  GTECH_AND2 C816 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[12]), .Z(N174)
         );
  GTECH_OR2 C817 ( .A(N175), .B(N176), .Z(m2stg_frac1_in[12]) );
  GTECH_AND2 C818 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[12]), .Z(N175)
         );
  GTECH_AND2 C819 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[11]), .Z(N176)
         );
  GTECH_OR2 C820 ( .A(N177), .B(N178), .Z(m2stg_frac1_in[11]) );
  GTECH_AND2 C821 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[11]), .Z(N177)
         );
  GTECH_AND2 C822 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[10]), .Z(N178)
         );
  GTECH_OR2 C823 ( .A(N179), .B(N180), .Z(m2stg_frac1_in[10]) );
  GTECH_AND2 C824 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[10]), .Z(N179)
         );
  GTECH_AND2 C825 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[9]), .Z(N180) );
  GTECH_OR2 C826 ( .A(N181), .B(N182), .Z(m2stg_frac1_in[9]) );
  GTECH_AND2 C827 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[9]), .Z(N181) );
  GTECH_AND2 C828 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[8]), .Z(N182) );
  GTECH_OR2 C829 ( .A(N183), .B(N184), .Z(m2stg_frac1_in[8]) );
  GTECH_AND2 C830 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[8]), .Z(N183) );
  GTECH_AND2 C831 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[7]), .Z(N184) );
  GTECH_OR2 C832 ( .A(N185), .B(N186), .Z(m2stg_frac1_in[7]) );
  GTECH_AND2 C833 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[7]), .Z(N185) );
  GTECH_AND2 C834 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[6]), .Z(N186) );
  GTECH_OR2 C835 ( .A(N187), .B(N188), .Z(m2stg_frac1_in[6]) );
  GTECH_AND2 C836 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[6]), .Z(N187) );
  GTECH_AND2 C837 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[5]), .Z(N188) );
  GTECH_OR2 C838 ( .A(N189), .B(N190), .Z(m2stg_frac1_in[5]) );
  GTECH_AND2 C839 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[5]), .Z(N189) );
  GTECH_AND2 C840 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[4]), .Z(N190) );
  GTECH_OR2 C841 ( .A(N191), .B(N192), .Z(m2stg_frac1_in[4]) );
  GTECH_AND2 C842 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[4]), .Z(N191) );
  GTECH_AND2 C843 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[3]), .Z(N192) );
  GTECH_OR2 C844 ( .A(N193), .B(N194), .Z(m2stg_frac1_in[3]) );
  GTECH_AND2 C845 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[3]), .Z(N193) );
  GTECH_AND2 C846 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[2]), .Z(N194) );
  GTECH_OR2 C847 ( .A(N195), .B(N196), .Z(m2stg_frac1_in[2]) );
  GTECH_AND2 C848 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[2]), .Z(N195) );
  GTECH_AND2 C849 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[1]), .Z(N196) );
  GTECH_OR2 C850 ( .A(N197), .B(N198), .Z(m2stg_frac1_in[1]) );
  GTECH_AND2 C851 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[1]), .Z(N197) );
  GTECH_AND2 C852 ( .A(m2stg_frac1_dbl_dnrm), .B(mul_frac_in1[0]), .Z(N198) );
  GTECH_AND2 C853 ( .A(m2stg_frac1_dbl_norm), .B(mul_frac_in1[0]), .Z(
        m2stg_frac1_in[0]) );
  GTECH_NOT I_1 ( .A(m2stg_frac1_in[52]), .Z(m2stg_frac1_array_in[52]) );
  GTECH_NOT I_2 ( .A(m2stg_frac1_in[51]), .Z(m2stg_frac1_array_in[51]) );
  GTECH_NOT I_3 ( .A(m2stg_frac1_in[50]), .Z(m2stg_frac1_array_in[50]) );
  GTECH_NOT I_4 ( .A(m2stg_frac1_in[49]), .Z(m2stg_frac1_array_in[49]) );
  GTECH_NOT I_5 ( .A(m2stg_frac1_in[48]), .Z(m2stg_frac1_array_in[48]) );
  GTECH_NOT I_6 ( .A(m2stg_frac1_in[47]), .Z(m2stg_frac1_array_in[47]) );
  GTECH_NOT I_7 ( .A(m2stg_frac1_in[46]), .Z(m2stg_frac1_array_in[46]) );
  GTECH_NOT I_8 ( .A(m2stg_frac1_in[45]), .Z(m2stg_frac1_array_in[45]) );
  GTECH_NOT I_9 ( .A(m2stg_frac1_in[44]), .Z(m2stg_frac1_array_in[44]) );
  GTECH_NOT I_10 ( .A(m2stg_frac1_in[43]), .Z(m2stg_frac1_array_in[43]) );
  GTECH_NOT I_11 ( .A(m2stg_frac1_in[42]), .Z(m2stg_frac1_array_in[42]) );
  GTECH_NOT I_12 ( .A(m2stg_frac1_in[41]), .Z(m2stg_frac1_array_in[41]) );
  GTECH_NOT I_13 ( .A(m2stg_frac1_in[40]), .Z(m2stg_frac1_array_in[40]) );
  GTECH_NOT I_14 ( .A(m2stg_frac1_in[39]), .Z(m2stg_frac1_array_in[39]) );
  GTECH_NOT I_15 ( .A(m2stg_frac1_in[38]), .Z(m2stg_frac1_array_in[38]) );
  GTECH_NOT I_16 ( .A(m2stg_frac1_in[37]), .Z(m2stg_frac1_array_in[37]) );
  GTECH_NOT I_17 ( .A(m2stg_frac1_in[36]), .Z(m2stg_frac1_array_in[36]) );
  GTECH_NOT I_18 ( .A(m2stg_frac1_in[35]), .Z(m2stg_frac1_array_in[35]) );
  GTECH_NOT I_19 ( .A(m2stg_frac1_in[34]), .Z(m2stg_frac1_array_in[34]) );
  GTECH_NOT I_20 ( .A(m2stg_frac1_in[33]), .Z(m2stg_frac1_array_in[33]) );
  GTECH_NOT I_21 ( .A(m2stg_frac1_in[32]), .Z(m2stg_frac1_array_in[32]) );
  GTECH_NOT I_22 ( .A(m2stg_frac1_in[31]), .Z(m2stg_frac1_array_in[31]) );
  GTECH_NOT I_23 ( .A(m2stg_frac1_in[30]), .Z(m2stg_frac1_array_in[30]) );
  GTECH_NOT I_24 ( .A(m2stg_frac1_in[29]), .Z(m2stg_frac1_array_in[29]) );
  GTECH_NOT I_25 ( .A(m2stg_frac1_in[28]), .Z(m2stg_frac1_array_in[28]) );
  GTECH_NOT I_26 ( .A(m2stg_frac1_in[27]), .Z(m2stg_frac1_array_in[27]) );
  GTECH_NOT I_27 ( .A(m2stg_frac1_in[26]), .Z(m2stg_frac1_array_in[26]) );
  GTECH_NOT I_28 ( .A(m2stg_frac1_in[25]), .Z(m2stg_frac1_array_in[25]) );
  GTECH_NOT I_29 ( .A(m2stg_frac1_in[24]), .Z(m2stg_frac1_array_in[24]) );
  GTECH_NOT I_30 ( .A(m2stg_frac1_in[23]), .Z(m2stg_frac1_array_in[23]) );
  GTECH_NOT I_31 ( .A(m2stg_frac1_in[22]), .Z(m2stg_frac1_array_in[22]) );
  GTECH_NOT I_32 ( .A(m2stg_frac1_in[21]), .Z(m2stg_frac1_array_in[21]) );
  GTECH_NOT I_33 ( .A(m2stg_frac1_in[20]), .Z(m2stg_frac1_array_in[20]) );
  GTECH_NOT I_34 ( .A(m2stg_frac1_in[19]), .Z(m2stg_frac1_array_in[19]) );
  GTECH_NOT I_35 ( .A(m2stg_frac1_in[18]), .Z(m2stg_frac1_array_in[18]) );
  GTECH_NOT I_36 ( .A(m2stg_frac1_in[17]), .Z(m2stg_frac1_array_in[17]) );
  GTECH_NOT I_37 ( .A(m2stg_frac1_in[16]), .Z(m2stg_frac1_array_in[16]) );
  GTECH_NOT I_38 ( .A(m2stg_frac1_in[15]), .Z(m2stg_frac1_array_in[15]) );
  GTECH_NOT I_39 ( .A(m2stg_frac1_in[14]), .Z(m2stg_frac1_array_in[14]) );
  GTECH_NOT I_40 ( .A(m2stg_frac1_in[13]), .Z(m2stg_frac1_array_in[13]) );
  GTECH_NOT I_41 ( .A(m2stg_frac1_in[12]), .Z(m2stg_frac1_array_in[12]) );
  GTECH_NOT I_42 ( .A(m2stg_frac1_in[11]), .Z(m2stg_frac1_array_in[11]) );
  GTECH_NOT I_43 ( .A(m2stg_frac1_in[10]), .Z(m2stg_frac1_array_in[10]) );
  GTECH_NOT I_44 ( .A(m2stg_frac1_in[9]), .Z(m2stg_frac1_array_in[9]) );
  GTECH_NOT I_45 ( .A(m2stg_frac1_in[8]), .Z(m2stg_frac1_array_in[8]) );
  GTECH_NOT I_46 ( .A(m2stg_frac1_in[7]), .Z(m2stg_frac1_array_in[7]) );
  GTECH_NOT I_47 ( .A(m2stg_frac1_in[6]), .Z(m2stg_frac1_array_in[6]) );
  GTECH_NOT I_48 ( .A(m2stg_frac1_in[5]), .Z(m2stg_frac1_array_in[5]) );
  GTECH_NOT I_49 ( .A(m2stg_frac1_in[4]), .Z(m2stg_frac1_array_in[4]) );
  GTECH_NOT I_50 ( .A(m2stg_frac1_in[3]), .Z(m2stg_frac1_array_in[3]) );
  GTECH_NOT I_51 ( .A(m2stg_frac1_in[2]), .Z(m2stg_frac1_array_in[2]) );
  GTECH_NOT I_52 ( .A(m2stg_frac1_in[1]), .Z(m2stg_frac1_array_in[1]) );
  GTECH_NOT I_53 ( .A(m2stg_frac1_in[0]), .Z(m2stg_frac1_array_in[0]) );
  GTECH_OR2 C907 ( .A(N203), .B(m2stg_frac2_inf), .Z(m2stg_frac2_array_in[52])
         );
  GTECH_OR2 C908 ( .A(N201), .B(N202), .Z(N203) );
  GTECH_OR2 C909 ( .A(N200), .B(m2stg_frac2_sng_norm), .Z(N201) );
  GTECH_OR2 C910 ( .A(m2stg_frac2_dbl_norm), .B(N199), .Z(N200) );
  GTECH_AND2 C911 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[51]), .Z(N199)
         );
  GTECH_AND2 C912 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[54]), .Z(N202)
         );
  GTECH_OR2 C913 ( .A(N212), .B(N213), .Z(m2stg_frac2_array_in[51]) );
  GTECH_OR2 C914 ( .A(N210), .B(N211), .Z(N212) );
  GTECH_OR2 C915 ( .A(N207), .B(N209), .Z(N210) );
  GTECH_OR2 C916 ( .A(N205), .B(N206), .Z(N207) );
  GTECH_AND2 C917 ( .A(m2stg_frac2_dbl_norm), .B(N204), .Z(N205) );
  GTECH_OR2 C918 ( .A(mul_frac_in2[51]), .B(m1stg_snan_dbl_in2), .Z(N204) );
  GTECH_AND2 C919 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[50]), .Z(N206)
         );
  GTECH_AND2 C920 ( .A(m2stg_frac2_sng_norm), .B(N208), .Z(N209) );
  GTECH_OR2 C921 ( .A(mul_frac_in2[54]), .B(m1stg_snan_sng_in2), .Z(N208) );
  GTECH_AND2 C922 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[53]), .Z(N211)
         );
  GTECH_AND2 C923 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N213) );
  GTECH_OR2 C924 ( .A(N220), .B(N221), .Z(m2stg_frac2_array_in[50]) );
  GTECH_OR2 C925 ( .A(N218), .B(N219), .Z(N220) );
  GTECH_OR2 C926 ( .A(N216), .B(N217), .Z(N218) );
  GTECH_OR2 C927 ( .A(N214), .B(N215), .Z(N216) );
  GTECH_AND2 C928 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[50]), .Z(N214)
         );
  GTECH_AND2 C929 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[49]), .Z(N215)
         );
  GTECH_AND2 C930 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[53]), .Z(N217)
         );
  GTECH_AND2 C931 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[52]), .Z(N219)
         );
  GTECH_AND2 C932 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N221) );
  GTECH_OR2 C933 ( .A(N228), .B(N229), .Z(m2stg_frac2_array_in[49]) );
  GTECH_OR2 C934 ( .A(N226), .B(N227), .Z(N228) );
  GTECH_OR2 C935 ( .A(N224), .B(N225), .Z(N226) );
  GTECH_OR2 C936 ( .A(N222), .B(N223), .Z(N224) );
  GTECH_AND2 C937 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[49]), .Z(N222)
         );
  GTECH_AND2 C938 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[48]), .Z(N223)
         );
  GTECH_AND2 C939 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[52]), .Z(N225)
         );
  GTECH_AND2 C940 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[51]), .Z(N227)
         );
  GTECH_AND2 C941 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N229) );
  GTECH_OR2 C942 ( .A(N236), .B(N237), .Z(m2stg_frac2_array_in[48]) );
  GTECH_OR2 C943 ( .A(N234), .B(N235), .Z(N236) );
  GTECH_OR2 C944 ( .A(N232), .B(N233), .Z(N234) );
  GTECH_OR2 C945 ( .A(N230), .B(N231), .Z(N232) );
  GTECH_AND2 C946 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[48]), .Z(N230)
         );
  GTECH_AND2 C947 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[47]), .Z(N231)
         );
  GTECH_AND2 C948 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[51]), .Z(N233)
         );
  GTECH_AND2 C949 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[50]), .Z(N235)
         );
  GTECH_AND2 C950 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N237) );
  GTECH_OR2 C951 ( .A(N244), .B(N245), .Z(m2stg_frac2_array_in[47]) );
  GTECH_OR2 C952 ( .A(N242), .B(N243), .Z(N244) );
  GTECH_OR2 C953 ( .A(N240), .B(N241), .Z(N242) );
  GTECH_OR2 C954 ( .A(N238), .B(N239), .Z(N240) );
  GTECH_AND2 C955 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[47]), .Z(N238)
         );
  GTECH_AND2 C956 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[46]), .Z(N239)
         );
  GTECH_AND2 C957 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[50]), .Z(N241)
         );
  GTECH_AND2 C958 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[49]), .Z(N243)
         );
  GTECH_AND2 C959 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N245) );
  GTECH_OR2 C960 ( .A(N252), .B(N253), .Z(m2stg_frac2_array_in[46]) );
  GTECH_OR2 C961 ( .A(N250), .B(N251), .Z(N252) );
  GTECH_OR2 C962 ( .A(N248), .B(N249), .Z(N250) );
  GTECH_OR2 C963 ( .A(N246), .B(N247), .Z(N248) );
  GTECH_AND2 C964 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[46]), .Z(N246)
         );
  GTECH_AND2 C965 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[45]), .Z(N247)
         );
  GTECH_AND2 C966 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[49]), .Z(N249)
         );
  GTECH_AND2 C967 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[48]), .Z(N251)
         );
  GTECH_AND2 C968 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N253) );
  GTECH_OR2 C969 ( .A(N260), .B(N261), .Z(m2stg_frac2_array_in[45]) );
  GTECH_OR2 C970 ( .A(N258), .B(N259), .Z(N260) );
  GTECH_OR2 C971 ( .A(N256), .B(N257), .Z(N258) );
  GTECH_OR2 C972 ( .A(N254), .B(N255), .Z(N256) );
  GTECH_AND2 C973 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[45]), .Z(N254)
         );
  GTECH_AND2 C974 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[44]), .Z(N255)
         );
  GTECH_AND2 C975 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[48]), .Z(N257)
         );
  GTECH_AND2 C976 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[47]), .Z(N259)
         );
  GTECH_AND2 C977 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N261) );
  GTECH_OR2 C978 ( .A(N268), .B(N269), .Z(m2stg_frac2_array_in[44]) );
  GTECH_OR2 C979 ( .A(N266), .B(N267), .Z(N268) );
  GTECH_OR2 C980 ( .A(N264), .B(N265), .Z(N266) );
  GTECH_OR2 C981 ( .A(N262), .B(N263), .Z(N264) );
  GTECH_AND2 C982 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[44]), .Z(N262)
         );
  GTECH_AND2 C983 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[43]), .Z(N263)
         );
  GTECH_AND2 C984 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[47]), .Z(N265)
         );
  GTECH_AND2 C985 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[46]), .Z(N267)
         );
  GTECH_AND2 C986 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N269) );
  GTECH_OR2 C987 ( .A(N276), .B(N277), .Z(m2stg_frac2_array_in[43]) );
  GTECH_OR2 C988 ( .A(N274), .B(N275), .Z(N276) );
  GTECH_OR2 C989 ( .A(N272), .B(N273), .Z(N274) );
  GTECH_OR2 C990 ( .A(N270), .B(N271), .Z(N272) );
  GTECH_AND2 C991 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[43]), .Z(N270)
         );
  GTECH_AND2 C992 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[42]), .Z(N271)
         );
  GTECH_AND2 C993 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[46]), .Z(N273)
         );
  GTECH_AND2 C994 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[45]), .Z(N275)
         );
  GTECH_AND2 C995 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N277) );
  GTECH_OR2 C996 ( .A(N284), .B(N285), .Z(m2stg_frac2_array_in[42]) );
  GTECH_OR2 C997 ( .A(N282), .B(N283), .Z(N284) );
  GTECH_OR2 C998 ( .A(N280), .B(N281), .Z(N282) );
  GTECH_OR2 C999 ( .A(N278), .B(N279), .Z(N280) );
  GTECH_AND2 C1000 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[42]), .Z(N278)
         );
  GTECH_AND2 C1001 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[41]), .Z(N279)
         );
  GTECH_AND2 C1002 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[45]), .Z(N281)
         );
  GTECH_AND2 C1003 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[44]), .Z(N283)
         );
  GTECH_AND2 C1004 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N285) );
  GTECH_OR2 C1005 ( .A(N292), .B(N293), .Z(m2stg_frac2_array_in[41]) );
  GTECH_OR2 C1006 ( .A(N290), .B(N291), .Z(N292) );
  GTECH_OR2 C1007 ( .A(N288), .B(N289), .Z(N290) );
  GTECH_OR2 C1008 ( .A(N286), .B(N287), .Z(N288) );
  GTECH_AND2 C1009 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[41]), .Z(N286)
         );
  GTECH_AND2 C1010 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[40]), .Z(N287)
         );
  GTECH_AND2 C1011 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[44]), .Z(N289)
         );
  GTECH_AND2 C1012 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[43]), .Z(N291)
         );
  GTECH_AND2 C1013 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N293) );
  GTECH_OR2 C1014 ( .A(N300), .B(N301), .Z(m2stg_frac2_array_in[40]) );
  GTECH_OR2 C1015 ( .A(N298), .B(N299), .Z(N300) );
  GTECH_OR2 C1016 ( .A(N296), .B(N297), .Z(N298) );
  GTECH_OR2 C1017 ( .A(N294), .B(N295), .Z(N296) );
  GTECH_AND2 C1018 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[40]), .Z(N294)
         );
  GTECH_AND2 C1019 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[39]), .Z(N295)
         );
  GTECH_AND2 C1020 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[43]), .Z(N297)
         );
  GTECH_AND2 C1021 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[42]), .Z(N299)
         );
  GTECH_AND2 C1022 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N301) );
  GTECH_OR2 C1023 ( .A(N308), .B(N309), .Z(m2stg_frac2_array_in[39]) );
  GTECH_OR2 C1024 ( .A(N306), .B(N307), .Z(N308) );
  GTECH_OR2 C1025 ( .A(N304), .B(N305), .Z(N306) );
  GTECH_OR2 C1026 ( .A(N302), .B(N303), .Z(N304) );
  GTECH_AND2 C1027 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[39]), .Z(N302)
         );
  GTECH_AND2 C1028 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[38]), .Z(N303)
         );
  GTECH_AND2 C1029 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[42]), .Z(N305)
         );
  GTECH_AND2 C1030 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[41]), .Z(N307)
         );
  GTECH_AND2 C1031 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N309) );
  GTECH_OR2 C1032 ( .A(N316), .B(N317), .Z(m2stg_frac2_array_in[38]) );
  GTECH_OR2 C1033 ( .A(N314), .B(N315), .Z(N316) );
  GTECH_OR2 C1034 ( .A(N312), .B(N313), .Z(N314) );
  GTECH_OR2 C1035 ( .A(N310), .B(N311), .Z(N312) );
  GTECH_AND2 C1036 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[38]), .Z(N310)
         );
  GTECH_AND2 C1037 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[37]), .Z(N311)
         );
  GTECH_AND2 C1038 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[41]), .Z(N313)
         );
  GTECH_AND2 C1039 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[40]), .Z(N315)
         );
  GTECH_AND2 C1040 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N317) );
  GTECH_OR2 C1041 ( .A(N324), .B(N325), .Z(m2stg_frac2_array_in[37]) );
  GTECH_OR2 C1042 ( .A(N322), .B(N323), .Z(N324) );
  GTECH_OR2 C1043 ( .A(N320), .B(N321), .Z(N322) );
  GTECH_OR2 C1044 ( .A(N318), .B(N319), .Z(N320) );
  GTECH_AND2 C1045 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[37]), .Z(N318)
         );
  GTECH_AND2 C1046 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[36]), .Z(N319)
         );
  GTECH_AND2 C1047 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[40]), .Z(N321)
         );
  GTECH_AND2 C1048 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[39]), .Z(N323)
         );
  GTECH_AND2 C1049 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N325) );
  GTECH_OR2 C1050 ( .A(N332), .B(N333), .Z(m2stg_frac2_array_in[36]) );
  GTECH_OR2 C1051 ( .A(N330), .B(N331), .Z(N332) );
  GTECH_OR2 C1052 ( .A(N328), .B(N329), .Z(N330) );
  GTECH_OR2 C1053 ( .A(N326), .B(N327), .Z(N328) );
  GTECH_AND2 C1054 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[36]), .Z(N326)
         );
  GTECH_AND2 C1055 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[35]), .Z(N327)
         );
  GTECH_AND2 C1056 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[39]), .Z(N329)
         );
  GTECH_AND2 C1057 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[38]), .Z(N331)
         );
  GTECH_AND2 C1058 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N333) );
  GTECH_OR2 C1059 ( .A(N340), .B(N341), .Z(m2stg_frac2_array_in[35]) );
  GTECH_OR2 C1060 ( .A(N338), .B(N339), .Z(N340) );
  GTECH_OR2 C1061 ( .A(N336), .B(N337), .Z(N338) );
  GTECH_OR2 C1062 ( .A(N334), .B(N335), .Z(N336) );
  GTECH_AND2 C1063 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[35]), .Z(N334)
         );
  GTECH_AND2 C1064 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[34]), .Z(N335)
         );
  GTECH_AND2 C1065 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[38]), .Z(N337)
         );
  GTECH_AND2 C1066 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[37]), .Z(N339)
         );
  GTECH_AND2 C1067 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N341) );
  GTECH_OR2 C1068 ( .A(N348), .B(N349), .Z(m2stg_frac2_array_in[34]) );
  GTECH_OR2 C1069 ( .A(N346), .B(N347), .Z(N348) );
  GTECH_OR2 C1070 ( .A(N344), .B(N345), .Z(N346) );
  GTECH_OR2 C1071 ( .A(N342), .B(N343), .Z(N344) );
  GTECH_AND2 C1072 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[34]), .Z(N342)
         );
  GTECH_AND2 C1073 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[33]), .Z(N343)
         );
  GTECH_AND2 C1074 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[37]), .Z(N345)
         );
  GTECH_AND2 C1075 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[36]), .Z(N347)
         );
  GTECH_AND2 C1076 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N349) );
  GTECH_OR2 C1077 ( .A(N356), .B(N357), .Z(m2stg_frac2_array_in[33]) );
  GTECH_OR2 C1078 ( .A(N354), .B(N355), .Z(N356) );
  GTECH_OR2 C1079 ( .A(N352), .B(N353), .Z(N354) );
  GTECH_OR2 C1080 ( .A(N350), .B(N351), .Z(N352) );
  GTECH_AND2 C1081 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[33]), .Z(N350)
         );
  GTECH_AND2 C1082 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[32]), .Z(N351)
         );
  GTECH_AND2 C1083 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[36]), .Z(N353)
         );
  GTECH_AND2 C1084 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[35]), .Z(N355)
         );
  GTECH_AND2 C1085 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N357) );
  GTECH_OR2 C1086 ( .A(N364), .B(N365), .Z(m2stg_frac2_array_in[32]) );
  GTECH_OR2 C1087 ( .A(N362), .B(N363), .Z(N364) );
  GTECH_OR2 C1088 ( .A(N360), .B(N361), .Z(N362) );
  GTECH_OR2 C1089 ( .A(N358), .B(N359), .Z(N360) );
  GTECH_AND2 C1090 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[32]), .Z(N358)
         );
  GTECH_AND2 C1091 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[31]), .Z(N359)
         );
  GTECH_AND2 C1092 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[35]), .Z(N361)
         );
  GTECH_AND2 C1093 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[34]), .Z(N363)
         );
  GTECH_AND2 C1094 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N365) );
  GTECH_OR2 C1095 ( .A(N372), .B(N373), .Z(m2stg_frac2_array_in[31]) );
  GTECH_OR2 C1096 ( .A(N370), .B(N371), .Z(N372) );
  GTECH_OR2 C1097 ( .A(N368), .B(N369), .Z(N370) );
  GTECH_OR2 C1098 ( .A(N366), .B(N367), .Z(N368) );
  GTECH_AND2 C1099 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[31]), .Z(N366)
         );
  GTECH_AND2 C1100 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[30]), .Z(N367)
         );
  GTECH_AND2 C1101 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[34]), .Z(N369)
         );
  GTECH_AND2 C1102 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[33]), .Z(N371)
         );
  GTECH_AND2 C1103 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N373) );
  GTECH_OR2 C1104 ( .A(N380), .B(N381), .Z(m2stg_frac2_array_in[30]) );
  GTECH_OR2 C1105 ( .A(N378), .B(N379), .Z(N380) );
  GTECH_OR2 C1106 ( .A(N376), .B(N377), .Z(N378) );
  GTECH_OR2 C1107 ( .A(N374), .B(N375), .Z(N376) );
  GTECH_AND2 C1108 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[30]), .Z(N374)
         );
  GTECH_AND2 C1109 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[29]), .Z(N375)
         );
  GTECH_AND2 C1110 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[33]), .Z(N377)
         );
  GTECH_AND2 C1111 ( .A(m2stg_frac2_sng_dnrm), .B(mul_frac_in2[32]), .Z(N379)
         );
  GTECH_AND2 C1112 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N381) );
  GTECH_OR2 C1113 ( .A(N386), .B(N387), .Z(m2stg_frac2_array_in[29]) );
  GTECH_OR2 C1114 ( .A(N384), .B(N385), .Z(N386) );
  GTECH_OR2 C1115 ( .A(N382), .B(N383), .Z(N384) );
  GTECH_AND2 C1116 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[29]), .Z(N382)
         );
  GTECH_AND2 C1117 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[28]), .Z(N383)
         );
  GTECH_AND2 C1118 ( .A(m2stg_frac2_sng_norm), .B(mul_frac_in2[32]), .Z(N385)
         );
  GTECH_AND2 C1119 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in), .Z(N387) );
  GTECH_OR2 C1120 ( .A(N390), .B(N391), .Z(m2stg_frac2_array_in[28]) );
  GTECH_OR2 C1121 ( .A(N388), .B(N389), .Z(N390) );
  GTECH_AND2 C1122 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[28]), .Z(N388)
         );
  GTECH_AND2 C1123 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[27]), .Z(N389)
         );
  GTECH_AND2 C1124 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N391)
         );
  GTECH_OR2 C1125 ( .A(N394), .B(N395), .Z(m2stg_frac2_array_in[27]) );
  GTECH_OR2 C1126 ( .A(N392), .B(N393), .Z(N394) );
  GTECH_AND2 C1127 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[27]), .Z(N392)
         );
  GTECH_AND2 C1128 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[26]), .Z(N393)
         );
  GTECH_AND2 C1129 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N395)
         );
  GTECH_OR2 C1130 ( .A(N398), .B(N399), .Z(m2stg_frac2_array_in[26]) );
  GTECH_OR2 C1131 ( .A(N396), .B(N397), .Z(N398) );
  GTECH_AND2 C1132 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[26]), .Z(N396)
         );
  GTECH_AND2 C1133 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[25]), .Z(N397)
         );
  GTECH_AND2 C1134 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N399)
         );
  GTECH_OR2 C1135 ( .A(N402), .B(N403), .Z(m2stg_frac2_array_in[25]) );
  GTECH_OR2 C1136 ( .A(N400), .B(N401), .Z(N402) );
  GTECH_AND2 C1137 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[25]), .Z(N400)
         );
  GTECH_AND2 C1138 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[24]), .Z(N401)
         );
  GTECH_AND2 C1139 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N403)
         );
  GTECH_OR2 C1140 ( .A(N406), .B(N407), .Z(m2stg_frac2_array_in[24]) );
  GTECH_OR2 C1141 ( .A(N404), .B(N405), .Z(N406) );
  GTECH_AND2 C1142 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[24]), .Z(N404)
         );
  GTECH_AND2 C1143 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[23]), .Z(N405)
         );
  GTECH_AND2 C1144 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N407)
         );
  GTECH_OR2 C1145 ( .A(N410), .B(N411), .Z(m2stg_frac2_array_in[23]) );
  GTECH_OR2 C1146 ( .A(N408), .B(N409), .Z(N410) );
  GTECH_AND2 C1147 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[23]), .Z(N408)
         );
  GTECH_AND2 C1148 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[22]), .Z(N409)
         );
  GTECH_AND2 C1149 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N411)
         );
  GTECH_OR2 C1150 ( .A(N414), .B(N415), .Z(m2stg_frac2_array_in[22]) );
  GTECH_OR2 C1151 ( .A(N412), .B(N413), .Z(N414) );
  GTECH_AND2 C1152 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[22]), .Z(N412)
         );
  GTECH_AND2 C1153 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[21]), .Z(N413)
         );
  GTECH_AND2 C1154 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N415)
         );
  GTECH_OR2 C1155 ( .A(N418), .B(N419), .Z(m2stg_frac2_array_in[21]) );
  GTECH_OR2 C1156 ( .A(N416), .B(N417), .Z(N418) );
  GTECH_AND2 C1157 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[21]), .Z(N416)
         );
  GTECH_AND2 C1158 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[20]), .Z(N417)
         );
  GTECH_AND2 C1159 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N419)
         );
  GTECH_OR2 C1160 ( .A(N422), .B(N423), .Z(m2stg_frac2_array_in[20]) );
  GTECH_OR2 C1161 ( .A(N420), .B(N421), .Z(N422) );
  GTECH_AND2 C1162 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[20]), .Z(N420)
         );
  GTECH_AND2 C1163 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[19]), .Z(N421)
         );
  GTECH_AND2 C1164 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N423)
         );
  GTECH_OR2 C1165 ( .A(N426), .B(N427), .Z(m2stg_frac2_array_in[19]) );
  GTECH_OR2 C1166 ( .A(N424), .B(N425), .Z(N426) );
  GTECH_AND2 C1167 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[19]), .Z(N424)
         );
  GTECH_AND2 C1168 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[18]), .Z(N425)
         );
  GTECH_AND2 C1169 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N427)
         );
  GTECH_OR2 C1170 ( .A(N430), .B(N431), .Z(m2stg_frac2_array_in[18]) );
  GTECH_OR2 C1171 ( .A(N428), .B(N429), .Z(N430) );
  GTECH_AND2 C1172 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[18]), .Z(N428)
         );
  GTECH_AND2 C1173 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[17]), .Z(N429)
         );
  GTECH_AND2 C1174 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N431)
         );
  GTECH_OR2 C1175 ( .A(N434), .B(N435), .Z(m2stg_frac2_array_in[17]) );
  GTECH_OR2 C1176 ( .A(N432), .B(N433), .Z(N434) );
  GTECH_AND2 C1177 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[17]), .Z(N432)
         );
  GTECH_AND2 C1178 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[16]), .Z(N433)
         );
  GTECH_AND2 C1179 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N435)
         );
  GTECH_OR2 C1180 ( .A(N438), .B(N439), .Z(m2stg_frac2_array_in[16]) );
  GTECH_OR2 C1181 ( .A(N436), .B(N437), .Z(N438) );
  GTECH_AND2 C1182 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[16]), .Z(N436)
         );
  GTECH_AND2 C1183 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[15]), .Z(N437)
         );
  GTECH_AND2 C1184 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N439)
         );
  GTECH_OR2 C1185 ( .A(N442), .B(N443), .Z(m2stg_frac2_array_in[15]) );
  GTECH_OR2 C1186 ( .A(N440), .B(N441), .Z(N442) );
  GTECH_AND2 C1187 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[15]), .Z(N440)
         );
  GTECH_AND2 C1188 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[14]), .Z(N441)
         );
  GTECH_AND2 C1189 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N443)
         );
  GTECH_OR2 C1190 ( .A(N446), .B(N447), .Z(m2stg_frac2_array_in[14]) );
  GTECH_OR2 C1191 ( .A(N444), .B(N445), .Z(N446) );
  GTECH_AND2 C1192 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[14]), .Z(N444)
         );
  GTECH_AND2 C1193 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[13]), .Z(N445)
         );
  GTECH_AND2 C1194 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N447)
         );
  GTECH_OR2 C1195 ( .A(N450), .B(N451), .Z(m2stg_frac2_array_in[13]) );
  GTECH_OR2 C1196 ( .A(N448), .B(N449), .Z(N450) );
  GTECH_AND2 C1197 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[13]), .Z(N448)
         );
  GTECH_AND2 C1198 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[12]), .Z(N449)
         );
  GTECH_AND2 C1199 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N451)
         );
  GTECH_OR2 C1200 ( .A(N454), .B(N455), .Z(m2stg_frac2_array_in[12]) );
  GTECH_OR2 C1201 ( .A(N452), .B(N453), .Z(N454) );
  GTECH_AND2 C1202 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[12]), .Z(N452)
         );
  GTECH_AND2 C1203 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[11]), .Z(N453)
         );
  GTECH_AND2 C1204 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N455)
         );
  GTECH_OR2 C1205 ( .A(N458), .B(N459), .Z(m2stg_frac2_array_in[11]) );
  GTECH_OR2 C1206 ( .A(N456), .B(N457), .Z(N458) );
  GTECH_AND2 C1207 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[11]), .Z(N456)
         );
  GTECH_AND2 C1208 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[10]), .Z(N457)
         );
  GTECH_AND2 C1209 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N459)
         );
  GTECH_OR2 C1210 ( .A(N462), .B(N463), .Z(m2stg_frac2_array_in[10]) );
  GTECH_OR2 C1211 ( .A(N460), .B(N461), .Z(N462) );
  GTECH_AND2 C1212 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[10]), .Z(N460)
         );
  GTECH_AND2 C1213 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[9]), .Z(N461)
         );
  GTECH_AND2 C1214 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N463)
         );
  GTECH_OR2 C1215 ( .A(N466), .B(N467), .Z(m2stg_frac2_array_in[9]) );
  GTECH_OR2 C1216 ( .A(N464), .B(N465), .Z(N466) );
  GTECH_AND2 C1217 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[9]), .Z(N464)
         );
  GTECH_AND2 C1218 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[8]), .Z(N465)
         );
  GTECH_AND2 C1219 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N467)
         );
  GTECH_OR2 C1220 ( .A(N470), .B(N471), .Z(m2stg_frac2_array_in[8]) );
  GTECH_OR2 C1221 ( .A(N468), .B(N469), .Z(N470) );
  GTECH_AND2 C1222 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[8]), .Z(N468)
         );
  GTECH_AND2 C1223 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[7]), .Z(N469)
         );
  GTECH_AND2 C1224 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N471)
         );
  GTECH_OR2 C1225 ( .A(N474), .B(N475), .Z(m2stg_frac2_array_in[7]) );
  GTECH_OR2 C1226 ( .A(N472), .B(N473), .Z(N474) );
  GTECH_AND2 C1227 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[7]), .Z(N472)
         );
  GTECH_AND2 C1228 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[6]), .Z(N473)
         );
  GTECH_AND2 C1229 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N475)
         );
  GTECH_OR2 C1230 ( .A(N478), .B(N479), .Z(m2stg_frac2_array_in[6]) );
  GTECH_OR2 C1231 ( .A(N476), .B(N477), .Z(N478) );
  GTECH_AND2 C1232 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[6]), .Z(N476)
         );
  GTECH_AND2 C1233 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[5]), .Z(N477)
         );
  GTECH_AND2 C1234 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N479)
         );
  GTECH_OR2 C1235 ( .A(N482), .B(N483), .Z(m2stg_frac2_array_in[5]) );
  GTECH_OR2 C1236 ( .A(N480), .B(N481), .Z(N482) );
  GTECH_AND2 C1237 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[5]), .Z(N480)
         );
  GTECH_AND2 C1238 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[4]), .Z(N481)
         );
  GTECH_AND2 C1239 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N483)
         );
  GTECH_OR2 C1240 ( .A(N486), .B(N487), .Z(m2stg_frac2_array_in[4]) );
  GTECH_OR2 C1241 ( .A(N484), .B(N485), .Z(N486) );
  GTECH_AND2 C1242 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[4]), .Z(N484)
         );
  GTECH_AND2 C1243 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[3]), .Z(N485)
         );
  GTECH_AND2 C1244 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N487)
         );
  GTECH_OR2 C1245 ( .A(N490), .B(N491), .Z(m2stg_frac2_array_in[3]) );
  GTECH_OR2 C1246 ( .A(N488), .B(N489), .Z(N490) );
  GTECH_AND2 C1247 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[3]), .Z(N488)
         );
  GTECH_AND2 C1248 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[2]), .Z(N489)
         );
  GTECH_AND2 C1249 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N491)
         );
  GTECH_OR2 C1250 ( .A(N494), .B(N495), .Z(m2stg_frac2_array_in[2]) );
  GTECH_OR2 C1251 ( .A(N492), .B(N493), .Z(N494) );
  GTECH_AND2 C1252 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[2]), .Z(N492)
         );
  GTECH_AND2 C1253 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[1]), .Z(N493)
         );
  GTECH_AND2 C1254 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N495)
         );
  GTECH_OR2 C1255 ( .A(N498), .B(N499), .Z(m2stg_frac2_array_in[1]) );
  GTECH_OR2 C1256 ( .A(N496), .B(N497), .Z(N498) );
  GTECH_AND2 C1257 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[1]), .Z(N496)
         );
  GTECH_AND2 C1258 ( .A(m2stg_frac2_dbl_dnrm), .B(mul_frac_in2[0]), .Z(N497)
         );
  GTECH_AND2 C1259 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N499)
         );
  GTECH_OR2 C1260 ( .A(N500), .B(N501), .Z(m2stg_frac2_array_in[0]) );
  GTECH_AND2 C1261 ( .A(m2stg_frac2_dbl_norm), .B(mul_frac_in2[0]), .Z(N500)
         );
  GTECH_AND2 C1262 ( .A(m2stg_frac2_inf), .B(m1stg_inf_zero_in_dbl), .Z(N501)
         );
  GTECH_OR2 C1263 ( .A(N502), .B(N503), .Z(m1stg_ld0_1_din[52]) );
  GTECH_AND2 C1264 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[54]), .Z(N502) );
  GTECH_AND2 C1265 ( .A(m1stg_dblop), .B(mul_frac_in1[51]), .Z(N503) );
  GTECH_OR2 C1266 ( .A(N504), .B(N505), .Z(m1stg_ld0_1_din[51]) );
  GTECH_AND2 C1267 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[53]), .Z(N504) );
  GTECH_AND2 C1268 ( .A(m1stg_dblop), .B(mul_frac_in1[50]), .Z(N505) );
  GTECH_OR2 C1269 ( .A(N506), .B(N507), .Z(m1stg_ld0_1_din[50]) );
  GTECH_AND2 C1270 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[52]), .Z(N506) );
  GTECH_AND2 C1271 ( .A(m1stg_dblop), .B(mul_frac_in1[49]), .Z(N507) );
  GTECH_OR2 C1272 ( .A(N508), .B(N509), .Z(m1stg_ld0_1_din[49]) );
  GTECH_AND2 C1273 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[51]), .Z(N508) );
  GTECH_AND2 C1274 ( .A(m1stg_dblop), .B(mul_frac_in1[48]), .Z(N509) );
  GTECH_OR2 C1275 ( .A(N510), .B(N511), .Z(m1stg_ld0_1_din[48]) );
  GTECH_AND2 C1276 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[50]), .Z(N510) );
  GTECH_AND2 C1277 ( .A(m1stg_dblop), .B(mul_frac_in1[47]), .Z(N511) );
  GTECH_OR2 C1278 ( .A(N512), .B(N513), .Z(m1stg_ld0_1_din[47]) );
  GTECH_AND2 C1279 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[49]), .Z(N512) );
  GTECH_AND2 C1280 ( .A(m1stg_dblop), .B(mul_frac_in1[46]), .Z(N513) );
  GTECH_OR2 C1281 ( .A(N514), .B(N515), .Z(m1stg_ld0_1_din[46]) );
  GTECH_AND2 C1282 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[48]), .Z(N514) );
  GTECH_AND2 C1283 ( .A(m1stg_dblop), .B(mul_frac_in1[45]), .Z(N515) );
  GTECH_OR2 C1284 ( .A(N516), .B(N517), .Z(m1stg_ld0_1_din[45]) );
  GTECH_AND2 C1285 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[47]), .Z(N516) );
  GTECH_AND2 C1286 ( .A(m1stg_dblop), .B(mul_frac_in1[44]), .Z(N517) );
  GTECH_OR2 C1287 ( .A(N518), .B(N519), .Z(m1stg_ld0_1_din[44]) );
  GTECH_AND2 C1288 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[46]), .Z(N518) );
  GTECH_AND2 C1289 ( .A(m1stg_dblop), .B(mul_frac_in1[43]), .Z(N519) );
  GTECH_OR2 C1290 ( .A(N520), .B(N521), .Z(m1stg_ld0_1_din[43]) );
  GTECH_AND2 C1291 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[45]), .Z(N520) );
  GTECH_AND2 C1292 ( .A(m1stg_dblop), .B(mul_frac_in1[42]), .Z(N521) );
  GTECH_OR2 C1293 ( .A(N522), .B(N523), .Z(m1stg_ld0_1_din[42]) );
  GTECH_AND2 C1294 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[44]), .Z(N522) );
  GTECH_AND2 C1295 ( .A(m1stg_dblop), .B(mul_frac_in1[41]), .Z(N523) );
  GTECH_OR2 C1296 ( .A(N524), .B(N525), .Z(m1stg_ld0_1_din[41]) );
  GTECH_AND2 C1297 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[43]), .Z(N524) );
  GTECH_AND2 C1298 ( .A(m1stg_dblop), .B(mul_frac_in1[40]), .Z(N525) );
  GTECH_OR2 C1299 ( .A(N526), .B(N527), .Z(m1stg_ld0_1_din[40]) );
  GTECH_AND2 C1300 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[42]), .Z(N526) );
  GTECH_AND2 C1301 ( .A(m1stg_dblop), .B(mul_frac_in1[39]), .Z(N527) );
  GTECH_OR2 C1302 ( .A(N528), .B(N529), .Z(m1stg_ld0_1_din[39]) );
  GTECH_AND2 C1303 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[41]), .Z(N528) );
  GTECH_AND2 C1304 ( .A(m1stg_dblop), .B(mul_frac_in1[38]), .Z(N529) );
  GTECH_OR2 C1305 ( .A(N530), .B(N531), .Z(m1stg_ld0_1_din[38]) );
  GTECH_AND2 C1306 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[40]), .Z(N530) );
  GTECH_AND2 C1307 ( .A(m1stg_dblop), .B(mul_frac_in1[37]), .Z(N531) );
  GTECH_OR2 C1308 ( .A(N532), .B(N533), .Z(m1stg_ld0_1_din[37]) );
  GTECH_AND2 C1309 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[39]), .Z(N532) );
  GTECH_AND2 C1310 ( .A(m1stg_dblop), .B(mul_frac_in1[36]), .Z(N533) );
  GTECH_OR2 C1311 ( .A(N534), .B(N535), .Z(m1stg_ld0_1_din[36]) );
  GTECH_AND2 C1312 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[38]), .Z(N534) );
  GTECH_AND2 C1313 ( .A(m1stg_dblop), .B(mul_frac_in1[35]), .Z(N535) );
  GTECH_OR2 C1314 ( .A(N536), .B(N537), .Z(m1stg_ld0_1_din[35]) );
  GTECH_AND2 C1315 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[37]), .Z(N536) );
  GTECH_AND2 C1316 ( .A(m1stg_dblop), .B(mul_frac_in1[34]), .Z(N537) );
  GTECH_OR2 C1317 ( .A(N538), .B(N539), .Z(m1stg_ld0_1_din[34]) );
  GTECH_AND2 C1318 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[36]), .Z(N538) );
  GTECH_AND2 C1319 ( .A(m1stg_dblop), .B(mul_frac_in1[33]), .Z(N539) );
  GTECH_OR2 C1320 ( .A(N540), .B(N541), .Z(m1stg_ld0_1_din[33]) );
  GTECH_AND2 C1321 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[35]), .Z(N540) );
  GTECH_AND2 C1322 ( .A(m1stg_dblop), .B(mul_frac_in1[32]), .Z(N541) );
  GTECH_OR2 C1323 ( .A(N542), .B(N543), .Z(m1stg_ld0_1_din[32]) );
  GTECH_AND2 C1324 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[34]), .Z(N542) );
  GTECH_AND2 C1325 ( .A(m1stg_dblop), .B(mul_frac_in1[31]), .Z(N543) );
  GTECH_OR2 C1326 ( .A(N544), .B(N545), .Z(m1stg_ld0_1_din[31]) );
  GTECH_AND2 C1327 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[33]), .Z(N544) );
  GTECH_AND2 C1328 ( .A(m1stg_dblop), .B(mul_frac_in1[30]), .Z(N545) );
  GTECH_OR2 C1329 ( .A(N546), .B(N547), .Z(m1stg_ld0_1_din[30]) );
  GTECH_AND2 C1330 ( .A(m1stg_dblop_inv), .B(mul_frac_in1[32]), .Z(N546) );
  GTECH_AND2 C1331 ( .A(m1stg_dblop), .B(mul_frac_in1[29]), .Z(N547) );
  GTECH_AND2 C1332 ( .A(m1stg_dblop), .B(mul_frac_in1[28]), .Z(
        m1stg_ld0_1_din[29]) );
  GTECH_AND2 C1333 ( .A(m1stg_dblop), .B(mul_frac_in1[27]), .Z(
        m1stg_ld0_1_din[28]) );
  GTECH_AND2 C1334 ( .A(m1stg_dblop), .B(mul_frac_in1[26]), .Z(
        m1stg_ld0_1_din[27]) );
  GTECH_AND2 C1335 ( .A(m1stg_dblop), .B(mul_frac_in1[25]), .Z(
        m1stg_ld0_1_din[26]) );
  GTECH_AND2 C1336 ( .A(m1stg_dblop), .B(mul_frac_in1[24]), .Z(
        m1stg_ld0_1_din[25]) );
  GTECH_AND2 C1337 ( .A(m1stg_dblop), .B(mul_frac_in1[23]), .Z(
        m1stg_ld0_1_din[24]) );
  GTECH_AND2 C1338 ( .A(m1stg_dblop), .B(mul_frac_in1[22]), .Z(
        m1stg_ld0_1_din[23]) );
  GTECH_AND2 C1339 ( .A(m1stg_dblop), .B(mul_frac_in1[21]), .Z(
        m1stg_ld0_1_din[22]) );
  GTECH_AND2 C1340 ( .A(m1stg_dblop), .B(mul_frac_in1[20]), .Z(
        m1stg_ld0_1_din[21]) );
  GTECH_AND2 C1341 ( .A(m1stg_dblop), .B(mul_frac_in1[19]), .Z(
        m1stg_ld0_1_din[20]) );
  GTECH_AND2 C1342 ( .A(m1stg_dblop), .B(mul_frac_in1[18]), .Z(
        m1stg_ld0_1_din[19]) );
  GTECH_AND2 C1343 ( .A(m1stg_dblop), .B(mul_frac_in1[17]), .Z(
        m1stg_ld0_1_din[18]) );
  GTECH_AND2 C1344 ( .A(m1stg_dblop), .B(mul_frac_in1[16]), .Z(
        m1stg_ld0_1_din[17]) );
  GTECH_AND2 C1345 ( .A(m1stg_dblop), .B(mul_frac_in1[15]), .Z(
        m1stg_ld0_1_din[16]) );
  GTECH_AND2 C1346 ( .A(m1stg_dblop), .B(mul_frac_in1[14]), .Z(
        m1stg_ld0_1_din[15]) );
  GTECH_AND2 C1347 ( .A(m1stg_dblop), .B(mul_frac_in1[13]), .Z(
        m1stg_ld0_1_din[14]) );
  GTECH_AND2 C1348 ( .A(m1stg_dblop), .B(mul_frac_in1[12]), .Z(
        m1stg_ld0_1_din[13]) );
  GTECH_AND2 C1349 ( .A(m1stg_dblop), .B(mul_frac_in1[11]), .Z(
        m1stg_ld0_1_din[12]) );
  GTECH_AND2 C1350 ( .A(m1stg_dblop), .B(mul_frac_in1[10]), .Z(
        m1stg_ld0_1_din[11]) );
  GTECH_AND2 C1351 ( .A(m1stg_dblop), .B(mul_frac_in1[9]), .Z(
        m1stg_ld0_1_din[10]) );
  GTECH_AND2 C1352 ( .A(m1stg_dblop), .B(mul_frac_in1[8]), .Z(
        m1stg_ld0_1_din[9]) );
  GTECH_AND2 C1353 ( .A(m1stg_dblop), .B(mul_frac_in1[7]), .Z(
        m1stg_ld0_1_din[8]) );
  GTECH_AND2 C1354 ( .A(m1stg_dblop), .B(mul_frac_in1[6]), .Z(
        m1stg_ld0_1_din[7]) );
  GTECH_AND2 C1355 ( .A(m1stg_dblop), .B(mul_frac_in1[5]), .Z(
        m1stg_ld0_1_din[6]) );
  GTECH_AND2 C1356 ( .A(m1stg_dblop), .B(mul_frac_in1[4]), .Z(
        m1stg_ld0_1_din[5]) );
  GTECH_AND2 C1357 ( .A(m1stg_dblop), .B(mul_frac_in1[3]), .Z(
        m1stg_ld0_1_din[4]) );
  GTECH_AND2 C1358 ( .A(m1stg_dblop), .B(mul_frac_in1[2]), .Z(
        m1stg_ld0_1_din[3]) );
  GTECH_AND2 C1359 ( .A(m1stg_dblop), .B(mul_frac_in1[1]), .Z(
        m1stg_ld0_1_din[2]) );
  GTECH_AND2 C1360 ( .A(m1stg_dblop), .B(mul_frac_in1[0]), .Z(
        m1stg_ld0_1_din[1]) );
  GTECH_OR2 C1361 ( .A(N548), .B(N549), .Z(m1stg_ld0_2_din[52]) );
  GTECH_AND2 C1362 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[54]), .Z(N548) );
  GTECH_AND2 C1363 ( .A(m1stg_dblop), .B(mul_frac_in2[51]), .Z(N549) );
  GTECH_OR2 C1364 ( .A(N550), .B(N551), .Z(m1stg_ld0_2_din[51]) );
  GTECH_AND2 C1365 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[53]), .Z(N550) );
  GTECH_AND2 C1366 ( .A(m1stg_dblop), .B(mul_frac_in2[50]), .Z(N551) );
  GTECH_OR2 C1367 ( .A(N552), .B(N553), .Z(m1stg_ld0_2_din[50]) );
  GTECH_AND2 C1368 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[52]), .Z(N552) );
  GTECH_AND2 C1369 ( .A(m1stg_dblop), .B(mul_frac_in2[49]), .Z(N553) );
  GTECH_OR2 C1370 ( .A(N554), .B(N555), .Z(m1stg_ld0_2_din[49]) );
  GTECH_AND2 C1371 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[51]), .Z(N554) );
  GTECH_AND2 C1372 ( .A(m1stg_dblop), .B(mul_frac_in2[48]), .Z(N555) );
  GTECH_OR2 C1373 ( .A(N556), .B(N557), .Z(m1stg_ld0_2_din[48]) );
  GTECH_AND2 C1374 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[50]), .Z(N556) );
  GTECH_AND2 C1375 ( .A(m1stg_dblop), .B(mul_frac_in2[47]), .Z(N557) );
  GTECH_OR2 C1376 ( .A(N558), .B(N559), .Z(m1stg_ld0_2_din[47]) );
  GTECH_AND2 C1377 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[49]), .Z(N558) );
  GTECH_AND2 C1378 ( .A(m1stg_dblop), .B(mul_frac_in2[46]), .Z(N559) );
  GTECH_OR2 C1379 ( .A(N560), .B(N561), .Z(m1stg_ld0_2_din[46]) );
  GTECH_AND2 C1380 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[48]), .Z(N560) );
  GTECH_AND2 C1381 ( .A(m1stg_dblop), .B(mul_frac_in2[45]), .Z(N561) );
  GTECH_OR2 C1382 ( .A(N562), .B(N563), .Z(m1stg_ld0_2_din[45]) );
  GTECH_AND2 C1383 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[47]), .Z(N562) );
  GTECH_AND2 C1384 ( .A(m1stg_dblop), .B(mul_frac_in2[44]), .Z(N563) );
  GTECH_OR2 C1385 ( .A(N564), .B(N565), .Z(m1stg_ld0_2_din[44]) );
  GTECH_AND2 C1386 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[46]), .Z(N564) );
  GTECH_AND2 C1387 ( .A(m1stg_dblop), .B(mul_frac_in2[43]), .Z(N565) );
  GTECH_OR2 C1388 ( .A(N566), .B(N567), .Z(m1stg_ld0_2_din[43]) );
  GTECH_AND2 C1389 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[45]), .Z(N566) );
  GTECH_AND2 C1390 ( .A(m1stg_dblop), .B(mul_frac_in2[42]), .Z(N567) );
  GTECH_OR2 C1391 ( .A(N568), .B(N569), .Z(m1stg_ld0_2_din[42]) );
  GTECH_AND2 C1392 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[44]), .Z(N568) );
  GTECH_AND2 C1393 ( .A(m1stg_dblop), .B(mul_frac_in2[41]), .Z(N569) );
  GTECH_OR2 C1394 ( .A(N570), .B(N571), .Z(m1stg_ld0_2_din[41]) );
  GTECH_AND2 C1395 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[43]), .Z(N570) );
  GTECH_AND2 C1396 ( .A(m1stg_dblop), .B(mul_frac_in2[40]), .Z(N571) );
  GTECH_OR2 C1397 ( .A(N572), .B(N573), .Z(m1stg_ld0_2_din[40]) );
  GTECH_AND2 C1398 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[42]), .Z(N572) );
  GTECH_AND2 C1399 ( .A(m1stg_dblop), .B(mul_frac_in2[39]), .Z(N573) );
  GTECH_OR2 C1400 ( .A(N574), .B(N575), .Z(m1stg_ld0_2_din[39]) );
  GTECH_AND2 C1401 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[41]), .Z(N574) );
  GTECH_AND2 C1402 ( .A(m1stg_dblop), .B(mul_frac_in2[38]), .Z(N575) );
  GTECH_OR2 C1403 ( .A(N576), .B(N577), .Z(m1stg_ld0_2_din[38]) );
  GTECH_AND2 C1404 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[40]), .Z(N576) );
  GTECH_AND2 C1405 ( .A(m1stg_dblop), .B(mul_frac_in2[37]), .Z(N577) );
  GTECH_OR2 C1406 ( .A(N578), .B(N579), .Z(m1stg_ld0_2_din[37]) );
  GTECH_AND2 C1407 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[39]), .Z(N578) );
  GTECH_AND2 C1408 ( .A(m1stg_dblop), .B(mul_frac_in2[36]), .Z(N579) );
  GTECH_OR2 C1409 ( .A(N580), .B(N581), .Z(m1stg_ld0_2_din[36]) );
  GTECH_AND2 C1410 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[38]), .Z(N580) );
  GTECH_AND2 C1411 ( .A(m1stg_dblop), .B(mul_frac_in2[35]), .Z(N581) );
  GTECH_OR2 C1412 ( .A(N582), .B(N583), .Z(m1stg_ld0_2_din[35]) );
  GTECH_AND2 C1413 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[37]), .Z(N582) );
  GTECH_AND2 C1414 ( .A(m1stg_dblop), .B(mul_frac_in2[34]), .Z(N583) );
  GTECH_OR2 C1415 ( .A(N584), .B(N585), .Z(m1stg_ld0_2_din[34]) );
  GTECH_AND2 C1416 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[36]), .Z(N584) );
  GTECH_AND2 C1417 ( .A(m1stg_dblop), .B(mul_frac_in2[33]), .Z(N585) );
  GTECH_OR2 C1418 ( .A(N586), .B(N587), .Z(m1stg_ld0_2_din[33]) );
  GTECH_AND2 C1419 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[35]), .Z(N586) );
  GTECH_AND2 C1420 ( .A(m1stg_dblop), .B(mul_frac_in2[32]), .Z(N587) );
  GTECH_OR2 C1421 ( .A(N588), .B(N589), .Z(m1stg_ld0_2_din[32]) );
  GTECH_AND2 C1422 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[34]), .Z(N588) );
  GTECH_AND2 C1423 ( .A(m1stg_dblop), .B(mul_frac_in2[31]), .Z(N589) );
  GTECH_OR2 C1424 ( .A(N590), .B(N591), .Z(m1stg_ld0_2_din[31]) );
  GTECH_AND2 C1425 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[33]), .Z(N590) );
  GTECH_AND2 C1426 ( .A(m1stg_dblop), .B(mul_frac_in2[30]), .Z(N591) );
  GTECH_OR2 C1427 ( .A(N592), .B(N593), .Z(m1stg_ld0_2_din[30]) );
  GTECH_AND2 C1428 ( .A(m1stg_dblop_inv), .B(mul_frac_in2[32]), .Z(N592) );
  GTECH_AND2 C1429 ( .A(m1stg_dblop), .B(mul_frac_in2[29]), .Z(N593) );
  GTECH_AND2 C1430 ( .A(m1stg_dblop), .B(mul_frac_in2[28]), .Z(
        m1stg_ld0_2_din[29]) );
  GTECH_AND2 C1431 ( .A(m1stg_dblop), .B(mul_frac_in2[27]), .Z(
        m1stg_ld0_2_din[28]) );
  GTECH_AND2 C1432 ( .A(m1stg_dblop), .B(mul_frac_in2[26]), .Z(
        m1stg_ld0_2_din[27]) );
  GTECH_AND2 C1433 ( .A(m1stg_dblop), .B(mul_frac_in2[25]), .Z(
        m1stg_ld0_2_din[26]) );
  GTECH_AND2 C1434 ( .A(m1stg_dblop), .B(mul_frac_in2[24]), .Z(
        m1stg_ld0_2_din[25]) );
  GTECH_AND2 C1435 ( .A(m1stg_dblop), .B(mul_frac_in2[23]), .Z(
        m1stg_ld0_2_din[24]) );
  GTECH_AND2 C1436 ( .A(m1stg_dblop), .B(mul_frac_in2[22]), .Z(
        m1stg_ld0_2_din[23]) );
  GTECH_AND2 C1437 ( .A(m1stg_dblop), .B(mul_frac_in2[21]), .Z(
        m1stg_ld0_2_din[22]) );
  GTECH_AND2 C1438 ( .A(m1stg_dblop), .B(mul_frac_in2[20]), .Z(
        m1stg_ld0_2_din[21]) );
  GTECH_AND2 C1439 ( .A(m1stg_dblop), .B(mul_frac_in2[19]), .Z(
        m1stg_ld0_2_din[20]) );
  GTECH_AND2 C1440 ( .A(m1stg_dblop), .B(mul_frac_in2[18]), .Z(
        m1stg_ld0_2_din[19]) );
  GTECH_AND2 C1441 ( .A(m1stg_dblop), .B(mul_frac_in2[17]), .Z(
        m1stg_ld0_2_din[18]) );
  GTECH_AND2 C1442 ( .A(m1stg_dblop), .B(mul_frac_in2[16]), .Z(
        m1stg_ld0_2_din[17]) );
  GTECH_AND2 C1443 ( .A(m1stg_dblop), .B(mul_frac_in2[15]), .Z(
        m1stg_ld0_2_din[16]) );
  GTECH_AND2 C1444 ( .A(m1stg_dblop), .B(mul_frac_in2[14]), .Z(
        m1stg_ld0_2_din[15]) );
  GTECH_AND2 C1445 ( .A(m1stg_dblop), .B(mul_frac_in2[13]), .Z(
        m1stg_ld0_2_din[14]) );
  GTECH_AND2 C1446 ( .A(m1stg_dblop), .B(mul_frac_in2[12]), .Z(
        m1stg_ld0_2_din[13]) );
  GTECH_AND2 C1447 ( .A(m1stg_dblop), .B(mul_frac_in2[11]), .Z(
        m1stg_ld0_2_din[12]) );
  GTECH_AND2 C1448 ( .A(m1stg_dblop), .B(mul_frac_in2[10]), .Z(
        m1stg_ld0_2_din[11]) );
  GTECH_AND2 C1449 ( .A(m1stg_dblop), .B(mul_frac_in2[9]), .Z(
        m1stg_ld0_2_din[10]) );
  GTECH_AND2 C1450 ( .A(m1stg_dblop), .B(mul_frac_in2[8]), .Z(
        m1stg_ld0_2_din[9]) );
  GTECH_AND2 C1451 ( .A(m1stg_dblop), .B(mul_frac_in2[7]), .Z(
        m1stg_ld0_2_din[8]) );
  GTECH_AND2 C1452 ( .A(m1stg_dblop), .B(mul_frac_in2[6]), .Z(
        m1stg_ld0_2_din[7]) );
  GTECH_AND2 C1453 ( .A(m1stg_dblop), .B(mul_frac_in2[5]), .Z(
        m1stg_ld0_2_din[6]) );
  GTECH_AND2 C1454 ( .A(m1stg_dblop), .B(mul_frac_in2[4]), .Z(
        m1stg_ld0_2_din[5]) );
  GTECH_AND2 C1455 ( .A(m1stg_dblop), .B(mul_frac_in2[3]), .Z(
        m1stg_ld0_2_din[4]) );
  GTECH_AND2 C1456 ( .A(m1stg_dblop), .B(mul_frac_in2[2]), .Z(
        m1stg_ld0_2_din[3]) );
  GTECH_AND2 C1457 ( .A(m1stg_dblop), .B(mul_frac_in2[1]), .Z(
        m1stg_ld0_2_din[2]) );
  GTECH_AND2 C1458 ( .A(m1stg_dblop), .B(mul_frac_in2[0]), .Z(
        m1stg_ld0_2_din[1]) );
  GTECH_OR2 C1459 ( .A(N642), .B(m4stg_shl_tmp[63]), .Z(m4stg_shl[0]) );
  GTECH_OR2 C1460 ( .A(N641), .B(m4stg_shl_tmp[64]), .Z(N642) );
  GTECH_OR2 C1461 ( .A(N640), .B(m4stg_shl_tmp[65]), .Z(N641) );
  GTECH_OR2 C1462 ( .A(N639), .B(m4stg_shl_tmp[66]), .Z(N640) );
  GTECH_OR2 C1463 ( .A(N638), .B(m4stg_shl_tmp[67]), .Z(N639) );
  GTECH_OR2 C1464 ( .A(N637), .B(m4stg_shl_tmp[68]), .Z(N638) );
  GTECH_OR2 C1465 ( .A(N636), .B(m4stg_shl_tmp[69]), .Z(N637) );
  GTECH_OR2 C1466 ( .A(N635), .B(m4stg_shl_tmp[70]), .Z(N636) );
  GTECH_OR2 C1467 ( .A(N634), .B(m4stg_shl_tmp[71]), .Z(N635) );
  GTECH_OR2 C1468 ( .A(N633), .B(m4stg_shl_tmp[72]), .Z(N634) );
  GTECH_OR2 C1469 ( .A(N632), .B(m4stg_shl_tmp[73]), .Z(N633) );
  GTECH_OR2 C1470 ( .A(N631), .B(m4stg_shl_tmp[74]), .Z(N632) );
  GTECH_OR2 C1471 ( .A(N630), .B(m4stg_shl_tmp[75]), .Z(N631) );
  GTECH_OR2 C1472 ( .A(N629), .B(m4stg_shl_tmp[76]), .Z(N630) );
  GTECH_OR2 C1473 ( .A(N628), .B(m4stg_shl_tmp[77]), .Z(N629) );
  GTECH_OR2 C1474 ( .A(N627), .B(m4stg_shl_tmp[78]), .Z(N628) );
  GTECH_OR2 C1475 ( .A(N626), .B(m4stg_shl_tmp[79]), .Z(N627) );
  GTECH_OR2 C1476 ( .A(N625), .B(m4stg_shl_tmp[80]), .Z(N626) );
  GTECH_OR2 C1477 ( .A(N624), .B(m4stg_shl_tmp[81]), .Z(N625) );
  GTECH_OR2 C1478 ( .A(N623), .B(m4stg_shl_tmp[82]), .Z(N624) );
  GTECH_OR2 C1479 ( .A(N622), .B(m4stg_shl_tmp[83]), .Z(N623) );
  GTECH_OR2 C1480 ( .A(N621), .B(m4stg_shl_tmp[84]), .Z(N622) );
  GTECH_OR2 C1481 ( .A(N620), .B(m4stg_shl_tmp[85]), .Z(N621) );
  GTECH_OR2 C1482 ( .A(N619), .B(m4stg_shl_tmp[86]), .Z(N620) );
  GTECH_OR2 C1483 ( .A(N618), .B(m4stg_shl_tmp[87]), .Z(N619) );
  GTECH_OR2 C1484 ( .A(N617), .B(m4stg_shl_tmp[88]), .Z(N618) );
  GTECH_OR2 C1485 ( .A(N616), .B(m4stg_shl_tmp[89]), .Z(N617) );
  GTECH_OR2 C1486 ( .A(N615), .B(m4stg_shl_tmp[90]), .Z(N616) );
  GTECH_OR2 C1487 ( .A(N614), .B(m4stg_shl_tmp[91]), .Z(N615) );
  GTECH_OR2 C1488 ( .A(N613), .B(m4stg_shl_tmp[92]), .Z(N614) );
  GTECH_OR2 C1489 ( .A(N612), .B(m4stg_shl_tmp[93]), .Z(N613) );
  GTECH_OR2 C1490 ( .A(N611), .B(m4stg_shl_tmp[94]), .Z(N612) );
  GTECH_OR2 C1491 ( .A(N610), .B(m4stg_shl_tmp[95]), .Z(N611) );
  GTECH_OR2 C1492 ( .A(N609), .B(m4stg_shl_tmp[96]), .Z(N610) );
  GTECH_OR2 C1493 ( .A(N608), .B(m4stg_shl_tmp[97]), .Z(N609) );
  GTECH_OR2 C1494 ( .A(N607), .B(m4stg_shl_tmp[98]), .Z(N608) );
  GTECH_OR2 C1495 ( .A(N606), .B(m4stg_shl_tmp[99]), .Z(N607) );
  GTECH_OR2 C1496 ( .A(N605), .B(m4stg_shl_tmp[100]), .Z(N606) );
  GTECH_OR2 C1497 ( .A(N604), .B(m4stg_shl_tmp[101]), .Z(N605) );
  GTECH_OR2 C1498 ( .A(N603), .B(m4stg_shl_tmp[102]), .Z(N604) );
  GTECH_OR2 C1499 ( .A(N602), .B(m4stg_shl_tmp[103]), .Z(N603) );
  GTECH_OR2 C1500 ( .A(N601), .B(m4stg_shl_tmp[104]), .Z(N602) );
  GTECH_OR2 C1501 ( .A(N600), .B(m4stg_shl_tmp[105]), .Z(N601) );
  GTECH_OR2 C1502 ( .A(N599), .B(m4stg_shl_tmp[106]), .Z(N600) );
  GTECH_OR2 C1503 ( .A(N598), .B(m4stg_shl_tmp[107]), .Z(N599) );
  GTECH_OR2 C1504 ( .A(N597), .B(m4stg_shl_tmp[108]), .Z(N598) );
  GTECH_OR2 C1505 ( .A(N596), .B(m4stg_shl_tmp[109]), .Z(N597) );
  GTECH_OR2 C1506 ( .A(N595), .B(m4stg_shl_tmp[110]), .Z(N596) );
  GTECH_OR2 C1507 ( .A(N594), .B(m4stg_shl_tmp[111]), .Z(N595) );
  GTECH_OR2 C1508 ( .A(m4stg_shl_tmp[113]), .B(m4stg_shl_tmp[112]), .Z(N594)
         );
  GTECH_OR2 C1509 ( .A(N754), .B(m4stg_shr_tmp[0]), .Z(m4stg_shr[0]) );
  GTECH_OR2 C1510 ( .A(N753), .B(m4stg_shr_tmp[1]), .Z(N754) );
  GTECH_OR2 C1511 ( .A(N752), .B(m4stg_shr_tmp[2]), .Z(N753) );
  GTECH_OR2 C1512 ( .A(N751), .B(m4stg_shr_tmp[3]), .Z(N752) );
  GTECH_OR2 C1513 ( .A(N750), .B(m4stg_shr_tmp[4]), .Z(N751) );
  GTECH_OR2 C1514 ( .A(N749), .B(m4stg_shr_tmp[5]), .Z(N750) );
  GTECH_OR2 C1515 ( .A(N748), .B(m4stg_shr_tmp[6]), .Z(N749) );
  GTECH_OR2 C1516 ( .A(N747), .B(m4stg_shr_tmp[7]), .Z(N748) );
  GTECH_OR2 C1517 ( .A(N746), .B(m4stg_shr_tmp[8]), .Z(N747) );
  GTECH_OR2 C1518 ( .A(N745), .B(m4stg_shr_tmp[9]), .Z(N746) );
  GTECH_OR2 C1519 ( .A(N744), .B(m4stg_shr_tmp[10]), .Z(N745) );
  GTECH_OR2 C1520 ( .A(N743), .B(m4stg_shr_tmp[11]), .Z(N744) );
  GTECH_OR2 C1521 ( .A(N742), .B(m4stg_shr_tmp[12]), .Z(N743) );
  GTECH_OR2 C1522 ( .A(N741), .B(m4stg_shr_tmp[13]), .Z(N742) );
  GTECH_OR2 C1523 ( .A(N740), .B(m4stg_shr_tmp[14]), .Z(N741) );
  GTECH_OR2 C1524 ( .A(N739), .B(m4stg_shr_tmp[15]), .Z(N740) );
  GTECH_OR2 C1525 ( .A(N738), .B(m4stg_shr_tmp[16]), .Z(N739) );
  GTECH_OR2 C1526 ( .A(N737), .B(m4stg_shr_tmp[17]), .Z(N738) );
  GTECH_OR2 C1527 ( .A(N736), .B(m4stg_shr_tmp[18]), .Z(N737) );
  GTECH_OR2 C1528 ( .A(N735), .B(m4stg_shr_tmp[19]), .Z(N736) );
  GTECH_OR2 C1529 ( .A(N734), .B(m4stg_shr_tmp[20]), .Z(N735) );
  GTECH_OR2 C1530 ( .A(N733), .B(m4stg_shr_tmp[21]), .Z(N734) );
  GTECH_OR2 C1531 ( .A(N732), .B(m4stg_shr_tmp[22]), .Z(N733) );
  GTECH_OR2 C1532 ( .A(N731), .B(m4stg_shr_tmp[23]), .Z(N732) );
  GTECH_OR2 C1533 ( .A(N730), .B(m4stg_shr_tmp[24]), .Z(N731) );
  GTECH_OR2 C1534 ( .A(N729), .B(m4stg_shr_tmp[25]), .Z(N730) );
  GTECH_OR2 C1535 ( .A(N728), .B(m4stg_shr_tmp[26]), .Z(N729) );
  GTECH_OR2 C1536 ( .A(N727), .B(m4stg_shr_tmp[27]), .Z(N728) );
  GTECH_OR2 C1537 ( .A(N726), .B(m4stg_shr_tmp[28]), .Z(N727) );
  GTECH_OR2 C1538 ( .A(N725), .B(m4stg_shr_tmp[29]), .Z(N726) );
  GTECH_OR2 C1539 ( .A(N724), .B(m4stg_shr_tmp[30]), .Z(N725) );
  GTECH_OR2 C1540 ( .A(N723), .B(m4stg_shr_tmp[31]), .Z(N724) );
  GTECH_OR2 C1541 ( .A(N722), .B(m4stg_shr_tmp[32]), .Z(N723) );
  GTECH_OR2 C1542 ( .A(N721), .B(m4stg_shr_tmp[33]), .Z(N722) );
  GTECH_OR2 C1543 ( .A(N720), .B(m4stg_shr_tmp[34]), .Z(N721) );
  GTECH_OR2 C1544 ( .A(N719), .B(m4stg_shr_tmp[35]), .Z(N720) );
  GTECH_OR2 C1545 ( .A(N718), .B(m4stg_shr_tmp[36]), .Z(N719) );
  GTECH_OR2 C1546 ( .A(N717), .B(m4stg_shr_tmp[37]), .Z(N718) );
  GTECH_OR2 C1547 ( .A(N716), .B(m4stg_shr_tmp[38]), .Z(N717) );
  GTECH_OR2 C1548 ( .A(N715), .B(m4stg_shr_tmp[39]), .Z(N716) );
  GTECH_OR2 C1549 ( .A(N714), .B(m4stg_shr_tmp[40]), .Z(N715) );
  GTECH_OR2 C1550 ( .A(N713), .B(m4stg_shr_tmp[41]), .Z(N714) );
  GTECH_OR2 C1551 ( .A(N712), .B(m4stg_shr_tmp[42]), .Z(N713) );
  GTECH_OR2 C1552 ( .A(N711), .B(m4stg_shr_tmp[43]), .Z(N712) );
  GTECH_OR2 C1553 ( .A(N710), .B(m4stg_shr_tmp[44]), .Z(N711) );
  GTECH_OR2 C1554 ( .A(N709), .B(m4stg_shr_tmp[45]), .Z(N710) );
  GTECH_OR2 C1555 ( .A(N708), .B(m4stg_shr_tmp[46]), .Z(N709) );
  GTECH_OR2 C1556 ( .A(N707), .B(m4stg_shr_tmp[47]), .Z(N708) );
  GTECH_OR2 C1557 ( .A(N706), .B(m4stg_shr_tmp[48]), .Z(N707) );
  GTECH_OR2 C1558 ( .A(N705), .B(m4stg_shr_tmp[49]), .Z(N706) );
  GTECH_OR2 C1559 ( .A(N704), .B(m4stg_shr_tmp[50]), .Z(N705) );
  GTECH_OR2 C1560 ( .A(N703), .B(m4stg_shr_tmp[51]), .Z(N704) );
  GTECH_OR2 C1561 ( .A(N702), .B(m4stg_shr_tmp[52]), .Z(N703) );
  GTECH_OR2 C1562 ( .A(N701), .B(m4stg_shr_tmp[53]), .Z(N702) );
  GTECH_OR2 C1563 ( .A(N700), .B(m4stg_shr_tmp[54]), .Z(N701) );
  GTECH_OR2 C1564 ( .A(N699), .B(m4stg_shr_tmp[55]), .Z(N700) );
  GTECH_OR2 C1565 ( .A(N698), .B(m4stg_shr_tmp[56]), .Z(N699) );
  GTECH_OR2 C1566 ( .A(N697), .B(m4stg_shr_tmp[57]), .Z(N698) );
  GTECH_OR2 C1567 ( .A(N696), .B(m4stg_shr_tmp[58]), .Z(N697) );
  GTECH_OR2 C1568 ( .A(N695), .B(m4stg_shr_tmp[59]), .Z(N696) );
  GTECH_OR2 C1569 ( .A(N694), .B(m4stg_shr_tmp[60]), .Z(N695) );
  GTECH_OR2 C1570 ( .A(N693), .B(m4stg_shr_tmp[61]), .Z(N694) );
  GTECH_OR2 C1571 ( .A(N692), .B(m4stg_shr_tmp[62]), .Z(N693) );
  GTECH_OR2 C1572 ( .A(N691), .B(m4stg_shr_tmp[63]), .Z(N692) );
  GTECH_OR2 C1573 ( .A(N690), .B(m4stg_shr_tmp[64]), .Z(N691) );
  GTECH_OR2 C1574 ( .A(N689), .B(m4stg_shr_tmp[65]), .Z(N690) );
  GTECH_OR2 C1575 ( .A(N688), .B(m4stg_shr_tmp[66]), .Z(N689) );
  GTECH_OR2 C1576 ( .A(N687), .B(m4stg_shr_tmp[67]), .Z(N688) );
  GTECH_OR2 C1577 ( .A(N686), .B(m4stg_shr_tmp[68]), .Z(N687) );
  GTECH_OR2 C1578 ( .A(N685), .B(m4stg_shr_tmp[69]), .Z(N686) );
  GTECH_OR2 C1579 ( .A(N684), .B(m4stg_shr_tmp[70]), .Z(N685) );
  GTECH_OR2 C1580 ( .A(N683), .B(m4stg_shr_tmp[71]), .Z(N684) );
  GTECH_OR2 C1581 ( .A(N682), .B(m4stg_shr_tmp[72]), .Z(N683) );
  GTECH_OR2 C1582 ( .A(N681), .B(m4stg_shr_tmp[73]), .Z(N682) );
  GTECH_OR2 C1583 ( .A(N680), .B(m4stg_shr_tmp[74]), .Z(N681) );
  GTECH_OR2 C1584 ( .A(N679), .B(m4stg_shr_tmp[75]), .Z(N680) );
  GTECH_OR2 C1585 ( .A(N678), .B(m4stg_shr_tmp[76]), .Z(N679) );
  GTECH_OR2 C1586 ( .A(N677), .B(m4stg_shr_tmp[77]), .Z(N678) );
  GTECH_OR2 C1587 ( .A(N676), .B(m4stg_shr_tmp[78]), .Z(N677) );
  GTECH_OR2 C1588 ( .A(N675), .B(m4stg_shr_tmp[79]), .Z(N676) );
  GTECH_OR2 C1589 ( .A(N674), .B(m4stg_shr_tmp[80]), .Z(N675) );
  GTECH_OR2 C1590 ( .A(N673), .B(m4stg_shr_tmp[81]), .Z(N674) );
  GTECH_OR2 C1591 ( .A(N672), .B(m4stg_shr_tmp[82]), .Z(N673) );
  GTECH_OR2 C1592 ( .A(N671), .B(m4stg_shr_tmp[83]), .Z(N672) );
  GTECH_OR2 C1593 ( .A(N670), .B(m4stg_shr_tmp[84]), .Z(N671) );
  GTECH_OR2 C1594 ( .A(N669), .B(m4stg_shr_tmp[85]), .Z(N670) );
  GTECH_OR2 C1595 ( .A(N668), .B(m4stg_shr_tmp[86]), .Z(N669) );
  GTECH_OR2 C1596 ( .A(N667), .B(m4stg_shr_tmp[87]), .Z(N668) );
  GTECH_OR2 C1597 ( .A(N666), .B(m4stg_shr_tmp[88]), .Z(N667) );
  GTECH_OR2 C1598 ( .A(N665), .B(m4stg_shr_tmp[89]), .Z(N666) );
  GTECH_OR2 C1599 ( .A(N664), .B(m4stg_shr_tmp[90]), .Z(N665) );
  GTECH_OR2 C1600 ( .A(N663), .B(m4stg_shr_tmp[91]), .Z(N664) );
  GTECH_OR2 C1601 ( .A(N662), .B(m4stg_shr_tmp[92]), .Z(N663) );
  GTECH_OR2 C1602 ( .A(N661), .B(m4stg_shr_tmp[93]), .Z(N662) );
  GTECH_OR2 C1603 ( .A(N660), .B(m4stg_shr_tmp[94]), .Z(N661) );
  GTECH_OR2 C1604 ( .A(N659), .B(m4stg_shr_tmp[95]), .Z(N660) );
  GTECH_OR2 C1605 ( .A(N658), .B(m4stg_shr_tmp[96]), .Z(N659) );
  GTECH_OR2 C1606 ( .A(N657), .B(m4stg_shr_tmp[97]), .Z(N658) );
  GTECH_OR2 C1607 ( .A(N656), .B(m4stg_shr_tmp[98]), .Z(N657) );
  GTECH_OR2 C1608 ( .A(N655), .B(m4stg_shr_tmp[99]), .Z(N656) );
  GTECH_OR2 C1609 ( .A(N654), .B(m4stg_shr_tmp[100]), .Z(N655) );
  GTECH_OR2 C1610 ( .A(N653), .B(m4stg_shr_tmp[101]), .Z(N654) );
  GTECH_OR2 C1611 ( .A(N652), .B(m4stg_shr_tmp[102]), .Z(N653) );
  GTECH_OR2 C1612 ( .A(N651), .B(m4stg_shr_tmp[103]), .Z(N652) );
  GTECH_OR2 C1613 ( .A(N650), .B(m4stg_shr_tmp[104]), .Z(N651) );
  GTECH_OR2 C1614 ( .A(N649), .B(m4stg_shr_tmp[105]), .Z(N650) );
  GTECH_OR2 C1615 ( .A(N648), .B(m4stg_shr_tmp[106]), .Z(N649) );
  GTECH_OR2 C1616 ( .A(N647), .B(m4stg_shr_tmp[107]), .Z(N648) );
  GTECH_OR2 C1617 ( .A(N646), .B(m4stg_shr_tmp[108]), .Z(N647) );
  GTECH_OR2 C1618 ( .A(N645), .B(m4stg_shr_tmp[109]), .Z(N646) );
  GTECH_OR2 C1619 ( .A(N644), .B(m4stg_shr_tmp[110]), .Z(N645) );
  GTECH_OR2 C1620 ( .A(N643), .B(m4stg_shr_tmp[111]), .Z(N644) );
  GTECH_OR2 C1621 ( .A(m4stg_shr_tmp[113]), .B(m4stg_shr_tmp[112]), .Z(N643)
         );
  GTECH_NOT I_54 ( .A(N759), .Z(m5stg_frac_pre1_in[54]) );
  GTECH_OR2 C1623 ( .A(N756), .B(N758), .Z(N759) );
  GTECH_AND2 C1624 ( .A(N755), .B(m4stg_shl_54), .Z(N756) );
  GTECH_AND2 C1625 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N755) );
  GTECH_AND2 C1626 ( .A(N757), .B(m5stg_frac_54_33[54]), .Z(N758) );
  GTECH_NOT I_55 ( .A(m6stg_step), .Z(N757) );
  GTECH_NOT I_56 ( .A(N764), .Z(m5stg_frac_pre1_in[53]) );
  GTECH_OR2 C1629 ( .A(N761), .B(N763), .Z(N764) );
  GTECH_AND2 C1630 ( .A(N760), .B(m4stg_shl_tmp[166]), .Z(N761) );
  GTECH_AND2 C1631 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N760) );
  GTECH_AND2 C1632 ( .A(N762), .B(m5stg_frac_54_33[53]), .Z(N763) );
  GTECH_NOT I_57 ( .A(m6stg_step), .Z(N762) );
  GTECH_NOT I_58 ( .A(N769), .Z(m5stg_frac_pre1_in[52]) );
  GTECH_OR2 C1635 ( .A(N766), .B(N768), .Z(N769) );
  GTECH_AND2 C1636 ( .A(N765), .B(m4stg_shl_tmp[165]), .Z(N766) );
  GTECH_AND2 C1637 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N765) );
  GTECH_AND2 C1638 ( .A(N767), .B(m5stg_frac_54_33[52]), .Z(N768) );
  GTECH_NOT I_59 ( .A(m6stg_step), .Z(N767) );
  GTECH_NOT I_60 ( .A(N774), .Z(m5stg_frac_pre1_in[51]) );
  GTECH_OR2 C1641 ( .A(N771), .B(N773), .Z(N774) );
  GTECH_AND2 C1642 ( .A(N770), .B(m4stg_shl_tmp[164]), .Z(N771) );
  GTECH_AND2 C1643 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N770) );
  GTECH_AND2 C1644 ( .A(N772), .B(m5stg_frac_54_33[51]), .Z(N773) );
  GTECH_NOT I_61 ( .A(m6stg_step), .Z(N772) );
  GTECH_NOT I_62 ( .A(N779), .Z(m5stg_frac_pre1_in[50]) );
  GTECH_OR2 C1647 ( .A(N776), .B(N778), .Z(N779) );
  GTECH_AND2 C1648 ( .A(N775), .B(m4stg_shl_tmp[163]), .Z(N776) );
  GTECH_AND2 C1649 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N775) );
  GTECH_AND2 C1650 ( .A(N777), .B(m5stg_frac_54_33[50]), .Z(N778) );
  GTECH_NOT I_63 ( .A(m6stg_step), .Z(N777) );
  GTECH_NOT I_64 ( .A(N784), .Z(m5stg_frac_pre1_in[49]) );
  GTECH_OR2 C1653 ( .A(N781), .B(N783), .Z(N784) );
  GTECH_AND2 C1654 ( .A(N780), .B(m4stg_shl_tmp[162]), .Z(N781) );
  GTECH_AND2 C1655 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N780) );
  GTECH_AND2 C1656 ( .A(N782), .B(m5stg_frac_54_33[49]), .Z(N783) );
  GTECH_NOT I_65 ( .A(m6stg_step), .Z(N782) );
  GTECH_NOT I_66 ( .A(N789), .Z(m5stg_frac_pre1_in[48]) );
  GTECH_OR2 C1659 ( .A(N786), .B(N788), .Z(N789) );
  GTECH_AND2 C1660 ( .A(N785), .B(m4stg_shl_tmp[161]), .Z(N786) );
  GTECH_AND2 C1661 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N785) );
  GTECH_AND2 C1662 ( .A(N787), .B(m5stg_frac_54_33[48]), .Z(N788) );
  GTECH_NOT I_67 ( .A(m6stg_step), .Z(N787) );
  GTECH_NOT I_68 ( .A(N794), .Z(m5stg_frac_pre1_in[47]) );
  GTECH_OR2 C1665 ( .A(N791), .B(N793), .Z(N794) );
  GTECH_AND2 C1666 ( .A(N790), .B(m4stg_shl_tmp[160]), .Z(N791) );
  GTECH_AND2 C1667 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N790) );
  GTECH_AND2 C1668 ( .A(N792), .B(m5stg_frac_54_33[47]), .Z(N793) );
  GTECH_NOT I_69 ( .A(m6stg_step), .Z(N792) );
  GTECH_NOT I_70 ( .A(N799), .Z(m5stg_frac_pre1_in[46]) );
  GTECH_OR2 C1671 ( .A(N796), .B(N798), .Z(N799) );
  GTECH_AND2 C1672 ( .A(N795), .B(m4stg_shl_tmp[159]), .Z(N796) );
  GTECH_AND2 C1673 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N795) );
  GTECH_AND2 C1674 ( .A(N797), .B(m5stg_frac_54_33[46]), .Z(N798) );
  GTECH_NOT I_71 ( .A(m6stg_step), .Z(N797) );
  GTECH_NOT I_72 ( .A(N804), .Z(m5stg_frac_pre1_in[45]) );
  GTECH_OR2 C1677 ( .A(N801), .B(N803), .Z(N804) );
  GTECH_AND2 C1678 ( .A(N800), .B(m4stg_shl_tmp[158]), .Z(N801) );
  GTECH_AND2 C1679 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N800) );
  GTECH_AND2 C1680 ( .A(N802), .B(m5stg_frac_54_33[45]), .Z(N803) );
  GTECH_NOT I_73 ( .A(m6stg_step), .Z(N802) );
  GTECH_NOT I_74 ( .A(N809), .Z(m5stg_frac_pre1_in[44]) );
  GTECH_OR2 C1683 ( .A(N806), .B(N808), .Z(N809) );
  GTECH_AND2 C1684 ( .A(N805), .B(m4stg_shl_tmp[157]), .Z(N806) );
  GTECH_AND2 C1685 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N805) );
  GTECH_AND2 C1686 ( .A(N807), .B(m5stg_frac_54_33[44]), .Z(N808) );
  GTECH_NOT I_75 ( .A(m6stg_step), .Z(N807) );
  GTECH_NOT I_76 ( .A(N814), .Z(m5stg_frac_pre1_in[43]) );
  GTECH_OR2 C1689 ( .A(N811), .B(N813), .Z(N814) );
  GTECH_AND2 C1690 ( .A(N810), .B(m4stg_shl_tmp[156]), .Z(N811) );
  GTECH_AND2 C1691 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N810) );
  GTECH_AND2 C1692 ( .A(N812), .B(m5stg_frac_54_33[43]), .Z(N813) );
  GTECH_NOT I_77 ( .A(m6stg_step), .Z(N812) );
  GTECH_NOT I_78 ( .A(N819), .Z(m5stg_frac_pre1_in[42]) );
  GTECH_OR2 C1695 ( .A(N816), .B(N818), .Z(N819) );
  GTECH_AND2 C1696 ( .A(N815), .B(m4stg_shl_tmp[155]), .Z(N816) );
  GTECH_AND2 C1697 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N815) );
  GTECH_AND2 C1698 ( .A(N817), .B(m5stg_frac_54_33[42]), .Z(N818) );
  GTECH_NOT I_79 ( .A(m6stg_step), .Z(N817) );
  GTECH_NOT I_80 ( .A(N824), .Z(m5stg_frac_pre1_in[41]) );
  GTECH_OR2 C1701 ( .A(N821), .B(N823), .Z(N824) );
  GTECH_AND2 C1702 ( .A(N820), .B(m4stg_shl_tmp[154]), .Z(N821) );
  GTECH_AND2 C1703 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N820) );
  GTECH_AND2 C1704 ( .A(N822), .B(m5stg_frac_54_33[41]), .Z(N823) );
  GTECH_NOT I_81 ( .A(m6stg_step), .Z(N822) );
  GTECH_NOT I_82 ( .A(N829), .Z(m5stg_frac_pre1_in[40]) );
  GTECH_OR2 C1707 ( .A(N826), .B(N828), .Z(N829) );
  GTECH_AND2 C1708 ( .A(N825), .B(m4stg_shl_tmp[153]), .Z(N826) );
  GTECH_AND2 C1709 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N825) );
  GTECH_AND2 C1710 ( .A(N827), .B(m5stg_frac_54_33[40]), .Z(N828) );
  GTECH_NOT I_83 ( .A(m6stg_step), .Z(N827) );
  GTECH_NOT I_84 ( .A(N834), .Z(m5stg_frac_pre1_in[39]) );
  GTECH_OR2 C1713 ( .A(N831), .B(N833), .Z(N834) );
  GTECH_AND2 C1714 ( .A(N830), .B(m4stg_shl_tmp[152]), .Z(N831) );
  GTECH_AND2 C1715 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N830) );
  GTECH_AND2 C1716 ( .A(N832), .B(m5stg_frac_54_33[39]), .Z(N833) );
  GTECH_NOT I_85 ( .A(m6stg_step), .Z(N832) );
  GTECH_NOT I_86 ( .A(N839), .Z(m5stg_frac_pre1_in[38]) );
  GTECH_OR2 C1719 ( .A(N836), .B(N838), .Z(N839) );
  GTECH_AND2 C1720 ( .A(N835), .B(m4stg_shl_tmp[151]), .Z(N836) );
  GTECH_AND2 C1721 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N835) );
  GTECH_AND2 C1722 ( .A(N837), .B(m5stg_frac_54_33[38]), .Z(N838) );
  GTECH_NOT I_87 ( .A(m6stg_step), .Z(N837) );
  GTECH_NOT I_88 ( .A(N844), .Z(m5stg_frac_pre1_in[37]) );
  GTECH_OR2 C1725 ( .A(N841), .B(N843), .Z(N844) );
  GTECH_AND2 C1726 ( .A(N840), .B(m4stg_shl_tmp[150]), .Z(N841) );
  GTECH_AND2 C1727 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N840) );
  GTECH_AND2 C1728 ( .A(N842), .B(m5stg_frac_54_33[37]), .Z(N843) );
  GTECH_NOT I_89 ( .A(m6stg_step), .Z(N842) );
  GTECH_NOT I_90 ( .A(N849), .Z(m5stg_frac_pre1_in[36]) );
  GTECH_OR2 C1731 ( .A(N846), .B(N848), .Z(N849) );
  GTECH_AND2 C1732 ( .A(N845), .B(m4stg_shl_tmp[149]), .Z(N846) );
  GTECH_AND2 C1733 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N845) );
  GTECH_AND2 C1734 ( .A(N847), .B(m5stg_frac_54_33[36]), .Z(N848) );
  GTECH_NOT I_91 ( .A(m6stg_step), .Z(N847) );
  GTECH_NOT I_92 ( .A(N854), .Z(m5stg_frac_pre1_in[35]) );
  GTECH_OR2 C1737 ( .A(N851), .B(N853), .Z(N854) );
  GTECH_AND2 C1738 ( .A(N850), .B(m4stg_shl_tmp[148]), .Z(N851) );
  GTECH_AND2 C1739 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N850) );
  GTECH_AND2 C1740 ( .A(N852), .B(m5stg_frac_54_33[35]), .Z(N853) );
  GTECH_NOT I_93 ( .A(m6stg_step), .Z(N852) );
  GTECH_NOT I_94 ( .A(N859), .Z(m5stg_frac_pre1_in[34]) );
  GTECH_OR2 C1743 ( .A(N856), .B(N858), .Z(N859) );
  GTECH_AND2 C1744 ( .A(N855), .B(m4stg_shl_tmp[147]), .Z(N856) );
  GTECH_AND2 C1745 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N855) );
  GTECH_AND2 C1746 ( .A(N857), .B(m5stg_frac_54_33[34]), .Z(N858) );
  GTECH_NOT I_95 ( .A(m6stg_step), .Z(N857) );
  GTECH_NOT I_96 ( .A(N864), .Z(m5stg_frac_pre1_in[33]) );
  GTECH_OR2 C1749 ( .A(N861), .B(N863), .Z(N864) );
  GTECH_AND2 C1750 ( .A(N860), .B(m4stg_shl_tmp[146]), .Z(N861) );
  GTECH_AND2 C1751 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N860) );
  GTECH_AND2 C1752 ( .A(N862), .B(m5stg_frac_54_33[33]), .Z(N863) );
  GTECH_NOT I_97 ( .A(m6stg_step), .Z(N862) );
  GTECH_NOT I_98 ( .A(N869), .Z(m5stg_frac_pre1_in[32]) );
  GTECH_OR2 C1755 ( .A(N866), .B(N868), .Z(N869) );
  GTECH_AND2 C1756 ( .A(N865), .B(m4stg_shl_tmp[145]), .Z(N866) );
  GTECH_AND2 C1757 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N865) );
  GTECH_AND2 C1758 ( .A(N867), .B(m5stg_frac_32_0[32]), .Z(N868) );
  GTECH_NOT I_99 ( .A(m6stg_step), .Z(N867) );
  GTECH_NOT I_100 ( .A(N874), .Z(m5stg_frac_pre1_in[31]) );
  GTECH_OR2 C1761 ( .A(N871), .B(N873), .Z(N874) );
  GTECH_AND2 C1762 ( .A(N870), .B(m4stg_shl_tmp[144]), .Z(N871) );
  GTECH_AND2 C1763 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N870) );
  GTECH_AND2 C1764 ( .A(N872), .B(m5stg_frac_32_0[31]), .Z(N873) );
  GTECH_NOT I_101 ( .A(m6stg_step), .Z(N872) );
  GTECH_NOT I_102 ( .A(N879), .Z(m5stg_frac_pre1_in[30]) );
  GTECH_OR2 C1767 ( .A(N876), .B(N878), .Z(N879) );
  GTECH_AND2 C1768 ( .A(N875), .B(m4stg_shl_tmp[143]), .Z(N876) );
  GTECH_AND2 C1769 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N875) );
  GTECH_AND2 C1770 ( .A(N877), .B(m5stg_frac_32_0[30]), .Z(N878) );
  GTECH_NOT I_103 ( .A(m6stg_step), .Z(N877) );
  GTECH_NOT I_104 ( .A(N884), .Z(m5stg_frac_pre1_in[29]) );
  GTECH_OR2 C1773 ( .A(N881), .B(N883), .Z(N884) );
  GTECH_AND2 C1774 ( .A(N880), .B(m4stg_shl_tmp[142]), .Z(N881) );
  GTECH_AND2 C1775 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N880) );
  GTECH_AND2 C1776 ( .A(N882), .B(m5stg_frac_32_0[29]), .Z(N883) );
  GTECH_NOT I_105 ( .A(m6stg_step), .Z(N882) );
  GTECH_NOT I_106 ( .A(N889), .Z(m5stg_frac_pre1_in[28]) );
  GTECH_OR2 C1779 ( .A(N886), .B(N888), .Z(N889) );
  GTECH_AND2 C1780 ( .A(N885), .B(m4stg_shl_tmp[141]), .Z(N886) );
  GTECH_AND2 C1781 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N885) );
  GTECH_AND2 C1782 ( .A(N887), .B(m5stg_frac_32_0[28]), .Z(N888) );
  GTECH_NOT I_107 ( .A(m6stg_step), .Z(N887) );
  GTECH_NOT I_108 ( .A(N894), .Z(m5stg_frac_pre1_in[27]) );
  GTECH_OR2 C1785 ( .A(N891), .B(N893), .Z(N894) );
  GTECH_AND2 C1786 ( .A(N890), .B(m4stg_shl_tmp[140]), .Z(N891) );
  GTECH_AND2 C1787 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N890) );
  GTECH_AND2 C1788 ( .A(N892), .B(m5stg_frac_32_0[27]), .Z(N893) );
  GTECH_NOT I_109 ( .A(m6stg_step), .Z(N892) );
  GTECH_NOT I_110 ( .A(N899), .Z(m5stg_frac_pre1_in[26]) );
  GTECH_OR2 C1791 ( .A(N896), .B(N898), .Z(N899) );
  GTECH_AND2 C1792 ( .A(N895), .B(m4stg_shl_tmp[139]), .Z(N896) );
  GTECH_AND2 C1793 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N895) );
  GTECH_AND2 C1794 ( .A(N897), .B(m5stg_frac_32_0[26]), .Z(N898) );
  GTECH_NOT I_111 ( .A(m6stg_step), .Z(N897) );
  GTECH_NOT I_112 ( .A(N904), .Z(m5stg_frac_pre1_in[25]) );
  GTECH_OR2 C1797 ( .A(N901), .B(N903), .Z(N904) );
  GTECH_AND2 C1798 ( .A(N900), .B(m4stg_shl_tmp[138]), .Z(N901) );
  GTECH_AND2 C1799 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N900) );
  GTECH_AND2 C1800 ( .A(N902), .B(m5stg_frac_32_0[25]), .Z(N903) );
  GTECH_NOT I_113 ( .A(m6stg_step), .Z(N902) );
  GTECH_NOT I_114 ( .A(N909), .Z(m5stg_frac_pre1_in[24]) );
  GTECH_OR2 C1803 ( .A(N906), .B(N908), .Z(N909) );
  GTECH_AND2 C1804 ( .A(N905), .B(m4stg_shl_tmp[137]), .Z(N906) );
  GTECH_AND2 C1805 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N905) );
  GTECH_AND2 C1806 ( .A(N907), .B(m5stg_frac_32_0[24]), .Z(N908) );
  GTECH_NOT I_115 ( .A(m6stg_step), .Z(N907) );
  GTECH_NOT I_116 ( .A(N914), .Z(m5stg_frac_pre1_in[23]) );
  GTECH_OR2 C1809 ( .A(N911), .B(N913), .Z(N914) );
  GTECH_AND2 C1810 ( .A(N910), .B(m4stg_shl_tmp[136]), .Z(N911) );
  GTECH_AND2 C1811 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N910) );
  GTECH_AND2 C1812 ( .A(N912), .B(m5stg_frac_32_0[23]), .Z(N913) );
  GTECH_NOT I_117 ( .A(m6stg_step), .Z(N912) );
  GTECH_NOT I_118 ( .A(N919), .Z(m5stg_frac_pre1_in[22]) );
  GTECH_OR2 C1815 ( .A(N916), .B(N918), .Z(N919) );
  GTECH_AND2 C1816 ( .A(N915), .B(m4stg_shl_tmp[135]), .Z(N916) );
  GTECH_AND2 C1817 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N915) );
  GTECH_AND2 C1818 ( .A(N917), .B(m5stg_frac_32_0[22]), .Z(N918) );
  GTECH_NOT I_119 ( .A(m6stg_step), .Z(N917) );
  GTECH_NOT I_120 ( .A(N924), .Z(m5stg_frac_pre1_in[21]) );
  GTECH_OR2 C1821 ( .A(N921), .B(N923), .Z(N924) );
  GTECH_AND2 C1822 ( .A(N920), .B(m4stg_shl_tmp[134]), .Z(N921) );
  GTECH_AND2 C1823 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N920) );
  GTECH_AND2 C1824 ( .A(N922), .B(m5stg_frac_32_0[21]), .Z(N923) );
  GTECH_NOT I_121 ( .A(m6stg_step), .Z(N922) );
  GTECH_NOT I_122 ( .A(N929), .Z(m5stg_frac_pre1_in[20]) );
  GTECH_OR2 C1827 ( .A(N926), .B(N928), .Z(N929) );
  GTECH_AND2 C1828 ( .A(N925), .B(m4stg_shl_tmp[133]), .Z(N926) );
  GTECH_AND2 C1829 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N925) );
  GTECH_AND2 C1830 ( .A(N927), .B(m5stg_frac_32_0[20]), .Z(N928) );
  GTECH_NOT I_123 ( .A(m6stg_step), .Z(N927) );
  GTECH_NOT I_124 ( .A(N934), .Z(m5stg_frac_pre1_in[19]) );
  GTECH_OR2 C1833 ( .A(N931), .B(N933), .Z(N934) );
  GTECH_AND2 C1834 ( .A(N930), .B(m4stg_shl_tmp[132]), .Z(N931) );
  GTECH_AND2 C1835 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N930) );
  GTECH_AND2 C1836 ( .A(N932), .B(m5stg_frac_32_0[19]), .Z(N933) );
  GTECH_NOT I_125 ( .A(m6stg_step), .Z(N932) );
  GTECH_NOT I_126 ( .A(N939), .Z(m5stg_frac_pre1_in[18]) );
  GTECH_OR2 C1839 ( .A(N936), .B(N938), .Z(N939) );
  GTECH_AND2 C1840 ( .A(N935), .B(m4stg_shl_tmp[131]), .Z(N936) );
  GTECH_AND2 C1841 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N935) );
  GTECH_AND2 C1842 ( .A(N937), .B(m5stg_frac_32_0[18]), .Z(N938) );
  GTECH_NOT I_127 ( .A(m6stg_step), .Z(N937) );
  GTECH_NOT I_128 ( .A(N944), .Z(m5stg_frac_pre1_in[17]) );
  GTECH_OR2 C1845 ( .A(N941), .B(N943), .Z(N944) );
  GTECH_AND2 C1846 ( .A(N940), .B(m4stg_shl_tmp[130]), .Z(N941) );
  GTECH_AND2 C1847 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N940) );
  GTECH_AND2 C1848 ( .A(N942), .B(m5stg_frac_32_0[17]), .Z(N943) );
  GTECH_NOT I_129 ( .A(m6stg_step), .Z(N942) );
  GTECH_NOT I_130 ( .A(N949), .Z(m5stg_frac_pre1_in[16]) );
  GTECH_OR2 C1851 ( .A(N946), .B(N948), .Z(N949) );
  GTECH_AND2 C1852 ( .A(N945), .B(m4stg_shl_tmp[129]), .Z(N946) );
  GTECH_AND2 C1853 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N945) );
  GTECH_AND2 C1854 ( .A(N947), .B(m5stg_frac_32_0[16]), .Z(N948) );
  GTECH_NOT I_131 ( .A(m6stg_step), .Z(N947) );
  GTECH_NOT I_132 ( .A(N954), .Z(m5stg_frac_pre1_in[15]) );
  GTECH_OR2 C1857 ( .A(N951), .B(N953), .Z(N954) );
  GTECH_AND2 C1858 ( .A(N950), .B(m4stg_shl_tmp[128]), .Z(N951) );
  GTECH_AND2 C1859 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N950) );
  GTECH_AND2 C1860 ( .A(N952), .B(m5stg_frac_32_0[15]), .Z(N953) );
  GTECH_NOT I_133 ( .A(m6stg_step), .Z(N952) );
  GTECH_NOT I_134 ( .A(N959), .Z(m5stg_frac_pre1_in[14]) );
  GTECH_OR2 C1863 ( .A(N956), .B(N958), .Z(N959) );
  GTECH_AND2 C1864 ( .A(N955), .B(m4stg_shl_tmp[127]), .Z(N956) );
  GTECH_AND2 C1865 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N955) );
  GTECH_AND2 C1866 ( .A(N957), .B(m5stg_frac_32_0[14]), .Z(N958) );
  GTECH_NOT I_135 ( .A(m6stg_step), .Z(N957) );
  GTECH_NOT I_136 ( .A(N964), .Z(m5stg_frac_pre1_in[13]) );
  GTECH_OR2 C1869 ( .A(N961), .B(N963), .Z(N964) );
  GTECH_AND2 C1870 ( .A(N960), .B(m4stg_shl_tmp[126]), .Z(N961) );
  GTECH_AND2 C1871 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N960) );
  GTECH_AND2 C1872 ( .A(N962), .B(m5stg_frac_32_0[13]), .Z(N963) );
  GTECH_NOT I_137 ( .A(m6stg_step), .Z(N962) );
  GTECH_NOT I_138 ( .A(N969), .Z(m5stg_frac_pre1_in[12]) );
  GTECH_OR2 C1875 ( .A(N966), .B(N968), .Z(N969) );
  GTECH_AND2 C1876 ( .A(N965), .B(m4stg_shl_tmp[125]), .Z(N966) );
  GTECH_AND2 C1877 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N965) );
  GTECH_AND2 C1878 ( .A(N967), .B(m5stg_frac_32_0[12]), .Z(N968) );
  GTECH_NOT I_139 ( .A(m6stg_step), .Z(N967) );
  GTECH_NOT I_140 ( .A(N974), .Z(m5stg_frac_pre1_in[11]) );
  GTECH_OR2 C1881 ( .A(N971), .B(N973), .Z(N974) );
  GTECH_AND2 C1882 ( .A(N970), .B(m4stg_shl_tmp[124]), .Z(N971) );
  GTECH_AND2 C1883 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N970) );
  GTECH_AND2 C1884 ( .A(N972), .B(m5stg_frac_32_0[11]), .Z(N973) );
  GTECH_NOT I_141 ( .A(m6stg_step), .Z(N972) );
  GTECH_NOT I_142 ( .A(N979), .Z(m5stg_frac_pre1_in[10]) );
  GTECH_OR2 C1887 ( .A(N976), .B(N978), .Z(N979) );
  GTECH_AND2 C1888 ( .A(N975), .B(m4stg_shl_tmp[123]), .Z(N976) );
  GTECH_AND2 C1889 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N975) );
  GTECH_AND2 C1890 ( .A(N977), .B(m5stg_frac_32_0[10]), .Z(N978) );
  GTECH_NOT I_143 ( .A(m6stg_step), .Z(N977) );
  GTECH_NOT I_144 ( .A(N984), .Z(m5stg_frac_pre1_in[9]) );
  GTECH_OR2 C1893 ( .A(N981), .B(N983), .Z(N984) );
  GTECH_AND2 C1894 ( .A(N980), .B(m4stg_shl_tmp[122]), .Z(N981) );
  GTECH_AND2 C1895 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N980) );
  GTECH_AND2 C1896 ( .A(N982), .B(m5stg_frac_32_0[9]), .Z(N983) );
  GTECH_NOT I_145 ( .A(m6stg_step), .Z(N982) );
  GTECH_NOT I_146 ( .A(N989), .Z(m5stg_frac_pre1_in[8]) );
  GTECH_OR2 C1899 ( .A(N986), .B(N988), .Z(N989) );
  GTECH_AND2 C1900 ( .A(N985), .B(m4stg_shl_tmp[121]), .Z(N986) );
  GTECH_AND2 C1901 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N985) );
  GTECH_AND2 C1902 ( .A(N987), .B(m5stg_frac_32_0[8]), .Z(N988) );
  GTECH_NOT I_147 ( .A(m6stg_step), .Z(N987) );
  GTECH_NOT I_148 ( .A(N994), .Z(m5stg_frac_pre1_in[7]) );
  GTECH_OR2 C1905 ( .A(N991), .B(N993), .Z(N994) );
  GTECH_AND2 C1906 ( .A(N990), .B(m4stg_shl_tmp[120]), .Z(N991) );
  GTECH_AND2 C1907 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N990) );
  GTECH_AND2 C1908 ( .A(N992), .B(m5stg_frac_32_0[7]), .Z(N993) );
  GTECH_NOT I_149 ( .A(m6stg_step), .Z(N992) );
  GTECH_NOT I_150 ( .A(N999), .Z(m5stg_frac_pre1_in[6]) );
  GTECH_OR2 C1911 ( .A(N996), .B(N998), .Z(N999) );
  GTECH_AND2 C1912 ( .A(N995), .B(m4stg_shl_tmp[119]), .Z(N996) );
  GTECH_AND2 C1913 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N995) );
  GTECH_AND2 C1914 ( .A(N997), .B(m5stg_frac_32_0[6]), .Z(N998) );
  GTECH_NOT I_151 ( .A(m6stg_step), .Z(N997) );
  GTECH_NOT I_152 ( .A(N1004), .Z(m5stg_frac_pre1_in[5]) );
  GTECH_OR2 C1917 ( .A(N1001), .B(N1003), .Z(N1004) );
  GTECH_AND2 C1918 ( .A(N1000), .B(m4stg_shl_tmp[118]), .Z(N1001) );
  GTECH_AND2 C1919 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1000) );
  GTECH_AND2 C1920 ( .A(N1002), .B(m5stg_frac_32_0[5]), .Z(N1003) );
  GTECH_NOT I_153 ( .A(m6stg_step), .Z(N1002) );
  GTECH_NOT I_154 ( .A(N1009), .Z(m5stg_frac_pre1_in[4]) );
  GTECH_OR2 C1923 ( .A(N1006), .B(N1008), .Z(N1009) );
  GTECH_AND2 C1924 ( .A(N1005), .B(m4stg_shl_tmp[117]), .Z(N1006) );
  GTECH_AND2 C1925 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1005) );
  GTECH_AND2 C1926 ( .A(N1007), .B(m5stg_frac_32_0[4]), .Z(N1008) );
  GTECH_NOT I_155 ( .A(m6stg_step), .Z(N1007) );
  GTECH_NOT I_156 ( .A(N1014), .Z(m5stg_frac_pre1_in[3]) );
  GTECH_OR2 C1929 ( .A(N1011), .B(N1013), .Z(N1014) );
  GTECH_AND2 C1930 ( .A(N1010), .B(m4stg_shl_tmp[116]), .Z(N1011) );
  GTECH_AND2 C1931 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1010) );
  GTECH_AND2 C1932 ( .A(N1012), .B(m5stg_frac_32_0[3]), .Z(N1013) );
  GTECH_NOT I_157 ( .A(m6stg_step), .Z(N1012) );
  GTECH_NOT I_158 ( .A(N1019), .Z(m5stg_frac_pre1_in[2]) );
  GTECH_OR2 C1935 ( .A(N1016), .B(N1018), .Z(N1019) );
  GTECH_AND2 C1936 ( .A(N1015), .B(m4stg_shl_tmp[115]), .Z(N1016) );
  GTECH_AND2 C1937 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1015) );
  GTECH_AND2 C1938 ( .A(N1017), .B(m5stg_frac_32_0[2]), .Z(N1018) );
  GTECH_NOT I_159 ( .A(m6stg_step), .Z(N1017) );
  GTECH_NOT I_160 ( .A(N1024), .Z(m5stg_frac_pre1_in[1]) );
  GTECH_OR2 C1941 ( .A(N1021), .B(N1023), .Z(N1024) );
  GTECH_AND2 C1942 ( .A(N1020), .B(m4stg_shl_tmp[114]), .Z(N1021) );
  GTECH_AND2 C1943 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1020) );
  GTECH_AND2 C1944 ( .A(N1022), .B(m5stg_frac_32_0[1]), .Z(N1023) );
  GTECH_NOT I_161 ( .A(m6stg_step), .Z(N1022) );
  GTECH_NOT I_162 ( .A(N1029), .Z(m5stg_frac_pre1_in[0]) );
  GTECH_OR2 C1947 ( .A(N1026), .B(N1028), .Z(N1029) );
  GTECH_AND2 C1948 ( .A(N1025), .B(m4stg_shl[0]), .Z(N1026) );
  GTECH_AND2 C1949 ( .A(m4stg_left_shift_step), .B(m4stg_shl_55), .Z(N1025) );
  GTECH_AND2 C1950 ( .A(N1027), .B(m5stg_frac_32_0[0]), .Z(N1028) );
  GTECH_NOT I_163 ( .A(m6stg_step), .Z(N1027) );
  GTECH_NOT I_164 ( .A(N1032), .Z(m5stg_frac_pre2_in[54]) );
  GTECH_AND2 C1953 ( .A(N1031), .B(m4stg_shl_tmp[166]), .Z(N1032) );
  GTECH_AND2 C1954 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1031) );
  GTECH_NOT I_165 ( .A(m4stg_shl_55), .Z(N1030) );
  GTECH_NOT I_166 ( .A(N1034), .Z(m5stg_frac_pre2_in[53]) );
  GTECH_AND2 C1957 ( .A(N1033), .B(m4stg_shl_tmp[165]), .Z(N1034) );
  GTECH_AND2 C1958 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1033) );
  GTECH_NOT I_167 ( .A(N1036), .Z(m5stg_frac_pre2_in[52]) );
  GTECH_AND2 C1961 ( .A(N1035), .B(m4stg_shl_tmp[164]), .Z(N1036) );
  GTECH_AND2 C1962 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1035) );
  GTECH_NOT I_168 ( .A(N1038), .Z(m5stg_frac_pre2_in[51]) );
  GTECH_AND2 C1965 ( .A(N1037), .B(m4stg_shl_tmp[163]), .Z(N1038) );
  GTECH_AND2 C1966 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1037) );
  GTECH_NOT I_169 ( .A(N1040), .Z(m5stg_frac_pre2_in[50]) );
  GTECH_AND2 C1969 ( .A(N1039), .B(m4stg_shl_tmp[162]), .Z(N1040) );
  GTECH_AND2 C1970 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1039) );
  GTECH_NOT I_170 ( .A(N1042), .Z(m5stg_frac_pre2_in[49]) );
  GTECH_AND2 C1973 ( .A(N1041), .B(m4stg_shl_tmp[161]), .Z(N1042) );
  GTECH_AND2 C1974 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1041) );
  GTECH_NOT I_171 ( .A(N1044), .Z(m5stg_frac_pre2_in[48]) );
  GTECH_AND2 C1977 ( .A(N1043), .B(m4stg_shl_tmp[160]), .Z(N1044) );
  GTECH_AND2 C1978 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1043) );
  GTECH_NOT I_172 ( .A(N1046), .Z(m5stg_frac_pre2_in[47]) );
  GTECH_AND2 C1981 ( .A(N1045), .B(m4stg_shl_tmp[159]), .Z(N1046) );
  GTECH_AND2 C1982 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1045) );
  GTECH_NOT I_173 ( .A(N1048), .Z(m5stg_frac_pre2_in[46]) );
  GTECH_AND2 C1985 ( .A(N1047), .B(m4stg_shl_tmp[158]), .Z(N1048) );
  GTECH_AND2 C1986 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1047) );
  GTECH_NOT I_174 ( .A(N1050), .Z(m5stg_frac_pre2_in[45]) );
  GTECH_AND2 C1989 ( .A(N1049), .B(m4stg_shl_tmp[157]), .Z(N1050) );
  GTECH_AND2 C1990 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1049) );
  GTECH_NOT I_175 ( .A(N1052), .Z(m5stg_frac_pre2_in[44]) );
  GTECH_AND2 C1993 ( .A(N1051), .B(m4stg_shl_tmp[156]), .Z(N1052) );
  GTECH_AND2 C1994 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1051) );
  GTECH_NOT I_176 ( .A(N1054), .Z(m5stg_frac_pre2_in[43]) );
  GTECH_AND2 C1997 ( .A(N1053), .B(m4stg_shl_tmp[155]), .Z(N1054) );
  GTECH_AND2 C1998 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1053) );
  GTECH_NOT I_177 ( .A(N1056), .Z(m5stg_frac_pre2_in[42]) );
  GTECH_AND2 C2001 ( .A(N1055), .B(m4stg_shl_tmp[154]), .Z(N1056) );
  GTECH_AND2 C2002 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1055) );
  GTECH_NOT I_178 ( .A(N1058), .Z(m5stg_frac_pre2_in[41]) );
  GTECH_AND2 C2005 ( .A(N1057), .B(m4stg_shl_tmp[153]), .Z(N1058) );
  GTECH_AND2 C2006 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1057) );
  GTECH_NOT I_179 ( .A(N1060), .Z(m5stg_frac_pre2_in[40]) );
  GTECH_AND2 C2009 ( .A(N1059), .B(m4stg_shl_tmp[152]), .Z(N1060) );
  GTECH_AND2 C2010 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1059) );
  GTECH_NOT I_180 ( .A(N1062), .Z(m5stg_frac_pre2_in[39]) );
  GTECH_AND2 C2013 ( .A(N1061), .B(m4stg_shl_tmp[151]), .Z(N1062) );
  GTECH_AND2 C2014 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1061) );
  GTECH_NOT I_181 ( .A(N1064), .Z(m5stg_frac_pre2_in[38]) );
  GTECH_AND2 C2017 ( .A(N1063), .B(m4stg_shl_tmp[150]), .Z(N1064) );
  GTECH_AND2 C2018 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1063) );
  GTECH_NOT I_182 ( .A(N1066), .Z(m5stg_frac_pre2_in[37]) );
  GTECH_AND2 C2021 ( .A(N1065), .B(m4stg_shl_tmp[149]), .Z(N1066) );
  GTECH_AND2 C2022 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1065) );
  GTECH_NOT I_183 ( .A(N1068), .Z(m5stg_frac_pre2_in[36]) );
  GTECH_AND2 C2025 ( .A(N1067), .B(m4stg_shl_tmp[148]), .Z(N1068) );
  GTECH_AND2 C2026 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1067) );
  GTECH_NOT I_184 ( .A(N1070), .Z(m5stg_frac_pre2_in[35]) );
  GTECH_AND2 C2029 ( .A(N1069), .B(m4stg_shl_tmp[147]), .Z(N1070) );
  GTECH_AND2 C2030 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1069) );
  GTECH_NOT I_185 ( .A(N1072), .Z(m5stg_frac_pre2_in[34]) );
  GTECH_AND2 C2033 ( .A(N1071), .B(m4stg_shl_tmp[146]), .Z(N1072) );
  GTECH_AND2 C2034 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1071) );
  GTECH_NOT I_186 ( .A(N1074), .Z(m5stg_frac_pre2_in[33]) );
  GTECH_AND2 C2037 ( .A(N1073), .B(m4stg_shl_tmp[145]), .Z(N1074) );
  GTECH_AND2 C2038 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1073) );
  GTECH_NOT I_187 ( .A(N1076), .Z(m5stg_frac_pre2_in[32]) );
  GTECH_AND2 C2041 ( .A(N1075), .B(m4stg_shl_tmp[144]), .Z(N1076) );
  GTECH_AND2 C2042 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1075) );
  GTECH_NOT I_188 ( .A(N1078), .Z(m5stg_frac_pre2_in[31]) );
  GTECH_AND2 C2045 ( .A(N1077), .B(m4stg_shl_tmp[143]), .Z(N1078) );
  GTECH_AND2 C2046 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1077) );
  GTECH_NOT I_189 ( .A(N1080), .Z(m5stg_frac_pre2_in[30]) );
  GTECH_AND2 C2049 ( .A(N1079), .B(m4stg_shl_tmp[142]), .Z(N1080) );
  GTECH_AND2 C2050 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1079) );
  GTECH_NOT I_190 ( .A(N1082), .Z(m5stg_frac_pre2_in[29]) );
  GTECH_AND2 C2053 ( .A(N1081), .B(m4stg_shl_tmp[141]), .Z(N1082) );
  GTECH_AND2 C2054 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1081) );
  GTECH_NOT I_191 ( .A(N1084), .Z(m5stg_frac_pre2_in[28]) );
  GTECH_AND2 C2057 ( .A(N1083), .B(m4stg_shl_tmp[140]), .Z(N1084) );
  GTECH_AND2 C2058 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1083) );
  GTECH_NOT I_192 ( .A(N1086), .Z(m5stg_frac_pre2_in[27]) );
  GTECH_AND2 C2061 ( .A(N1085), .B(m4stg_shl_tmp[139]), .Z(N1086) );
  GTECH_AND2 C2062 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1085) );
  GTECH_NOT I_193 ( .A(N1088), .Z(m5stg_frac_pre2_in[26]) );
  GTECH_AND2 C2065 ( .A(N1087), .B(m4stg_shl_tmp[138]), .Z(N1088) );
  GTECH_AND2 C2066 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1087) );
  GTECH_NOT I_194 ( .A(N1090), .Z(m5stg_frac_pre2_in[25]) );
  GTECH_AND2 C2069 ( .A(N1089), .B(m4stg_shl_tmp[137]), .Z(N1090) );
  GTECH_AND2 C2070 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1089) );
  GTECH_NOT I_195 ( .A(N1092), .Z(m5stg_frac_pre2_in[24]) );
  GTECH_AND2 C2073 ( .A(N1091), .B(m4stg_shl_tmp[136]), .Z(N1092) );
  GTECH_AND2 C2074 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1091) );
  GTECH_NOT I_196 ( .A(N1094), .Z(m5stg_frac_pre2_in[23]) );
  GTECH_AND2 C2077 ( .A(N1093), .B(m4stg_shl_tmp[135]), .Z(N1094) );
  GTECH_AND2 C2078 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1093) );
  GTECH_NOT I_197 ( .A(N1096), .Z(m5stg_frac_pre2_in[22]) );
  GTECH_AND2 C2081 ( .A(N1095), .B(m4stg_shl_tmp[134]), .Z(N1096) );
  GTECH_AND2 C2082 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1095) );
  GTECH_NOT I_198 ( .A(N1098), .Z(m5stg_frac_pre2_in[21]) );
  GTECH_AND2 C2085 ( .A(N1097), .B(m4stg_shl_tmp[133]), .Z(N1098) );
  GTECH_AND2 C2086 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1097) );
  GTECH_NOT I_199 ( .A(N1100), .Z(m5stg_frac_pre2_in[20]) );
  GTECH_AND2 C2089 ( .A(N1099), .B(m4stg_shl_tmp[132]), .Z(N1100) );
  GTECH_AND2 C2090 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1099) );
  GTECH_NOT I_200 ( .A(N1102), .Z(m5stg_frac_pre2_in[19]) );
  GTECH_AND2 C2093 ( .A(N1101), .B(m4stg_shl_tmp[131]), .Z(N1102) );
  GTECH_AND2 C2094 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1101) );
  GTECH_NOT I_201 ( .A(N1104), .Z(m5stg_frac_pre2_in[18]) );
  GTECH_AND2 C2097 ( .A(N1103), .B(m4stg_shl_tmp[130]), .Z(N1104) );
  GTECH_AND2 C2098 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1103) );
  GTECH_NOT I_202 ( .A(N1106), .Z(m5stg_frac_pre2_in[17]) );
  GTECH_AND2 C2101 ( .A(N1105), .B(m4stg_shl_tmp[129]), .Z(N1106) );
  GTECH_AND2 C2102 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1105) );
  GTECH_NOT I_203 ( .A(N1108), .Z(m5stg_frac_pre2_in[16]) );
  GTECH_AND2 C2105 ( .A(N1107), .B(m4stg_shl_tmp[128]), .Z(N1108) );
  GTECH_AND2 C2106 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1107) );
  GTECH_NOT I_204 ( .A(N1110), .Z(m5stg_frac_pre2_in[15]) );
  GTECH_AND2 C2109 ( .A(N1109), .B(m4stg_shl_tmp[127]), .Z(N1110) );
  GTECH_AND2 C2110 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1109) );
  GTECH_NOT I_205 ( .A(N1112), .Z(m5stg_frac_pre2_in[14]) );
  GTECH_AND2 C2113 ( .A(N1111), .B(m4stg_shl_tmp[126]), .Z(N1112) );
  GTECH_AND2 C2114 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1111) );
  GTECH_NOT I_206 ( .A(N1114), .Z(m5stg_frac_pre2_in[13]) );
  GTECH_AND2 C2117 ( .A(N1113), .B(m4stg_shl_tmp[125]), .Z(N1114) );
  GTECH_AND2 C2118 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1113) );
  GTECH_NOT I_207 ( .A(N1116), .Z(m5stg_frac_pre2_in[12]) );
  GTECH_AND2 C2121 ( .A(N1115), .B(m4stg_shl_tmp[124]), .Z(N1116) );
  GTECH_AND2 C2122 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1115) );
  GTECH_NOT I_208 ( .A(N1118), .Z(m5stg_frac_pre2_in[11]) );
  GTECH_AND2 C2125 ( .A(N1117), .B(m4stg_shl_tmp[123]), .Z(N1118) );
  GTECH_AND2 C2126 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1117) );
  GTECH_NOT I_209 ( .A(N1120), .Z(m5stg_frac_pre2_in[10]) );
  GTECH_AND2 C2129 ( .A(N1119), .B(m4stg_shl_tmp[122]), .Z(N1120) );
  GTECH_AND2 C2130 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1119) );
  GTECH_NOT I_210 ( .A(N1122), .Z(m5stg_frac_pre2_in[9]) );
  GTECH_AND2 C2133 ( .A(N1121), .B(m4stg_shl_tmp[121]), .Z(N1122) );
  GTECH_AND2 C2134 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1121) );
  GTECH_NOT I_211 ( .A(N1124), .Z(m5stg_frac_pre2_in[8]) );
  GTECH_AND2 C2137 ( .A(N1123), .B(m4stg_shl_tmp[120]), .Z(N1124) );
  GTECH_AND2 C2138 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1123) );
  GTECH_NOT I_212 ( .A(N1126), .Z(m5stg_frac_pre2_in[7]) );
  GTECH_AND2 C2141 ( .A(N1125), .B(m4stg_shl_tmp[119]), .Z(N1126) );
  GTECH_AND2 C2142 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1125) );
  GTECH_NOT I_213 ( .A(N1128), .Z(m5stg_frac_pre2_in[6]) );
  GTECH_AND2 C2145 ( .A(N1127), .B(m4stg_shl_tmp[118]), .Z(N1128) );
  GTECH_AND2 C2146 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1127) );
  GTECH_NOT I_214 ( .A(N1130), .Z(m5stg_frac_pre2_in[5]) );
  GTECH_AND2 C2149 ( .A(N1129), .B(m4stg_shl_tmp[117]), .Z(N1130) );
  GTECH_AND2 C2150 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1129) );
  GTECH_NOT I_215 ( .A(N1132), .Z(m5stg_frac_pre2_in[4]) );
  GTECH_AND2 C2153 ( .A(N1131), .B(m4stg_shl_tmp[116]), .Z(N1132) );
  GTECH_AND2 C2154 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1131) );
  GTECH_NOT I_216 ( .A(N1134), .Z(m5stg_frac_pre2_in[3]) );
  GTECH_AND2 C2157 ( .A(N1133), .B(m4stg_shl_tmp[115]), .Z(N1134) );
  GTECH_AND2 C2158 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1133) );
  GTECH_NOT I_217 ( .A(N1136), .Z(m5stg_frac_pre2_in[2]) );
  GTECH_AND2 C2161 ( .A(N1135), .B(m4stg_shl_tmp[114]), .Z(N1136) );
  GTECH_AND2 C2162 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1135) );
  GTECH_NOT I_218 ( .A(N1138), .Z(m5stg_frac_pre2_in[1]) );
  GTECH_AND2 C2165 ( .A(N1137), .B(m4stg_shl[0]), .Z(N1138) );
  GTECH_AND2 C2166 ( .A(m4stg_left_shift_step), .B(N1030), .Z(N1137) );
  GTECH_NOT I_219 ( .A(N1140), .Z(m5stg_frac_pre3_in[54]) );
  GTECH_AND2 C2169 ( .A(N1139), .B(m4stg_shr_tmp[167]), .Z(N1140) );
  GTECH_AND2 C2170 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1139) );
  GTECH_NOT I_220 ( .A(N1142), .Z(m5stg_frac_pre3_in[53]) );
  GTECH_AND2 C2172 ( .A(N1141), .B(m4stg_shr_tmp[166]), .Z(N1142) );
  GTECH_AND2 C2173 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1141) );
  GTECH_NOT I_221 ( .A(N1144), .Z(m5stg_frac_pre3_in[52]) );
  GTECH_AND2 C2175 ( .A(N1143), .B(m4stg_shr_tmp[165]), .Z(N1144) );
  GTECH_AND2 C2176 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1143) );
  GTECH_NOT I_222 ( .A(N1146), .Z(m5stg_frac_pre3_in[51]) );
  GTECH_AND2 C2178 ( .A(N1145), .B(m4stg_shr_tmp[164]), .Z(N1146) );
  GTECH_AND2 C2179 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1145) );
  GTECH_NOT I_223 ( .A(N1148), .Z(m5stg_frac_pre3_in[50]) );
  GTECH_AND2 C2181 ( .A(N1147), .B(m4stg_shr_tmp[163]), .Z(N1148) );
  GTECH_AND2 C2182 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1147) );
  GTECH_NOT I_224 ( .A(N1150), .Z(m5stg_frac_pre3_in[49]) );
  GTECH_AND2 C2184 ( .A(N1149), .B(m4stg_shr_tmp[162]), .Z(N1150) );
  GTECH_AND2 C2185 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1149) );
  GTECH_NOT I_225 ( .A(N1152), .Z(m5stg_frac_pre3_in[48]) );
  GTECH_AND2 C2187 ( .A(N1151), .B(m4stg_shr_tmp[161]), .Z(N1152) );
  GTECH_AND2 C2188 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1151) );
  GTECH_NOT I_226 ( .A(N1154), .Z(m5stg_frac_pre3_in[47]) );
  GTECH_AND2 C2190 ( .A(N1153), .B(m4stg_shr_tmp[160]), .Z(N1154) );
  GTECH_AND2 C2191 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1153) );
  GTECH_NOT I_227 ( .A(N1156), .Z(m5stg_frac_pre3_in[46]) );
  GTECH_AND2 C2193 ( .A(N1155), .B(m4stg_shr_tmp[159]), .Z(N1156) );
  GTECH_AND2 C2194 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1155) );
  GTECH_NOT I_228 ( .A(N1158), .Z(m5stg_frac_pre3_in[45]) );
  GTECH_AND2 C2196 ( .A(N1157), .B(m4stg_shr_tmp[158]), .Z(N1158) );
  GTECH_AND2 C2197 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1157) );
  GTECH_NOT I_229 ( .A(N1160), .Z(m5stg_frac_pre3_in[44]) );
  GTECH_AND2 C2199 ( .A(N1159), .B(m4stg_shr_tmp[157]), .Z(N1160) );
  GTECH_AND2 C2200 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1159) );
  GTECH_NOT I_230 ( .A(N1162), .Z(m5stg_frac_pre3_in[43]) );
  GTECH_AND2 C2202 ( .A(N1161), .B(m4stg_shr_tmp[156]), .Z(N1162) );
  GTECH_AND2 C2203 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1161) );
  GTECH_NOT I_231 ( .A(N1164), .Z(m5stg_frac_pre3_in[42]) );
  GTECH_AND2 C2205 ( .A(N1163), .B(m4stg_shr_tmp[155]), .Z(N1164) );
  GTECH_AND2 C2206 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1163) );
  GTECH_NOT I_232 ( .A(N1166), .Z(m5stg_frac_pre3_in[41]) );
  GTECH_AND2 C2208 ( .A(N1165), .B(m4stg_shr_tmp[154]), .Z(N1166) );
  GTECH_AND2 C2209 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1165) );
  GTECH_NOT I_233 ( .A(N1168), .Z(m5stg_frac_pre3_in[40]) );
  GTECH_AND2 C2211 ( .A(N1167), .B(m4stg_shr_tmp[153]), .Z(N1168) );
  GTECH_AND2 C2212 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1167) );
  GTECH_NOT I_234 ( .A(N1170), .Z(m5stg_frac_pre3_in[39]) );
  GTECH_AND2 C2214 ( .A(N1169), .B(m4stg_shr_tmp[152]), .Z(N1170) );
  GTECH_AND2 C2215 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1169) );
  GTECH_NOT I_235 ( .A(N1172), .Z(m5stg_frac_pre3_in[38]) );
  GTECH_AND2 C2217 ( .A(N1171), .B(m4stg_shr_tmp[151]), .Z(N1172) );
  GTECH_AND2 C2218 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1171) );
  GTECH_NOT I_236 ( .A(N1174), .Z(m5stg_frac_pre3_in[37]) );
  GTECH_AND2 C2220 ( .A(N1173), .B(m4stg_shr_tmp[150]), .Z(N1174) );
  GTECH_AND2 C2221 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1173) );
  GTECH_NOT I_237 ( .A(N1176), .Z(m5stg_frac_pre3_in[36]) );
  GTECH_AND2 C2223 ( .A(N1175), .B(m4stg_shr_tmp[149]), .Z(N1176) );
  GTECH_AND2 C2224 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1175) );
  GTECH_NOT I_238 ( .A(N1178), .Z(m5stg_frac_pre3_in[35]) );
  GTECH_AND2 C2226 ( .A(N1177), .B(m4stg_shr_tmp[148]), .Z(N1178) );
  GTECH_AND2 C2227 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1177) );
  GTECH_NOT I_239 ( .A(N1180), .Z(m5stg_frac_pre3_in[34]) );
  GTECH_AND2 C2229 ( .A(N1179), .B(m4stg_shr_tmp[147]), .Z(N1180) );
  GTECH_AND2 C2230 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1179) );
  GTECH_NOT I_240 ( .A(N1182), .Z(m5stg_frac_pre3_in[33]) );
  GTECH_AND2 C2232 ( .A(N1181), .B(m4stg_shr_tmp[146]), .Z(N1182) );
  GTECH_AND2 C2233 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1181) );
  GTECH_NOT I_241 ( .A(N1184), .Z(m5stg_frac_pre3_in[32]) );
  GTECH_AND2 C2235 ( .A(N1183), .B(m4stg_shr_tmp[145]), .Z(N1184) );
  GTECH_AND2 C2236 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1183) );
  GTECH_NOT I_242 ( .A(N1186), .Z(m5stg_frac_pre3_in[31]) );
  GTECH_AND2 C2238 ( .A(N1185), .B(m4stg_shr_tmp[144]), .Z(N1186) );
  GTECH_AND2 C2239 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1185) );
  GTECH_NOT I_243 ( .A(N1188), .Z(m5stg_frac_pre3_in[30]) );
  GTECH_AND2 C2241 ( .A(N1187), .B(m4stg_shr_tmp[143]), .Z(N1188) );
  GTECH_AND2 C2242 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1187) );
  GTECH_NOT I_244 ( .A(N1190), .Z(m5stg_frac_pre3_in[29]) );
  GTECH_AND2 C2244 ( .A(N1189), .B(m4stg_shr_tmp[142]), .Z(N1190) );
  GTECH_AND2 C2245 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1189) );
  GTECH_NOT I_245 ( .A(N1192), .Z(m5stg_frac_pre3_in[28]) );
  GTECH_AND2 C2247 ( .A(N1191), .B(m4stg_shr_tmp[141]), .Z(N1192) );
  GTECH_AND2 C2248 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1191) );
  GTECH_NOT I_246 ( .A(N1194), .Z(m5stg_frac_pre3_in[27]) );
  GTECH_AND2 C2250 ( .A(N1193), .B(m4stg_shr_tmp[140]), .Z(N1194) );
  GTECH_AND2 C2251 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1193) );
  GTECH_NOT I_247 ( .A(N1196), .Z(m5stg_frac_pre3_in[26]) );
  GTECH_AND2 C2253 ( .A(N1195), .B(m4stg_shr_tmp[139]), .Z(N1196) );
  GTECH_AND2 C2254 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1195) );
  GTECH_NOT I_248 ( .A(N1198), .Z(m5stg_frac_pre3_in[25]) );
  GTECH_AND2 C2256 ( .A(N1197), .B(m4stg_shr_tmp[138]), .Z(N1198) );
  GTECH_AND2 C2257 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1197) );
  GTECH_NOT I_249 ( .A(N1200), .Z(m5stg_frac_pre3_in[24]) );
  GTECH_AND2 C2259 ( .A(N1199), .B(m4stg_shr_tmp[137]), .Z(N1200) );
  GTECH_AND2 C2260 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1199) );
  GTECH_NOT I_250 ( .A(N1202), .Z(m5stg_frac_pre3_in[23]) );
  GTECH_AND2 C2262 ( .A(N1201), .B(m4stg_shr_tmp[136]), .Z(N1202) );
  GTECH_AND2 C2263 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1201) );
  GTECH_NOT I_251 ( .A(N1204), .Z(m5stg_frac_pre3_in[22]) );
  GTECH_AND2 C2265 ( .A(N1203), .B(m4stg_shr_tmp[135]), .Z(N1204) );
  GTECH_AND2 C2266 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1203) );
  GTECH_NOT I_252 ( .A(N1206), .Z(m5stg_frac_pre3_in[21]) );
  GTECH_AND2 C2268 ( .A(N1205), .B(m4stg_shr_tmp[134]), .Z(N1206) );
  GTECH_AND2 C2269 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1205) );
  GTECH_NOT I_253 ( .A(N1208), .Z(m5stg_frac_pre3_in[20]) );
  GTECH_AND2 C2271 ( .A(N1207), .B(m4stg_shr_tmp[133]), .Z(N1208) );
  GTECH_AND2 C2272 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1207) );
  GTECH_NOT I_254 ( .A(N1210), .Z(m5stg_frac_pre3_in[19]) );
  GTECH_AND2 C2274 ( .A(N1209), .B(m4stg_shr_tmp[132]), .Z(N1210) );
  GTECH_AND2 C2275 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1209) );
  GTECH_NOT I_255 ( .A(N1212), .Z(m5stg_frac_pre3_in[18]) );
  GTECH_AND2 C2277 ( .A(N1211), .B(m4stg_shr_tmp[131]), .Z(N1212) );
  GTECH_AND2 C2278 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1211) );
  GTECH_NOT I_256 ( .A(N1214), .Z(m5stg_frac_pre3_in[17]) );
  GTECH_AND2 C2280 ( .A(N1213), .B(m4stg_shr_tmp[130]), .Z(N1214) );
  GTECH_AND2 C2281 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1213) );
  GTECH_NOT I_257 ( .A(N1216), .Z(m5stg_frac_pre3_in[16]) );
  GTECH_AND2 C2283 ( .A(N1215), .B(m4stg_shr_tmp[129]), .Z(N1216) );
  GTECH_AND2 C2284 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1215) );
  GTECH_NOT I_258 ( .A(N1218), .Z(m5stg_frac_pre3_in[15]) );
  GTECH_AND2 C2286 ( .A(N1217), .B(m4stg_shr_tmp[128]), .Z(N1218) );
  GTECH_AND2 C2287 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1217) );
  GTECH_NOT I_259 ( .A(N1220), .Z(m5stg_frac_pre3_in[14]) );
  GTECH_AND2 C2289 ( .A(N1219), .B(m4stg_shr_tmp[127]), .Z(N1220) );
  GTECH_AND2 C2290 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1219) );
  GTECH_NOT I_260 ( .A(N1222), .Z(m5stg_frac_pre3_in[13]) );
  GTECH_AND2 C2292 ( .A(N1221), .B(m4stg_shr_tmp[126]), .Z(N1222) );
  GTECH_AND2 C2293 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1221) );
  GTECH_NOT I_261 ( .A(N1224), .Z(m5stg_frac_pre3_in[12]) );
  GTECH_AND2 C2295 ( .A(N1223), .B(m4stg_shr_tmp[125]), .Z(N1224) );
  GTECH_AND2 C2296 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1223) );
  GTECH_NOT I_262 ( .A(N1226), .Z(m5stg_frac_pre3_in[11]) );
  GTECH_AND2 C2298 ( .A(N1225), .B(m4stg_shr_tmp[124]), .Z(N1226) );
  GTECH_AND2 C2299 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1225) );
  GTECH_NOT I_263 ( .A(N1228), .Z(m5stg_frac_pre3_in[10]) );
  GTECH_AND2 C2301 ( .A(N1227), .B(m4stg_shr_tmp[123]), .Z(N1228) );
  GTECH_AND2 C2302 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1227) );
  GTECH_NOT I_264 ( .A(N1230), .Z(m5stg_frac_pre3_in[9]) );
  GTECH_AND2 C2304 ( .A(N1229), .B(m4stg_shr_tmp[122]), .Z(N1230) );
  GTECH_AND2 C2305 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1229) );
  GTECH_NOT I_265 ( .A(N1232), .Z(m5stg_frac_pre3_in[8]) );
  GTECH_AND2 C2307 ( .A(N1231), .B(m4stg_shr_tmp[121]), .Z(N1232) );
  GTECH_AND2 C2308 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1231) );
  GTECH_NOT I_266 ( .A(N1234), .Z(m5stg_frac_pre3_in[7]) );
  GTECH_AND2 C2310 ( .A(N1233), .B(m4stg_shr_tmp[120]), .Z(N1234) );
  GTECH_AND2 C2311 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1233) );
  GTECH_NOT I_267 ( .A(N1236), .Z(m5stg_frac_pre3_in[6]) );
  GTECH_AND2 C2313 ( .A(N1235), .B(m4stg_shr_tmp[119]), .Z(N1236) );
  GTECH_AND2 C2314 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1235) );
  GTECH_NOT I_268 ( .A(N1238), .Z(m5stg_frac_pre3_in[5]) );
  GTECH_AND2 C2316 ( .A(N1237), .B(m4stg_shr_tmp[118]), .Z(N1238) );
  GTECH_AND2 C2317 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1237) );
  GTECH_NOT I_269 ( .A(N1240), .Z(m5stg_frac_pre3_in[4]) );
  GTECH_AND2 C2319 ( .A(N1239), .B(m4stg_shr_tmp[117]), .Z(N1240) );
  GTECH_AND2 C2320 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1239) );
  GTECH_NOT I_270 ( .A(N1242), .Z(m5stg_frac_pre3_in[3]) );
  GTECH_AND2 C2322 ( .A(N1241), .B(m4stg_shr_tmp[116]), .Z(N1242) );
  GTECH_AND2 C2323 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1241) );
  GTECH_NOT I_271 ( .A(N1244), .Z(m5stg_frac_pre3_in[2]) );
  GTECH_AND2 C2325 ( .A(N1243), .B(m4stg_shr_tmp[115]), .Z(N1244) );
  GTECH_AND2 C2326 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1243) );
  GTECH_NOT I_272 ( .A(N1246), .Z(m5stg_frac_pre3_in[1]) );
  GTECH_AND2 C2328 ( .A(N1245), .B(m4stg_shr_tmp[114]), .Z(N1246) );
  GTECH_AND2 C2329 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1245) );
  GTECH_NOT I_273 ( .A(N1248), .Z(m5stg_frac_pre3_in[0]) );
  GTECH_AND2 C2331 ( .A(N1247), .B(m4stg_shr[0]), .Z(N1248) );
  GTECH_AND2 C2332 ( .A(m4stg_right_shift_step), .B(m4stg_shr_tmp[168]), .Z(
        N1247) );
  GTECH_NOT I_274 ( .A(N1251), .Z(m5stg_frac_pre4_in[54]) );
  GTECH_AND2 C2334 ( .A(N1250), .B(m4stg_shr_tmp[166]), .Z(N1251) );
  GTECH_AND2 C2335 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1250) );
  GTECH_NOT I_275 ( .A(m4stg_shr_tmp[168]), .Z(N1249) );
  GTECH_NOT I_276 ( .A(N1253), .Z(m5stg_frac_pre4_in[53]) );
  GTECH_AND2 C2338 ( .A(N1252), .B(m4stg_shr_tmp[165]), .Z(N1253) );
  GTECH_AND2 C2339 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1252) );
  GTECH_NOT I_277 ( .A(N1255), .Z(m5stg_frac_pre4_in[52]) );
  GTECH_AND2 C2342 ( .A(N1254), .B(m4stg_shr_tmp[164]), .Z(N1255) );
  GTECH_AND2 C2343 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1254) );
  GTECH_NOT I_278 ( .A(N1257), .Z(m5stg_frac_pre4_in[51]) );
  GTECH_AND2 C2346 ( .A(N1256), .B(m4stg_shr_tmp[163]), .Z(N1257) );
  GTECH_AND2 C2347 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1256) );
  GTECH_NOT I_279 ( .A(N1259), .Z(m5stg_frac_pre4_in[50]) );
  GTECH_AND2 C2350 ( .A(N1258), .B(m4stg_shr_tmp[162]), .Z(N1259) );
  GTECH_AND2 C2351 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1258) );
  GTECH_NOT I_280 ( .A(N1261), .Z(m5stg_frac_pre4_in[49]) );
  GTECH_AND2 C2354 ( .A(N1260), .B(m4stg_shr_tmp[161]), .Z(N1261) );
  GTECH_AND2 C2355 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1260) );
  GTECH_NOT I_281 ( .A(N1263), .Z(m5stg_frac_pre4_in[48]) );
  GTECH_AND2 C2358 ( .A(N1262), .B(m4stg_shr_tmp[160]), .Z(N1263) );
  GTECH_AND2 C2359 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1262) );
  GTECH_NOT I_282 ( .A(N1265), .Z(m5stg_frac_pre4_in[47]) );
  GTECH_AND2 C2362 ( .A(N1264), .B(m4stg_shr_tmp[159]), .Z(N1265) );
  GTECH_AND2 C2363 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1264) );
  GTECH_NOT I_283 ( .A(N1267), .Z(m5stg_frac_pre4_in[46]) );
  GTECH_AND2 C2366 ( .A(N1266), .B(m4stg_shr_tmp[158]), .Z(N1267) );
  GTECH_AND2 C2367 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1266) );
  GTECH_NOT I_284 ( .A(N1269), .Z(m5stg_frac_pre4_in[45]) );
  GTECH_AND2 C2370 ( .A(N1268), .B(m4stg_shr_tmp[157]), .Z(N1269) );
  GTECH_AND2 C2371 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1268) );
  GTECH_NOT I_285 ( .A(N1271), .Z(m5stg_frac_pre4_in[44]) );
  GTECH_AND2 C2374 ( .A(N1270), .B(m4stg_shr_tmp[156]), .Z(N1271) );
  GTECH_AND2 C2375 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1270) );
  GTECH_NOT I_286 ( .A(N1273), .Z(m5stg_frac_pre4_in[43]) );
  GTECH_AND2 C2378 ( .A(N1272), .B(m4stg_shr_tmp[155]), .Z(N1273) );
  GTECH_AND2 C2379 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1272) );
  GTECH_NOT I_287 ( .A(N1275), .Z(m5stg_frac_pre4_in[42]) );
  GTECH_AND2 C2382 ( .A(N1274), .B(m4stg_shr_tmp[154]), .Z(N1275) );
  GTECH_AND2 C2383 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1274) );
  GTECH_NOT I_288 ( .A(N1277), .Z(m5stg_frac_pre4_in[41]) );
  GTECH_AND2 C2386 ( .A(N1276), .B(m4stg_shr_tmp[153]), .Z(N1277) );
  GTECH_AND2 C2387 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1276) );
  GTECH_NOT I_289 ( .A(N1279), .Z(m5stg_frac_pre4_in[40]) );
  GTECH_AND2 C2390 ( .A(N1278), .B(m4stg_shr_tmp[152]), .Z(N1279) );
  GTECH_AND2 C2391 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1278) );
  GTECH_NOT I_290 ( .A(N1281), .Z(m5stg_frac_pre4_in[39]) );
  GTECH_AND2 C2394 ( .A(N1280), .B(m4stg_shr_tmp[151]), .Z(N1281) );
  GTECH_AND2 C2395 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1280) );
  GTECH_NOT I_291 ( .A(N1283), .Z(m5stg_frac_pre4_in[38]) );
  GTECH_AND2 C2398 ( .A(N1282), .B(m4stg_shr_tmp[150]), .Z(N1283) );
  GTECH_AND2 C2399 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1282) );
  GTECH_NOT I_292 ( .A(N1285), .Z(m5stg_frac_pre4_in[37]) );
  GTECH_AND2 C2402 ( .A(N1284), .B(m4stg_shr_tmp[149]), .Z(N1285) );
  GTECH_AND2 C2403 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1284) );
  GTECH_NOT I_293 ( .A(N1287), .Z(m5stg_frac_pre4_in[36]) );
  GTECH_AND2 C2406 ( .A(N1286), .B(m4stg_shr_tmp[148]), .Z(N1287) );
  GTECH_AND2 C2407 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1286) );
  GTECH_NOT I_294 ( .A(N1289), .Z(m5stg_frac_pre4_in[35]) );
  GTECH_AND2 C2410 ( .A(N1288), .B(m4stg_shr_tmp[147]), .Z(N1289) );
  GTECH_AND2 C2411 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1288) );
  GTECH_NOT I_295 ( .A(N1291), .Z(m5stg_frac_pre4_in[34]) );
  GTECH_AND2 C2414 ( .A(N1290), .B(m4stg_shr_tmp[146]), .Z(N1291) );
  GTECH_AND2 C2415 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1290) );
  GTECH_NOT I_296 ( .A(N1293), .Z(m5stg_frac_pre4_in[33]) );
  GTECH_AND2 C2418 ( .A(N1292), .B(m4stg_shr_tmp[145]), .Z(N1293) );
  GTECH_AND2 C2419 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1292) );
  GTECH_NOT I_297 ( .A(N1295), .Z(m5stg_frac_pre4_in[32]) );
  GTECH_AND2 C2422 ( .A(N1294), .B(m4stg_shr_tmp[144]), .Z(N1295) );
  GTECH_AND2 C2423 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1294) );
  GTECH_NOT I_298 ( .A(N1297), .Z(m5stg_frac_pre4_in[31]) );
  GTECH_AND2 C2426 ( .A(N1296), .B(m4stg_shr_tmp[143]), .Z(N1297) );
  GTECH_AND2 C2427 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1296) );
  GTECH_NOT I_299 ( .A(N1299), .Z(m5stg_frac_pre4_in[30]) );
  GTECH_AND2 C2430 ( .A(N1298), .B(m4stg_shr_tmp[142]), .Z(N1299) );
  GTECH_AND2 C2431 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1298) );
  GTECH_NOT I_300 ( .A(N1301), .Z(m5stg_frac_pre4_in[29]) );
  GTECH_AND2 C2434 ( .A(N1300), .B(m4stg_shr_tmp[141]), .Z(N1301) );
  GTECH_AND2 C2435 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1300) );
  GTECH_NOT I_301 ( .A(N1303), .Z(m5stg_frac_pre4_in[28]) );
  GTECH_AND2 C2438 ( .A(N1302), .B(m4stg_shr_tmp[140]), .Z(N1303) );
  GTECH_AND2 C2439 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1302) );
  GTECH_NOT I_302 ( .A(N1305), .Z(m5stg_frac_pre4_in[27]) );
  GTECH_AND2 C2442 ( .A(N1304), .B(m4stg_shr_tmp[139]), .Z(N1305) );
  GTECH_AND2 C2443 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1304) );
  GTECH_NOT I_303 ( .A(N1307), .Z(m5stg_frac_pre4_in[26]) );
  GTECH_AND2 C2446 ( .A(N1306), .B(m4stg_shr_tmp[138]), .Z(N1307) );
  GTECH_AND2 C2447 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1306) );
  GTECH_NOT I_304 ( .A(N1309), .Z(m5stg_frac_pre4_in[25]) );
  GTECH_AND2 C2450 ( .A(N1308), .B(m4stg_shr_tmp[137]), .Z(N1309) );
  GTECH_AND2 C2451 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1308) );
  GTECH_NOT I_305 ( .A(N1311), .Z(m5stg_frac_pre4_in[24]) );
  GTECH_AND2 C2454 ( .A(N1310), .B(m4stg_shr_tmp[136]), .Z(N1311) );
  GTECH_AND2 C2455 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1310) );
  GTECH_NOT I_306 ( .A(N1313), .Z(m5stg_frac_pre4_in[23]) );
  GTECH_AND2 C2458 ( .A(N1312), .B(m4stg_shr_tmp[135]), .Z(N1313) );
  GTECH_AND2 C2459 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1312) );
  GTECH_NOT I_307 ( .A(N1315), .Z(m5stg_frac_pre4_in[22]) );
  GTECH_AND2 C2462 ( .A(N1314), .B(m4stg_shr_tmp[134]), .Z(N1315) );
  GTECH_AND2 C2463 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1314) );
  GTECH_NOT I_308 ( .A(N1317), .Z(m5stg_frac_pre4_in[21]) );
  GTECH_AND2 C2466 ( .A(N1316), .B(m4stg_shr_tmp[133]), .Z(N1317) );
  GTECH_AND2 C2467 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1316) );
  GTECH_NOT I_309 ( .A(N1319), .Z(m5stg_frac_pre4_in[20]) );
  GTECH_AND2 C2470 ( .A(N1318), .B(m4stg_shr_tmp[132]), .Z(N1319) );
  GTECH_AND2 C2471 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1318) );
  GTECH_NOT I_310 ( .A(N1321), .Z(m5stg_frac_pre4_in[19]) );
  GTECH_AND2 C2474 ( .A(N1320), .B(m4stg_shr_tmp[131]), .Z(N1321) );
  GTECH_AND2 C2475 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1320) );
  GTECH_NOT I_311 ( .A(N1323), .Z(m5stg_frac_pre4_in[18]) );
  GTECH_AND2 C2478 ( .A(N1322), .B(m4stg_shr_tmp[130]), .Z(N1323) );
  GTECH_AND2 C2479 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1322) );
  GTECH_NOT I_312 ( .A(N1325), .Z(m5stg_frac_pre4_in[17]) );
  GTECH_AND2 C2482 ( .A(N1324), .B(m4stg_shr_tmp[129]), .Z(N1325) );
  GTECH_AND2 C2483 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1324) );
  GTECH_NOT I_313 ( .A(N1327), .Z(m5stg_frac_pre4_in[16]) );
  GTECH_AND2 C2486 ( .A(N1326), .B(m4stg_shr_tmp[128]), .Z(N1327) );
  GTECH_AND2 C2487 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1326) );
  GTECH_NOT I_314 ( .A(N1329), .Z(m5stg_frac_pre4_in[15]) );
  GTECH_AND2 C2490 ( .A(N1328), .B(m4stg_shr_tmp[127]), .Z(N1329) );
  GTECH_AND2 C2491 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1328) );
  GTECH_NOT I_315 ( .A(N1331), .Z(m5stg_frac_pre4_in[14]) );
  GTECH_AND2 C2494 ( .A(N1330), .B(m4stg_shr_tmp[126]), .Z(N1331) );
  GTECH_AND2 C2495 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1330) );
  GTECH_NOT I_316 ( .A(N1333), .Z(m5stg_frac_pre4_in[13]) );
  GTECH_AND2 C2498 ( .A(N1332), .B(m4stg_shr_tmp[125]), .Z(N1333) );
  GTECH_AND2 C2499 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1332) );
  GTECH_NOT I_317 ( .A(N1335), .Z(m5stg_frac_pre4_in[12]) );
  GTECH_AND2 C2502 ( .A(N1334), .B(m4stg_shr_tmp[124]), .Z(N1335) );
  GTECH_AND2 C2503 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1334) );
  GTECH_NOT I_318 ( .A(N1337), .Z(m5stg_frac_pre4_in[11]) );
  GTECH_AND2 C2506 ( .A(N1336), .B(m4stg_shr_tmp[123]), .Z(N1337) );
  GTECH_AND2 C2507 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1336) );
  GTECH_NOT I_319 ( .A(N1339), .Z(m5stg_frac_pre4_in[10]) );
  GTECH_AND2 C2510 ( .A(N1338), .B(m4stg_shr_tmp[122]), .Z(N1339) );
  GTECH_AND2 C2511 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1338) );
  GTECH_NOT I_320 ( .A(N1341), .Z(m5stg_frac_pre4_in[9]) );
  GTECH_AND2 C2514 ( .A(N1340), .B(m4stg_shr_tmp[121]), .Z(N1341) );
  GTECH_AND2 C2515 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1340) );
  GTECH_NOT I_321 ( .A(N1343), .Z(m5stg_frac_pre4_in[8]) );
  GTECH_AND2 C2518 ( .A(N1342), .B(m4stg_shr_tmp[120]), .Z(N1343) );
  GTECH_AND2 C2519 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1342) );
  GTECH_NOT I_322 ( .A(N1345), .Z(m5stg_frac_pre4_in[7]) );
  GTECH_AND2 C2522 ( .A(N1344), .B(m4stg_shr_tmp[119]), .Z(N1345) );
  GTECH_AND2 C2523 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1344) );
  GTECH_NOT I_323 ( .A(N1347), .Z(m5stg_frac_pre4_in[6]) );
  GTECH_AND2 C2526 ( .A(N1346), .B(m4stg_shr_tmp[118]), .Z(N1347) );
  GTECH_AND2 C2527 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1346) );
  GTECH_NOT I_324 ( .A(N1349), .Z(m5stg_frac_pre4_in[5]) );
  GTECH_AND2 C2530 ( .A(N1348), .B(m4stg_shr_tmp[117]), .Z(N1349) );
  GTECH_AND2 C2531 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1348) );
  GTECH_NOT I_325 ( .A(N1351), .Z(m5stg_frac_pre4_in[4]) );
  GTECH_AND2 C2534 ( .A(N1350), .B(m4stg_shr_tmp[116]), .Z(N1351) );
  GTECH_AND2 C2535 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1350) );
  GTECH_NOT I_326 ( .A(N1353), .Z(m5stg_frac_pre4_in[3]) );
  GTECH_AND2 C2538 ( .A(N1352), .B(m4stg_shr_tmp[115]), .Z(N1353) );
  GTECH_AND2 C2539 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1352) );
  GTECH_NOT I_327 ( .A(N1355), .Z(m5stg_frac_pre4_in[2]) );
  GTECH_AND2 C2542 ( .A(N1354), .B(m4stg_shr_tmp[114]), .Z(N1355) );
  GTECH_AND2 C2543 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1354) );
  GTECH_NOT I_328 ( .A(N1357), .Z(m5stg_frac_pre4_in[1]) );
  GTECH_AND2 C2546 ( .A(N1356), .B(m4stg_shr[0]), .Z(N1357) );
  GTECH_AND2 C2547 ( .A(m4stg_right_shift_step), .B(N1249), .Z(N1356) );
  GTECH_NOT I_329 ( .A(N1360), .Z(m5stg_frac_54_33[54]) );
  GTECH_AND2 C2550 ( .A(N1359), .B(m5stg_frac_pre4[54]), .Z(N1360) );
  GTECH_AND2 C2551 ( .A(N1358), .B(m5stg_frac_pre3[54]), .Z(N1359) );
  GTECH_AND2 C2552 ( .A(m5stg_frac_pre1[54]), .B(m5stg_frac_pre2[54]), .Z(
        N1358) );
  GTECH_NOT I_330 ( .A(N1363), .Z(m5stg_frac_54_33[53]) );
  GTECH_AND2 C2554 ( .A(N1362), .B(m5stg_frac_pre4[53]), .Z(N1363) );
  GTECH_AND2 C2555 ( .A(N1361), .B(m5stg_frac_pre3[53]), .Z(N1362) );
  GTECH_AND2 C2556 ( .A(m5stg_frac_pre1[53]), .B(m5stg_frac_pre2[53]), .Z(
        N1361) );
  GTECH_NOT I_331 ( .A(N1366), .Z(m5stg_frac_54_33[52]) );
  GTECH_AND2 C2558 ( .A(N1365), .B(m5stg_frac_pre4[52]), .Z(N1366) );
  GTECH_AND2 C2559 ( .A(N1364), .B(m5stg_frac_pre3[52]), .Z(N1365) );
  GTECH_AND2 C2560 ( .A(m5stg_frac_pre1[52]), .B(m5stg_frac_pre2[52]), .Z(
        N1364) );
  GTECH_NOT I_332 ( .A(N1369), .Z(m5stg_frac_54_33[51]) );
  GTECH_AND2 C2562 ( .A(N1368), .B(m5stg_frac_pre4[51]), .Z(N1369) );
  GTECH_AND2 C2563 ( .A(N1367), .B(m5stg_frac_pre3[51]), .Z(N1368) );
  GTECH_AND2 C2564 ( .A(m5stg_frac_pre1[51]), .B(m5stg_frac_pre2[51]), .Z(
        N1367) );
  GTECH_NOT I_333 ( .A(N1372), .Z(m5stg_frac_54_33[50]) );
  GTECH_AND2 C2566 ( .A(N1371), .B(m5stg_frac_pre4[50]), .Z(N1372) );
  GTECH_AND2 C2567 ( .A(N1370), .B(m5stg_frac_pre3[50]), .Z(N1371) );
  GTECH_AND2 C2568 ( .A(m5stg_frac_pre1[50]), .B(m5stg_frac_pre2[50]), .Z(
        N1370) );
  GTECH_NOT I_334 ( .A(N1375), .Z(m5stg_frac_54_33[49]) );
  GTECH_AND2 C2570 ( .A(N1374), .B(m5stg_frac_pre4[49]), .Z(N1375) );
  GTECH_AND2 C2571 ( .A(N1373), .B(m5stg_frac_pre3[49]), .Z(N1374) );
  GTECH_AND2 C2572 ( .A(m5stg_frac_pre1[49]), .B(m5stg_frac_pre2[49]), .Z(
        N1373) );
  GTECH_NOT I_335 ( .A(N1378), .Z(m5stg_frac_54_33[48]) );
  GTECH_AND2 C2574 ( .A(N1377), .B(m5stg_frac_pre4[48]), .Z(N1378) );
  GTECH_AND2 C2575 ( .A(N1376), .B(m5stg_frac_pre3[48]), .Z(N1377) );
  GTECH_AND2 C2576 ( .A(m5stg_frac_pre1[48]), .B(m5stg_frac_pre2[48]), .Z(
        N1376) );
  GTECH_NOT I_336 ( .A(N1381), .Z(m5stg_frac_54_33[47]) );
  GTECH_AND2 C2578 ( .A(N1380), .B(m5stg_frac_pre4[47]), .Z(N1381) );
  GTECH_AND2 C2579 ( .A(N1379), .B(m5stg_frac_pre3[47]), .Z(N1380) );
  GTECH_AND2 C2580 ( .A(m5stg_frac_pre1[47]), .B(m5stg_frac_pre2[47]), .Z(
        N1379) );
  GTECH_NOT I_337 ( .A(N1384), .Z(m5stg_frac_54_33[46]) );
  GTECH_AND2 C2582 ( .A(N1383), .B(m5stg_frac_pre4[46]), .Z(N1384) );
  GTECH_AND2 C2583 ( .A(N1382), .B(m5stg_frac_pre3[46]), .Z(N1383) );
  GTECH_AND2 C2584 ( .A(m5stg_frac_pre1[46]), .B(m5stg_frac_pre2[46]), .Z(
        N1382) );
  GTECH_NOT I_338 ( .A(N1387), .Z(m5stg_frac_54_33[45]) );
  GTECH_AND2 C2586 ( .A(N1386), .B(m5stg_frac_pre4[45]), .Z(N1387) );
  GTECH_AND2 C2587 ( .A(N1385), .B(m5stg_frac_pre3[45]), .Z(N1386) );
  GTECH_AND2 C2588 ( .A(m5stg_frac_pre1[45]), .B(m5stg_frac_pre2[45]), .Z(
        N1385) );
  GTECH_NOT I_339 ( .A(N1390), .Z(m5stg_frac_54_33[44]) );
  GTECH_AND2 C2590 ( .A(N1389), .B(m5stg_frac_pre4[44]), .Z(N1390) );
  GTECH_AND2 C2591 ( .A(N1388), .B(m5stg_frac_pre3[44]), .Z(N1389) );
  GTECH_AND2 C2592 ( .A(m5stg_frac_pre1[44]), .B(m5stg_frac_pre2[44]), .Z(
        N1388) );
  GTECH_NOT I_340 ( .A(N1393), .Z(m5stg_frac_54_33[43]) );
  GTECH_AND2 C2594 ( .A(N1392), .B(m5stg_frac_pre4[43]), .Z(N1393) );
  GTECH_AND2 C2595 ( .A(N1391), .B(m5stg_frac_pre3[43]), .Z(N1392) );
  GTECH_AND2 C2596 ( .A(m5stg_frac_pre1[43]), .B(m5stg_frac_pre2[43]), .Z(
        N1391) );
  GTECH_NOT I_341 ( .A(N1396), .Z(m5stg_frac_54_33[42]) );
  GTECH_AND2 C2598 ( .A(N1395), .B(m5stg_frac_pre4[42]), .Z(N1396) );
  GTECH_AND2 C2599 ( .A(N1394), .B(m5stg_frac_pre3[42]), .Z(N1395) );
  GTECH_AND2 C2600 ( .A(m5stg_frac_pre1[42]), .B(m5stg_frac_pre2[42]), .Z(
        N1394) );
  GTECH_NOT I_342 ( .A(N1399), .Z(m5stg_frac_54_33[41]) );
  GTECH_AND2 C2602 ( .A(N1398), .B(m5stg_frac_pre4[41]), .Z(N1399) );
  GTECH_AND2 C2603 ( .A(N1397), .B(m5stg_frac_pre3[41]), .Z(N1398) );
  GTECH_AND2 C2604 ( .A(m5stg_frac_pre1[41]), .B(m5stg_frac_pre2[41]), .Z(
        N1397) );
  GTECH_NOT I_343 ( .A(N1402), .Z(m5stg_frac_54_33[40]) );
  GTECH_AND2 C2606 ( .A(N1401), .B(m5stg_frac_pre4[40]), .Z(N1402) );
  GTECH_AND2 C2607 ( .A(N1400), .B(m5stg_frac_pre3[40]), .Z(N1401) );
  GTECH_AND2 C2608 ( .A(m5stg_frac_pre1[40]), .B(m5stg_frac_pre2[40]), .Z(
        N1400) );
  GTECH_NOT I_344 ( .A(N1405), .Z(m5stg_frac_54_33[39]) );
  GTECH_AND2 C2610 ( .A(N1404), .B(m5stg_frac_pre4[39]), .Z(N1405) );
  GTECH_AND2 C2611 ( .A(N1403), .B(m5stg_frac_pre3[39]), .Z(N1404) );
  GTECH_AND2 C2612 ( .A(m5stg_frac_pre1[39]), .B(m5stg_frac_pre2[39]), .Z(
        N1403) );
  GTECH_NOT I_345 ( .A(N1408), .Z(m5stg_frac_54_33[38]) );
  GTECH_AND2 C2614 ( .A(N1407), .B(m5stg_frac_pre4[38]), .Z(N1408) );
  GTECH_AND2 C2615 ( .A(N1406), .B(m5stg_frac_pre3[38]), .Z(N1407) );
  GTECH_AND2 C2616 ( .A(m5stg_frac_pre1[38]), .B(m5stg_frac_pre2[38]), .Z(
        N1406) );
  GTECH_NOT I_346 ( .A(N1411), .Z(m5stg_frac_54_33[37]) );
  GTECH_AND2 C2618 ( .A(N1410), .B(m5stg_frac_pre4[37]), .Z(N1411) );
  GTECH_AND2 C2619 ( .A(N1409), .B(m5stg_frac_pre3[37]), .Z(N1410) );
  GTECH_AND2 C2620 ( .A(m5stg_frac_pre1[37]), .B(m5stg_frac_pre2[37]), .Z(
        N1409) );
  GTECH_NOT I_347 ( .A(N1414), .Z(m5stg_frac_54_33[36]) );
  GTECH_AND2 C2622 ( .A(N1413), .B(m5stg_frac_pre4[36]), .Z(N1414) );
  GTECH_AND2 C2623 ( .A(N1412), .B(m5stg_frac_pre3[36]), .Z(N1413) );
  GTECH_AND2 C2624 ( .A(m5stg_frac_pre1[36]), .B(m5stg_frac_pre2[36]), .Z(
        N1412) );
  GTECH_NOT I_348 ( .A(N1417), .Z(m5stg_frac_54_33[35]) );
  GTECH_AND2 C2626 ( .A(N1416), .B(m5stg_frac_pre4[35]), .Z(N1417) );
  GTECH_AND2 C2627 ( .A(N1415), .B(m5stg_frac_pre3[35]), .Z(N1416) );
  GTECH_AND2 C2628 ( .A(m5stg_frac_pre1[35]), .B(m5stg_frac_pre2[35]), .Z(
        N1415) );
  GTECH_NOT I_349 ( .A(N1420), .Z(m5stg_frac_54_33[34]) );
  GTECH_AND2 C2630 ( .A(N1419), .B(m5stg_frac_pre4[34]), .Z(N1420) );
  GTECH_AND2 C2631 ( .A(N1418), .B(m5stg_frac_pre3[34]), .Z(N1419) );
  GTECH_AND2 C2632 ( .A(m5stg_frac_pre1[34]), .B(m5stg_frac_pre2[34]), .Z(
        N1418) );
  GTECH_NOT I_350 ( .A(N1423), .Z(m5stg_frac_54_33[33]) );
  GTECH_AND2 C2634 ( .A(N1422), .B(m5stg_frac_pre4[33]), .Z(N1423) );
  GTECH_AND2 C2635 ( .A(N1421), .B(m5stg_frac_pre3[33]), .Z(N1422) );
  GTECH_AND2 C2636 ( .A(m5stg_frac_pre1[33]), .B(m5stg_frac_pre2[33]), .Z(
        N1421) );
  GTECH_NOT I_351 ( .A(N1426), .Z(m5stg_frac_32_0[32]) );
  GTECH_AND2 C2638 ( .A(N1425), .B(m5stg_frac_pre4[32]), .Z(N1426) );
  GTECH_AND2 C2639 ( .A(N1424), .B(m5stg_frac_pre3[32]), .Z(N1425) );
  GTECH_AND2 C2640 ( .A(m5stg_frac_pre1[32]), .B(m5stg_frac_pre2[32]), .Z(
        N1424) );
  GTECH_NOT I_352 ( .A(N1429), .Z(m5stg_frac_32_0[31]) );
  GTECH_AND2 C2642 ( .A(N1428), .B(m5stg_frac_pre4[31]), .Z(N1429) );
  GTECH_AND2 C2643 ( .A(N1427), .B(m5stg_frac_pre3[31]), .Z(N1428) );
  GTECH_AND2 C2644 ( .A(m5stg_frac_pre1[31]), .B(m5stg_frac_pre2[31]), .Z(
        N1427) );
  GTECH_NOT I_353 ( .A(N1432), .Z(m5stg_frac_32_0[30]) );
  GTECH_AND2 C2646 ( .A(N1431), .B(m5stg_frac_pre4[30]), .Z(N1432) );
  GTECH_AND2 C2647 ( .A(N1430), .B(m5stg_frac_pre3[30]), .Z(N1431) );
  GTECH_AND2 C2648 ( .A(m5stg_frac_pre1[30]), .B(m5stg_frac_pre2[30]), .Z(
        N1430) );
  GTECH_NOT I_354 ( .A(N1435), .Z(m5stg_frac_32_0[29]) );
  GTECH_AND2 C2650 ( .A(N1434), .B(m5stg_frac_pre4[29]), .Z(N1435) );
  GTECH_AND2 C2651 ( .A(N1433), .B(m5stg_frac_pre3[29]), .Z(N1434) );
  GTECH_AND2 C2652 ( .A(m5stg_frac_pre1[29]), .B(m5stg_frac_pre2[29]), .Z(
        N1433) );
  GTECH_NOT I_355 ( .A(N1438), .Z(m5stg_frac_32_0[28]) );
  GTECH_AND2 C2654 ( .A(N1437), .B(m5stg_frac_pre4[28]), .Z(N1438) );
  GTECH_AND2 C2655 ( .A(N1436), .B(m5stg_frac_pre3[28]), .Z(N1437) );
  GTECH_AND2 C2656 ( .A(m5stg_frac_pre1[28]), .B(m5stg_frac_pre2[28]), .Z(
        N1436) );
  GTECH_NOT I_356 ( .A(N1441), .Z(m5stg_frac_32_0[27]) );
  GTECH_AND2 C2658 ( .A(N1440), .B(m5stg_frac_pre4[27]), .Z(N1441) );
  GTECH_AND2 C2659 ( .A(N1439), .B(m5stg_frac_pre3[27]), .Z(N1440) );
  GTECH_AND2 C2660 ( .A(m5stg_frac_pre1[27]), .B(m5stg_frac_pre2[27]), .Z(
        N1439) );
  GTECH_NOT I_357 ( .A(N1444), .Z(m5stg_frac_32_0[26]) );
  GTECH_AND2 C2662 ( .A(N1443), .B(m5stg_frac_pre4[26]), .Z(N1444) );
  GTECH_AND2 C2663 ( .A(N1442), .B(m5stg_frac_pre3[26]), .Z(N1443) );
  GTECH_AND2 C2664 ( .A(m5stg_frac_pre1[26]), .B(m5stg_frac_pre2[26]), .Z(
        N1442) );
  GTECH_NOT I_358 ( .A(N1447), .Z(m5stg_frac_32_0[25]) );
  GTECH_AND2 C2666 ( .A(N1446), .B(m5stg_frac_pre4[25]), .Z(N1447) );
  GTECH_AND2 C2667 ( .A(N1445), .B(m5stg_frac_pre3[25]), .Z(N1446) );
  GTECH_AND2 C2668 ( .A(m5stg_frac_pre1[25]), .B(m5stg_frac_pre2[25]), .Z(
        N1445) );
  GTECH_NOT I_359 ( .A(N1450), .Z(m5stg_frac_32_0[24]) );
  GTECH_AND2 C2670 ( .A(N1449), .B(m5stg_frac_pre4[24]), .Z(N1450) );
  GTECH_AND2 C2671 ( .A(N1448), .B(m5stg_frac_pre3[24]), .Z(N1449) );
  GTECH_AND2 C2672 ( .A(m5stg_frac_pre1[24]), .B(m5stg_frac_pre2[24]), .Z(
        N1448) );
  GTECH_NOT I_360 ( .A(N1453), .Z(m5stg_frac_32_0[23]) );
  GTECH_AND2 C2674 ( .A(N1452), .B(m5stg_frac_pre4[23]), .Z(N1453) );
  GTECH_AND2 C2675 ( .A(N1451), .B(m5stg_frac_pre3[23]), .Z(N1452) );
  GTECH_AND2 C2676 ( .A(m5stg_frac_pre1[23]), .B(m5stg_frac_pre2[23]), .Z(
        N1451) );
  GTECH_NOT I_361 ( .A(N1456), .Z(m5stg_frac_32_0[22]) );
  GTECH_AND2 C2678 ( .A(N1455), .B(m5stg_frac_pre4[22]), .Z(N1456) );
  GTECH_AND2 C2679 ( .A(N1454), .B(m5stg_frac_pre3[22]), .Z(N1455) );
  GTECH_AND2 C2680 ( .A(m5stg_frac_pre1[22]), .B(m5stg_frac_pre2[22]), .Z(
        N1454) );
  GTECH_NOT I_362 ( .A(N1459), .Z(m5stg_frac_32_0[21]) );
  GTECH_AND2 C2682 ( .A(N1458), .B(m5stg_frac_pre4[21]), .Z(N1459) );
  GTECH_AND2 C2683 ( .A(N1457), .B(m5stg_frac_pre3[21]), .Z(N1458) );
  GTECH_AND2 C2684 ( .A(m5stg_frac_pre1[21]), .B(m5stg_frac_pre2[21]), .Z(
        N1457) );
  GTECH_NOT I_363 ( .A(N1462), .Z(m5stg_frac_32_0[20]) );
  GTECH_AND2 C2686 ( .A(N1461), .B(m5stg_frac_pre4[20]), .Z(N1462) );
  GTECH_AND2 C2687 ( .A(N1460), .B(m5stg_frac_pre3[20]), .Z(N1461) );
  GTECH_AND2 C2688 ( .A(m5stg_frac_pre1[20]), .B(m5stg_frac_pre2[20]), .Z(
        N1460) );
  GTECH_NOT I_364 ( .A(N1465), .Z(m5stg_frac_32_0[19]) );
  GTECH_AND2 C2690 ( .A(N1464), .B(m5stg_frac_pre4[19]), .Z(N1465) );
  GTECH_AND2 C2691 ( .A(N1463), .B(m5stg_frac_pre3[19]), .Z(N1464) );
  GTECH_AND2 C2692 ( .A(m5stg_frac_pre1[19]), .B(m5stg_frac_pre2[19]), .Z(
        N1463) );
  GTECH_NOT I_365 ( .A(N1468), .Z(m5stg_frac_32_0[18]) );
  GTECH_AND2 C2694 ( .A(N1467), .B(m5stg_frac_pre4[18]), .Z(N1468) );
  GTECH_AND2 C2695 ( .A(N1466), .B(m5stg_frac_pre3[18]), .Z(N1467) );
  GTECH_AND2 C2696 ( .A(m5stg_frac_pre1[18]), .B(m5stg_frac_pre2[18]), .Z(
        N1466) );
  GTECH_NOT I_366 ( .A(N1471), .Z(m5stg_frac_32_0[17]) );
  GTECH_AND2 C2698 ( .A(N1470), .B(m5stg_frac_pre4[17]), .Z(N1471) );
  GTECH_AND2 C2699 ( .A(N1469), .B(m5stg_frac_pre3[17]), .Z(N1470) );
  GTECH_AND2 C2700 ( .A(m5stg_frac_pre1[17]), .B(m5stg_frac_pre2[17]), .Z(
        N1469) );
  GTECH_NOT I_367 ( .A(N1474), .Z(m5stg_frac_32_0[16]) );
  GTECH_AND2 C2702 ( .A(N1473), .B(m5stg_frac_pre4[16]), .Z(N1474) );
  GTECH_AND2 C2703 ( .A(N1472), .B(m5stg_frac_pre3[16]), .Z(N1473) );
  GTECH_AND2 C2704 ( .A(m5stg_frac_pre1[16]), .B(m5stg_frac_pre2[16]), .Z(
        N1472) );
  GTECH_NOT I_368 ( .A(N1477), .Z(m5stg_frac_32_0[15]) );
  GTECH_AND2 C2706 ( .A(N1476), .B(m5stg_frac_pre4[15]), .Z(N1477) );
  GTECH_AND2 C2707 ( .A(N1475), .B(m5stg_frac_pre3[15]), .Z(N1476) );
  GTECH_AND2 C2708 ( .A(m5stg_frac_pre1[15]), .B(m5stg_frac_pre2[15]), .Z(
        N1475) );
  GTECH_NOT I_369 ( .A(N1480), .Z(m5stg_frac_32_0[14]) );
  GTECH_AND2 C2710 ( .A(N1479), .B(m5stg_frac_pre4[14]), .Z(N1480) );
  GTECH_AND2 C2711 ( .A(N1478), .B(m5stg_frac_pre3[14]), .Z(N1479) );
  GTECH_AND2 C2712 ( .A(m5stg_frac_pre1[14]), .B(m5stg_frac_pre2[14]), .Z(
        N1478) );
  GTECH_NOT I_370 ( .A(N1483), .Z(m5stg_frac_32_0[13]) );
  GTECH_AND2 C2714 ( .A(N1482), .B(m5stg_frac_pre4[13]), .Z(N1483) );
  GTECH_AND2 C2715 ( .A(N1481), .B(m5stg_frac_pre3[13]), .Z(N1482) );
  GTECH_AND2 C2716 ( .A(m5stg_frac_pre1[13]), .B(m5stg_frac_pre2[13]), .Z(
        N1481) );
  GTECH_NOT I_371 ( .A(N1486), .Z(m5stg_frac_32_0[12]) );
  GTECH_AND2 C2718 ( .A(N1485), .B(m5stg_frac_pre4[12]), .Z(N1486) );
  GTECH_AND2 C2719 ( .A(N1484), .B(m5stg_frac_pre3[12]), .Z(N1485) );
  GTECH_AND2 C2720 ( .A(m5stg_frac_pre1[12]), .B(m5stg_frac_pre2[12]), .Z(
        N1484) );
  GTECH_NOT I_372 ( .A(N1489), .Z(m5stg_frac_32_0[11]) );
  GTECH_AND2 C2722 ( .A(N1488), .B(m5stg_frac_pre4[11]), .Z(N1489) );
  GTECH_AND2 C2723 ( .A(N1487), .B(m5stg_frac_pre3[11]), .Z(N1488) );
  GTECH_AND2 C2724 ( .A(m5stg_frac_pre1[11]), .B(m5stg_frac_pre2[11]), .Z(
        N1487) );
  GTECH_NOT I_373 ( .A(N1492), .Z(m5stg_frac_32_0[10]) );
  GTECH_AND2 C2726 ( .A(N1491), .B(m5stg_frac_pre4[10]), .Z(N1492) );
  GTECH_AND2 C2727 ( .A(N1490), .B(m5stg_frac_pre3[10]), .Z(N1491) );
  GTECH_AND2 C2728 ( .A(m5stg_frac_pre1[10]), .B(m5stg_frac_pre2[10]), .Z(
        N1490) );
  GTECH_NOT I_374 ( .A(N1495), .Z(m5stg_frac_32_0[9]) );
  GTECH_AND2 C2730 ( .A(N1494), .B(m5stg_frac_pre4[9]), .Z(N1495) );
  GTECH_AND2 C2731 ( .A(N1493), .B(m5stg_frac_pre3[9]), .Z(N1494) );
  GTECH_AND2 C2732 ( .A(m5stg_frac_pre1[9]), .B(m5stg_frac_pre2[9]), .Z(N1493)
         );
  GTECH_NOT I_375 ( .A(N1498), .Z(m5stg_frac_32_0[8]) );
  GTECH_AND2 C2734 ( .A(N1497), .B(m5stg_frac_pre4[8]), .Z(N1498) );
  GTECH_AND2 C2735 ( .A(N1496), .B(m5stg_frac_pre3[8]), .Z(N1497) );
  GTECH_AND2 C2736 ( .A(m5stg_frac_pre1[8]), .B(m5stg_frac_pre2[8]), .Z(N1496)
         );
  GTECH_NOT I_376 ( .A(N1501), .Z(m5stg_frac_32_0[7]) );
  GTECH_AND2 C2738 ( .A(N1500), .B(m5stg_frac_pre4[7]), .Z(N1501) );
  GTECH_AND2 C2739 ( .A(N1499), .B(m5stg_frac_pre3[7]), .Z(N1500) );
  GTECH_AND2 C2740 ( .A(m5stg_frac_pre1[7]), .B(m5stg_frac_pre2[7]), .Z(N1499)
         );
  GTECH_NOT I_377 ( .A(N1504), .Z(m5stg_frac_32_0[6]) );
  GTECH_AND2 C2742 ( .A(N1503), .B(m5stg_frac_pre4[6]), .Z(N1504) );
  GTECH_AND2 C2743 ( .A(N1502), .B(m5stg_frac_pre3[6]), .Z(N1503) );
  GTECH_AND2 C2744 ( .A(m5stg_frac_pre1[6]), .B(m5stg_frac_pre2[6]), .Z(N1502)
         );
  GTECH_NOT I_378 ( .A(N1507), .Z(m5stg_frac_32_0[5]) );
  GTECH_AND2 C2746 ( .A(N1506), .B(m5stg_frac_pre4[5]), .Z(N1507) );
  GTECH_AND2 C2747 ( .A(N1505), .B(m5stg_frac_pre3[5]), .Z(N1506) );
  GTECH_AND2 C2748 ( .A(m5stg_frac_pre1[5]), .B(m5stg_frac_pre2[5]), .Z(N1505)
         );
  GTECH_NOT I_379 ( .A(N1510), .Z(m5stg_frac_32_0[4]) );
  GTECH_AND2 C2750 ( .A(N1509), .B(m5stg_frac_pre4[4]), .Z(N1510) );
  GTECH_AND2 C2751 ( .A(N1508), .B(m5stg_frac_pre3[4]), .Z(N1509) );
  GTECH_AND2 C2752 ( .A(m5stg_frac_pre1[4]), .B(m5stg_frac_pre2[4]), .Z(N1508)
         );
  GTECH_NOT I_380 ( .A(N1513), .Z(m5stg_frac_32_0[3]) );
  GTECH_AND2 C2754 ( .A(N1512), .B(m5stg_frac_pre4[3]), .Z(N1513) );
  GTECH_AND2 C2755 ( .A(N1511), .B(m5stg_frac_pre3[3]), .Z(N1512) );
  GTECH_AND2 C2756 ( .A(m5stg_frac_pre1[3]), .B(m5stg_frac_pre2[3]), .Z(N1511)
         );
  GTECH_NOT I_381 ( .A(N1516), .Z(m5stg_frac_32_0[2]) );
  GTECH_AND2 C2758 ( .A(N1515), .B(m5stg_frac_pre4[2]), .Z(N1516) );
  GTECH_AND2 C2759 ( .A(N1514), .B(m5stg_frac_pre3[2]), .Z(N1515) );
  GTECH_AND2 C2760 ( .A(m5stg_frac_pre1[2]), .B(m5stg_frac_pre2[2]), .Z(N1514)
         );
  GTECH_NOT I_382 ( .A(N1519), .Z(m5stg_frac_32_0[1]) );
  GTECH_AND2 C2762 ( .A(N1518), .B(m5stg_frac_pre4[1]), .Z(N1519) );
  GTECH_AND2 C2763 ( .A(N1517), .B(m5stg_frac_pre3[1]), .Z(N1518) );
  GTECH_AND2 C2764 ( .A(m5stg_frac_pre1[1]), .B(m5stg_frac_pre2[1]), .Z(N1517)
         );
  GTECH_NOT I_383 ( .A(N1522), .Z(m5stg_frac_32_0[0]) );
  GTECH_AND2 C2766 ( .A(N1521), .B(m5stg_frac_pre4[0]), .Z(N1522) );
  GTECH_AND2 C2767 ( .A(N1520), .B(m5stg_frac_pre3[0]), .Z(N1521) );
  GTECH_AND2 C2768 ( .A(m5stg_frac_pre1[0]), .B(m5stg_frac_pre2[0]), .Z(N1520)
         );
  GTECH_OR2 C2769 ( .A(N1523), .B(m5stg_frac_32_0[0]), .Z(m5stg_frac_dbl_nx)
         );
  GTECH_OR2 C2770 ( .A(m5stg_frac_32_0[2]), .B(m5stg_frac_32_0[1]), .Z(N1523)
         );
  GTECH_OR2 C2771 ( .A(m5stg_frac_dbl_nx), .B(N1551), .Z(m5stg_frac_sng_nx) );
  GTECH_OR2 C2772 ( .A(N1550), .B(m5stg_frac_32_0[3]), .Z(N1551) );
  GTECH_OR2 C2773 ( .A(N1549), .B(m5stg_frac_32_0[4]), .Z(N1550) );
  GTECH_OR2 C2774 ( .A(N1548), .B(m5stg_frac_32_0[5]), .Z(N1549) );
  GTECH_OR2 C2775 ( .A(N1547), .B(m5stg_frac_32_0[6]), .Z(N1548) );
  GTECH_OR2 C2776 ( .A(N1546), .B(m5stg_frac_32_0[7]), .Z(N1547) );
  GTECH_OR2 C2777 ( .A(N1545), .B(m5stg_frac_32_0[8]), .Z(N1546) );
  GTECH_OR2 C2778 ( .A(N1544), .B(m5stg_frac_32_0[9]), .Z(N1545) );
  GTECH_OR2 C2779 ( .A(N1543), .B(m5stg_frac_32_0[10]), .Z(N1544) );
  GTECH_OR2 C2780 ( .A(N1542), .B(m5stg_frac_32_0[11]), .Z(N1543) );
  GTECH_OR2 C2781 ( .A(N1541), .B(m5stg_frac_32_0[12]), .Z(N1542) );
  GTECH_OR2 C2782 ( .A(N1540), .B(m5stg_frac_32_0[13]), .Z(N1541) );
  GTECH_OR2 C2783 ( .A(N1539), .B(m5stg_frac_32_0[14]), .Z(N1540) );
  GTECH_OR2 C2784 ( .A(N1538), .B(m5stg_frac_32_0[15]), .Z(N1539) );
  GTECH_OR2 C2785 ( .A(N1537), .B(m5stg_frac_32_0[16]), .Z(N1538) );
  GTECH_OR2 C2786 ( .A(N1536), .B(m5stg_frac_32_0[17]), .Z(N1537) );
  GTECH_OR2 C2787 ( .A(N1535), .B(m5stg_frac_32_0[18]), .Z(N1536) );
  GTECH_OR2 C2788 ( .A(N1534), .B(m5stg_frac_32_0[19]), .Z(N1535) );
  GTECH_OR2 C2789 ( .A(N1533), .B(m5stg_frac_32_0[20]), .Z(N1534) );
  GTECH_OR2 C2790 ( .A(N1532), .B(m5stg_frac_32_0[21]), .Z(N1533) );
  GTECH_OR2 C2791 ( .A(N1531), .B(m5stg_frac_32_0[22]), .Z(N1532) );
  GTECH_OR2 C2792 ( .A(N1530), .B(m5stg_frac_32_0[23]), .Z(N1531) );
  GTECH_OR2 C2793 ( .A(N1529), .B(m5stg_frac_32_0[24]), .Z(N1530) );
  GTECH_OR2 C2794 ( .A(N1528), .B(m5stg_frac_32_0[25]), .Z(N1529) );
  GTECH_OR2 C2795 ( .A(N1527), .B(m5stg_frac_32_0[26]), .Z(N1528) );
  GTECH_OR2 C2796 ( .A(N1526), .B(m5stg_frac_32_0[27]), .Z(N1527) );
  GTECH_OR2 C2797 ( .A(N1525), .B(m5stg_frac_32_0[28]), .Z(N1526) );
  GTECH_OR2 C2798 ( .A(N1524), .B(m5stg_frac_32_0[29]), .Z(N1525) );
  GTECH_OR2 C2799 ( .A(m5stg_frac_32_0[31]), .B(m5stg_frac_32_0[30]), .Z(N1524) );
  GTECH_OR2 C2800 ( .A(m5stg_frac_sng_nx), .B(N1573), .Z(m5stg_frac_neq_0) );
  GTECH_OR2 C2801 ( .A(N1572), .B(m5stg_frac_32_0[32]), .Z(N1573) );
  GTECH_OR2 C2802 ( .A(N1571), .B(m5stg_frac_54_33[33]), .Z(N1572) );
  GTECH_OR2 C2803 ( .A(N1570), .B(m5stg_frac_54_33[34]), .Z(N1571) );
  GTECH_OR2 C2804 ( .A(N1569), .B(m5stg_frac_54_33[35]), .Z(N1570) );
  GTECH_OR2 C2805 ( .A(N1568), .B(m5stg_frac_54_33[36]), .Z(N1569) );
  GTECH_OR2 C2806 ( .A(N1567), .B(m5stg_frac_54_33[37]), .Z(N1568) );
  GTECH_OR2 C2807 ( .A(N1566), .B(m5stg_frac_54_33[38]), .Z(N1567) );
  GTECH_OR2 C2808 ( .A(N1565), .B(m5stg_frac_54_33[39]), .Z(N1566) );
  GTECH_OR2 C2809 ( .A(N1564), .B(m5stg_frac_54_33[40]), .Z(N1565) );
  GTECH_OR2 C2810 ( .A(N1563), .B(m5stg_frac_54_33[41]), .Z(N1564) );
  GTECH_OR2 C2811 ( .A(N1562), .B(m5stg_frac_54_33[42]), .Z(N1563) );
  GTECH_OR2 C2812 ( .A(N1561), .B(m5stg_frac_54_33[43]), .Z(N1562) );
  GTECH_OR2 C2813 ( .A(N1560), .B(m5stg_frac_54_33[44]), .Z(N1561) );
  GTECH_OR2 C2814 ( .A(N1559), .B(m5stg_frac_54_33[45]), .Z(N1560) );
  GTECH_OR2 C2815 ( .A(N1558), .B(m5stg_frac_54_33[46]), .Z(N1559) );
  GTECH_OR2 C2816 ( .A(N1557), .B(m5stg_frac_54_33[47]), .Z(N1558) );
  GTECH_OR2 C2817 ( .A(N1556), .B(m5stg_frac_54_33[48]), .Z(N1557) );
  GTECH_OR2 C2818 ( .A(N1555), .B(m5stg_frac_54_33[49]), .Z(N1556) );
  GTECH_OR2 C2819 ( .A(N1554), .B(m5stg_frac_54_33[50]), .Z(N1555) );
  GTECH_OR2 C2820 ( .A(N1553), .B(m5stg_frac_54_33[51]), .Z(N1554) );
  GTECH_OR2 C2821 ( .A(N1552), .B(m5stg_frac_54_33[52]), .Z(N1553) );
  GTECH_OR2 C2822 ( .A(m5stg_frac_54_33[54]), .B(m5stg_frac_54_33[53]), .Z(
        N1552) );
  GTECH_OR2 C2823 ( .A(N1576), .B(N1577), .Z(mul_frac_out_in[51]) );
  GTECH_OR2 C2824 ( .A(N1574), .B(N1575), .Z(N1576) );
  GTECH_AND2 C2825 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[51]), .Z(
        N1574) );
  GTECH_AND2 C2826 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[54]), .Z(N1575) );
  GTECH_AND2 C2827 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1577) );
  GTECH_OR2 C2828 ( .A(N1580), .B(N1581), .Z(mul_frac_out_in[50]) );
  GTECH_OR2 C2829 ( .A(N1578), .B(N1579), .Z(N1580) );
  GTECH_AND2 C2830 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[50]), .Z(
        N1578) );
  GTECH_AND2 C2831 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[53]), .Z(N1579) );
  GTECH_AND2 C2832 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1581) );
  GTECH_OR2 C2833 ( .A(N1584), .B(N1585), .Z(mul_frac_out_in[49]) );
  GTECH_OR2 C2834 ( .A(N1582), .B(N1583), .Z(N1584) );
  GTECH_AND2 C2835 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[49]), .Z(
        N1582) );
  GTECH_AND2 C2836 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[52]), .Z(N1583) );
  GTECH_AND2 C2837 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1585) );
  GTECH_OR2 C2838 ( .A(N1588), .B(N1589), .Z(mul_frac_out_in[48]) );
  GTECH_OR2 C2839 ( .A(N1586), .B(N1587), .Z(N1588) );
  GTECH_AND2 C2840 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[48]), .Z(
        N1586) );
  GTECH_AND2 C2841 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[51]), .Z(N1587) );
  GTECH_AND2 C2842 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1589) );
  GTECH_OR2 C2843 ( .A(N1592), .B(N1593), .Z(mul_frac_out_in[47]) );
  GTECH_OR2 C2844 ( .A(N1590), .B(N1591), .Z(N1592) );
  GTECH_AND2 C2845 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[47]), .Z(
        N1590) );
  GTECH_AND2 C2846 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[50]), .Z(N1591) );
  GTECH_AND2 C2847 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1593) );
  GTECH_OR2 C2848 ( .A(N1596), .B(N1597), .Z(mul_frac_out_in[46]) );
  GTECH_OR2 C2849 ( .A(N1594), .B(N1595), .Z(N1596) );
  GTECH_AND2 C2850 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[46]), .Z(
        N1594) );
  GTECH_AND2 C2851 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[49]), .Z(N1595) );
  GTECH_AND2 C2852 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1597) );
  GTECH_OR2 C2853 ( .A(N1600), .B(N1601), .Z(mul_frac_out_in[45]) );
  GTECH_OR2 C2854 ( .A(N1598), .B(N1599), .Z(N1600) );
  GTECH_AND2 C2855 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[45]), .Z(
        N1598) );
  GTECH_AND2 C2856 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[48]), .Z(N1599) );
  GTECH_AND2 C2857 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1601) );
  GTECH_OR2 C2858 ( .A(N1604), .B(N1605), .Z(mul_frac_out_in[44]) );
  GTECH_OR2 C2859 ( .A(N1602), .B(N1603), .Z(N1604) );
  GTECH_AND2 C2860 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[44]), .Z(
        N1602) );
  GTECH_AND2 C2861 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[47]), .Z(N1603) );
  GTECH_AND2 C2862 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1605) );
  GTECH_OR2 C2863 ( .A(N1608), .B(N1609), .Z(mul_frac_out_in[43]) );
  GTECH_OR2 C2864 ( .A(N1606), .B(N1607), .Z(N1608) );
  GTECH_AND2 C2865 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[43]), .Z(
        N1606) );
  GTECH_AND2 C2866 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[46]), .Z(N1607) );
  GTECH_AND2 C2867 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1609) );
  GTECH_OR2 C2868 ( .A(N1612), .B(N1613), .Z(mul_frac_out_in[42]) );
  GTECH_OR2 C2869 ( .A(N1610), .B(N1611), .Z(N1612) );
  GTECH_AND2 C2870 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[42]), .Z(
        N1610) );
  GTECH_AND2 C2871 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[45]), .Z(N1611) );
  GTECH_AND2 C2872 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1613) );
  GTECH_OR2 C2873 ( .A(N1616), .B(N1617), .Z(mul_frac_out_in[41]) );
  GTECH_OR2 C2874 ( .A(N1614), .B(N1615), .Z(N1616) );
  GTECH_AND2 C2875 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[41]), .Z(
        N1614) );
  GTECH_AND2 C2876 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[44]), .Z(N1615) );
  GTECH_AND2 C2877 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1617) );
  GTECH_OR2 C2878 ( .A(N1620), .B(N1621), .Z(mul_frac_out_in[40]) );
  GTECH_OR2 C2879 ( .A(N1618), .B(N1619), .Z(N1620) );
  GTECH_AND2 C2880 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[40]), .Z(
        N1618) );
  GTECH_AND2 C2881 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[43]), .Z(N1619) );
  GTECH_AND2 C2882 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1621) );
  GTECH_OR2 C2883 ( .A(N1624), .B(N1625), .Z(mul_frac_out_in[39]) );
  GTECH_OR2 C2884 ( .A(N1622), .B(N1623), .Z(N1624) );
  GTECH_AND2 C2885 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[39]), .Z(
        N1622) );
  GTECH_AND2 C2886 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[42]), .Z(N1623) );
  GTECH_AND2 C2887 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1625) );
  GTECH_OR2 C2888 ( .A(N1628), .B(N1629), .Z(mul_frac_out_in[38]) );
  GTECH_OR2 C2889 ( .A(N1626), .B(N1627), .Z(N1628) );
  GTECH_AND2 C2890 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[38]), .Z(
        N1626) );
  GTECH_AND2 C2891 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[41]), .Z(N1627) );
  GTECH_AND2 C2892 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1629) );
  GTECH_OR2 C2893 ( .A(N1632), .B(N1633), .Z(mul_frac_out_in[37]) );
  GTECH_OR2 C2894 ( .A(N1630), .B(N1631), .Z(N1632) );
  GTECH_AND2 C2895 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[37]), .Z(
        N1630) );
  GTECH_AND2 C2896 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[40]), .Z(N1631) );
  GTECH_AND2 C2897 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1633) );
  GTECH_OR2 C2898 ( .A(N1636), .B(N1637), .Z(mul_frac_out_in[36]) );
  GTECH_OR2 C2899 ( .A(N1634), .B(N1635), .Z(N1636) );
  GTECH_AND2 C2900 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[36]), .Z(
        N1634) );
  GTECH_AND2 C2901 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[39]), .Z(N1635) );
  GTECH_AND2 C2902 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1637) );
  GTECH_OR2 C2903 ( .A(N1640), .B(N1641), .Z(mul_frac_out_in[35]) );
  GTECH_OR2 C2904 ( .A(N1638), .B(N1639), .Z(N1640) );
  GTECH_AND2 C2905 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[35]), .Z(
        N1638) );
  GTECH_AND2 C2906 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[38]), .Z(N1639) );
  GTECH_AND2 C2907 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1641) );
  GTECH_OR2 C2908 ( .A(N1644), .B(N1645), .Z(mul_frac_out_in[34]) );
  GTECH_OR2 C2909 ( .A(N1642), .B(N1643), .Z(N1644) );
  GTECH_AND2 C2910 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[34]), .Z(
        N1642) );
  GTECH_AND2 C2911 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[37]), .Z(N1643) );
  GTECH_AND2 C2912 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1645) );
  GTECH_OR2 C2913 ( .A(N1648), .B(N1649), .Z(mul_frac_out_in[33]) );
  GTECH_OR2 C2914 ( .A(N1646), .B(N1647), .Z(N1648) );
  GTECH_AND2 C2915 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[33]), .Z(
        N1646) );
  GTECH_AND2 C2916 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[36]), .Z(N1647) );
  GTECH_AND2 C2917 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1649) );
  GTECH_OR2 C2918 ( .A(N1652), .B(N1653), .Z(mul_frac_out_in[32]) );
  GTECH_OR2 C2919 ( .A(N1650), .B(N1651), .Z(N1652) );
  GTECH_AND2 C2920 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[32]), .Z(
        N1650) );
  GTECH_AND2 C2921 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[35]), .Z(N1651) );
  GTECH_AND2 C2922 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1653) );
  GTECH_OR2 C2923 ( .A(N1656), .B(N1657), .Z(mul_frac_out_in[31]) );
  GTECH_OR2 C2924 ( .A(N1654), .B(N1655), .Z(N1656) );
  GTECH_AND2 C2925 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[31]), .Z(
        N1654) );
  GTECH_AND2 C2926 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[34]), .Z(N1655) );
  GTECH_AND2 C2927 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1657) );
  GTECH_OR2 C2928 ( .A(N1660), .B(N1661), .Z(mul_frac_out_in[30]) );
  GTECH_OR2 C2929 ( .A(N1658), .B(N1659), .Z(N1660) );
  GTECH_AND2 C2930 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[30]), .Z(
        N1658) );
  GTECH_AND2 C2931 ( .A(mul_frac_out_frac), .B(m5stg_frac_54_33[33]), .Z(N1659) );
  GTECH_AND2 C2932 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1661) );
  GTECH_OR2 C2933 ( .A(N1664), .B(N1665), .Z(mul_frac_out_in[29]) );
  GTECH_OR2 C2934 ( .A(N1662), .B(N1663), .Z(N1664) );
  GTECH_AND2 C2935 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[29]), .Z(
        N1662) );
  GTECH_AND2 C2936 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[32]), .Z(N1663)
         );
  GTECH_AND2 C2937 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1665) );
  GTECH_OR2 C2938 ( .A(N1668), .B(N1669), .Z(mul_frac_out_in[28]) );
  GTECH_OR2 C2939 ( .A(N1666), .B(N1667), .Z(N1668) );
  GTECH_AND2 C2940 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[28]), .Z(
        N1666) );
  GTECH_AND2 C2941 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[31]), .Z(N1667)
         );
  GTECH_AND2 C2942 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1669) );
  GTECH_OR2 C2943 ( .A(N1672), .B(N1673), .Z(mul_frac_out_in[27]) );
  GTECH_OR2 C2944 ( .A(N1670), .B(N1671), .Z(N1672) );
  GTECH_AND2 C2945 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[27]), .Z(
        N1670) );
  GTECH_AND2 C2946 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[30]), .Z(N1671)
         );
  GTECH_AND2 C2947 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1673) );
  GTECH_OR2 C2948 ( .A(N1676), .B(N1677), .Z(mul_frac_out_in[26]) );
  GTECH_OR2 C2949 ( .A(N1674), .B(N1675), .Z(N1676) );
  GTECH_AND2 C2950 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[26]), .Z(
        N1674) );
  GTECH_AND2 C2951 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[29]), .Z(N1675)
         );
  GTECH_AND2 C2952 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1677) );
  GTECH_OR2 C2953 ( .A(N1680), .B(N1681), .Z(mul_frac_out_in[25]) );
  GTECH_OR2 C2954 ( .A(N1678), .B(N1679), .Z(N1680) );
  GTECH_AND2 C2955 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[25]), .Z(
        N1678) );
  GTECH_AND2 C2956 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[28]), .Z(N1679)
         );
  GTECH_AND2 C2957 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1681) );
  GTECH_OR2 C2958 ( .A(N1684), .B(N1685), .Z(mul_frac_out_in[24]) );
  GTECH_OR2 C2959 ( .A(N1682), .B(N1683), .Z(N1684) );
  GTECH_AND2 C2960 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[24]), .Z(
        N1682) );
  GTECH_AND2 C2961 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[27]), .Z(N1683)
         );
  GTECH_AND2 C2962 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1685) );
  GTECH_OR2 C2963 ( .A(N1688), .B(N1689), .Z(mul_frac_out_in[23]) );
  GTECH_OR2 C2964 ( .A(N1686), .B(N1687), .Z(N1688) );
  GTECH_AND2 C2965 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[23]), .Z(
        N1686) );
  GTECH_AND2 C2966 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[26]), .Z(N1687)
         );
  GTECH_AND2 C2967 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1689) );
  GTECH_OR2 C2968 ( .A(N1692), .B(N1693), .Z(mul_frac_out_in[22]) );
  GTECH_OR2 C2969 ( .A(N1690), .B(N1691), .Z(N1692) );
  GTECH_AND2 C2970 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[22]), .Z(
        N1690) );
  GTECH_AND2 C2971 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[25]), .Z(N1691)
         );
  GTECH_AND2 C2972 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1693) );
  GTECH_OR2 C2973 ( .A(N1696), .B(N1697), .Z(mul_frac_out_in[21]) );
  GTECH_OR2 C2974 ( .A(N1694), .B(N1695), .Z(N1696) );
  GTECH_AND2 C2975 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[21]), .Z(
        N1694) );
  GTECH_AND2 C2976 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[24]), .Z(N1695)
         );
  GTECH_AND2 C2977 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1697) );
  GTECH_OR2 C2978 ( .A(N1700), .B(N1701), .Z(mul_frac_out_in[20]) );
  GTECH_OR2 C2979 ( .A(N1698), .B(N1699), .Z(N1700) );
  GTECH_AND2 C2980 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[20]), .Z(
        N1698) );
  GTECH_AND2 C2981 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[23]), .Z(N1699)
         );
  GTECH_AND2 C2982 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1701) );
  GTECH_OR2 C2983 ( .A(N1704), .B(N1705), .Z(mul_frac_out_in[19]) );
  GTECH_OR2 C2984 ( .A(N1702), .B(N1703), .Z(N1704) );
  GTECH_AND2 C2985 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[19]), .Z(
        N1702) );
  GTECH_AND2 C2986 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[22]), .Z(N1703)
         );
  GTECH_AND2 C2987 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1705) );
  GTECH_OR2 C2988 ( .A(N1708), .B(N1709), .Z(mul_frac_out_in[18]) );
  GTECH_OR2 C2989 ( .A(N1706), .B(N1707), .Z(N1708) );
  GTECH_AND2 C2990 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[18]), .Z(
        N1706) );
  GTECH_AND2 C2991 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[21]), .Z(N1707)
         );
  GTECH_AND2 C2992 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1709) );
  GTECH_OR2 C2993 ( .A(N1712), .B(N1713), .Z(mul_frac_out_in[17]) );
  GTECH_OR2 C2994 ( .A(N1710), .B(N1711), .Z(N1712) );
  GTECH_AND2 C2995 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[17]), .Z(
        N1710) );
  GTECH_AND2 C2996 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[20]), .Z(N1711)
         );
  GTECH_AND2 C2997 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1713) );
  GTECH_OR2 C2998 ( .A(N1716), .B(N1717), .Z(mul_frac_out_in[16]) );
  GTECH_OR2 C2999 ( .A(N1714), .B(N1715), .Z(N1716) );
  GTECH_AND2 C3000 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[16]), .Z(
        N1714) );
  GTECH_AND2 C3001 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[19]), .Z(N1715)
         );
  GTECH_AND2 C3002 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1717) );
  GTECH_OR2 C3003 ( .A(N1720), .B(N1721), .Z(mul_frac_out_in[15]) );
  GTECH_OR2 C3004 ( .A(N1718), .B(N1719), .Z(N1720) );
  GTECH_AND2 C3005 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[15]), .Z(
        N1718) );
  GTECH_AND2 C3006 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[18]), .Z(N1719)
         );
  GTECH_AND2 C3007 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1721) );
  GTECH_OR2 C3008 ( .A(N1724), .B(N1725), .Z(mul_frac_out_in[14]) );
  GTECH_OR2 C3009 ( .A(N1722), .B(N1723), .Z(N1724) );
  GTECH_AND2 C3010 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[14]), .Z(
        N1722) );
  GTECH_AND2 C3011 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[17]), .Z(N1723)
         );
  GTECH_AND2 C3012 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1725) );
  GTECH_OR2 C3013 ( .A(N1728), .B(N1729), .Z(mul_frac_out_in[13]) );
  GTECH_OR2 C3014 ( .A(N1726), .B(N1727), .Z(N1728) );
  GTECH_AND2 C3015 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[13]), .Z(
        N1726) );
  GTECH_AND2 C3016 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[16]), .Z(N1727)
         );
  GTECH_AND2 C3017 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1729) );
  GTECH_OR2 C3018 ( .A(N1732), .B(N1733), .Z(mul_frac_out_in[12]) );
  GTECH_OR2 C3019 ( .A(N1730), .B(N1731), .Z(N1732) );
  GTECH_AND2 C3020 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[12]), .Z(
        N1730) );
  GTECH_AND2 C3021 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[15]), .Z(N1731)
         );
  GTECH_AND2 C3022 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1733) );
  GTECH_OR2 C3023 ( .A(N1736), .B(N1737), .Z(mul_frac_out_in[11]) );
  GTECH_OR2 C3024 ( .A(N1734), .B(N1735), .Z(N1736) );
  GTECH_AND2 C3025 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[11]), .Z(
        N1734) );
  GTECH_AND2 C3026 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[14]), .Z(N1735)
         );
  GTECH_AND2 C3027 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1737) );
  GTECH_OR2 C3028 ( .A(N1740), .B(N1741), .Z(mul_frac_out_in[10]) );
  GTECH_OR2 C3029 ( .A(N1738), .B(N1739), .Z(N1740) );
  GTECH_AND2 C3030 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[10]), .Z(
        N1738) );
  GTECH_AND2 C3031 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[13]), .Z(N1739)
         );
  GTECH_AND2 C3032 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1741) );
  GTECH_OR2 C3033 ( .A(N1744), .B(N1745), .Z(mul_frac_out_in[9]) );
  GTECH_OR2 C3034 ( .A(N1742), .B(N1743), .Z(N1744) );
  GTECH_AND2 C3035 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[9]), .Z(
        N1742) );
  GTECH_AND2 C3036 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[12]), .Z(N1743)
         );
  GTECH_AND2 C3037 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1745) );
  GTECH_OR2 C3038 ( .A(N1748), .B(N1749), .Z(mul_frac_out_in[8]) );
  GTECH_OR2 C3039 ( .A(N1746), .B(N1747), .Z(N1748) );
  GTECH_AND2 C3040 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[8]), .Z(
        N1746) );
  GTECH_AND2 C3041 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[11]), .Z(N1747)
         );
  GTECH_AND2 C3042 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1749) );
  GTECH_OR2 C3043 ( .A(N1752), .B(N1753), .Z(mul_frac_out_in[7]) );
  GTECH_OR2 C3044 ( .A(N1750), .B(N1751), .Z(N1752) );
  GTECH_AND2 C3045 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[7]), .Z(
        N1750) );
  GTECH_AND2 C3046 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[10]), .Z(N1751)
         );
  GTECH_AND2 C3047 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1753) );
  GTECH_OR2 C3048 ( .A(N1756), .B(N1757), .Z(mul_frac_out_in[6]) );
  GTECH_OR2 C3049 ( .A(N1754), .B(N1755), .Z(N1756) );
  GTECH_AND2 C3050 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[6]), .Z(
        N1754) );
  GTECH_AND2 C3051 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[9]), .Z(N1755)
         );
  GTECH_AND2 C3052 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1757) );
  GTECH_OR2 C3053 ( .A(N1760), .B(N1761), .Z(mul_frac_out_in[5]) );
  GTECH_OR2 C3054 ( .A(N1758), .B(N1759), .Z(N1760) );
  GTECH_AND2 C3055 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[5]), .Z(
        N1758) );
  GTECH_AND2 C3056 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[8]), .Z(N1759)
         );
  GTECH_AND2 C3057 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1761) );
  GTECH_OR2 C3058 ( .A(N1764), .B(N1765), .Z(mul_frac_out_in[4]) );
  GTECH_OR2 C3059 ( .A(N1762), .B(N1763), .Z(N1764) );
  GTECH_AND2 C3060 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[4]), .Z(
        N1762) );
  GTECH_AND2 C3061 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[7]), .Z(N1763)
         );
  GTECH_AND2 C3062 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1765) );
  GTECH_OR2 C3063 ( .A(N1768), .B(N1769), .Z(mul_frac_out_in[3]) );
  GTECH_OR2 C3064 ( .A(N1766), .B(N1767), .Z(N1768) );
  GTECH_AND2 C3065 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[3]), .Z(
        N1766) );
  GTECH_AND2 C3066 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[6]), .Z(N1767)
         );
  GTECH_AND2 C3067 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1769) );
  GTECH_OR2 C3068 ( .A(N1772), .B(N1773), .Z(mul_frac_out_in[2]) );
  GTECH_OR2 C3069 ( .A(N1770), .B(N1771), .Z(N1772) );
  GTECH_AND2 C3070 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[2]), .Z(
        N1770) );
  GTECH_AND2 C3071 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[5]), .Z(N1771)
         );
  GTECH_AND2 C3072 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1773) );
  GTECH_OR2 C3073 ( .A(N1776), .B(N1777), .Z(mul_frac_out_in[1]) );
  GTECH_OR2 C3074 ( .A(N1774), .B(N1775), .Z(N1776) );
  GTECH_AND2 C3075 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[1]), .Z(
        N1774) );
  GTECH_AND2 C3076 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[4]), .Z(N1775)
         );
  GTECH_AND2 C3077 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1777) );
  GTECH_OR2 C3078 ( .A(N1780), .B(N1781), .Z(mul_frac_out_in[0]) );
  GTECH_OR2 C3079 ( .A(N1778), .B(N1779), .Z(N1780) );
  GTECH_AND2 C3080 ( .A(mul_frac_out_fracadd), .B(m5stg_fracadd_tmp[0]), .Z(
        N1778) );
  GTECH_AND2 C3081 ( .A(mul_frac_out_frac), .B(m5stg_frac_32_0[3]), .Z(N1779)
         );
  GTECH_AND2 C3082 ( .A(m5stg_in_of), .B(m5stg_to_0), .Z(N1781) );
endmodule


module mul_bodec ( x, b, b0, b1, b2, b3, b4, b5, b6, b7 );
  input [15:0] b;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  input x;
  wire   b_12, b_10, b_8, b_6, b_4, b_2, b_0, N0, N1, N2, N3, N4, N5, N6, N7,
         N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88;
  assign b_12 = b[12];
  assign b_10 = b[10];
  assign b_8 = b[8];
  assign b_6 = b[6];
  assign b_4 = b[4];
  assign b_2 = b[2];
  assign b_0 = b[0];
  assign b0[2] = b[1];
  assign b1[2] = b[3];
  assign b2[2] = b[5];
  assign b3[2] = b[7];
  assign b4[2] = b[9];
  assign b5[2] = b[11];
  assign b6[2] = b[13];
  assign b7[2] = b[15];

  GTECH_NOT I_0 ( .A(N7), .Z(b0[1]) );
  GTECH_OR2 C23 ( .A(N1), .B(N6), .Z(N7) );
  GTECH_AND2 C24 ( .A(N0), .B(x), .Z(N1) );
  GTECH_AND2 C25 ( .A(b0[2]), .B(b_0), .Z(N0) );
  GTECH_AND2 C26 ( .A(N4), .B(N5), .Z(N6) );
  GTECH_AND2 C27 ( .A(N2), .B(N3), .Z(N4) );
  GTECH_NOT I_1 ( .A(b0[2]), .Z(N2) );
  GTECH_NOT I_2 ( .A(b_0), .Z(N3) );
  GTECH_NOT I_3 ( .A(x), .Z(N5) );
  GTECH_OR2 C31 ( .A(N9), .B(N11), .Z(b0[0]) );
  GTECH_AND2 C32 ( .A(N8), .B(x), .Z(N9) );
  GTECH_AND2 C33 ( .A(N2), .B(b_0), .Z(N8) );
  GTECH_AND2 C35 ( .A(N10), .B(N5), .Z(N11) );
  GTECH_AND2 C36 ( .A(b0[2]), .B(N3), .Z(N10) );
  GTECH_NOT I_4 ( .A(N18), .Z(b1[1]) );
  GTECH_OR2 C40 ( .A(N13), .B(N17), .Z(N18) );
  GTECH_AND2 C41 ( .A(N12), .B(b0[2]), .Z(N13) );
  GTECH_AND2 C42 ( .A(b1[2]), .B(b_2), .Z(N12) );
  GTECH_AND2 C43 ( .A(N16), .B(N2), .Z(N17) );
  GTECH_AND2 C44 ( .A(N14), .B(N15), .Z(N16) );
  GTECH_NOT I_5 ( .A(b1[2]), .Z(N14) );
  GTECH_NOT I_6 ( .A(b_2), .Z(N15) );
  GTECH_OR2 C48 ( .A(N20), .B(N22), .Z(b1[0]) );
  GTECH_AND2 C49 ( .A(N19), .B(b0[2]), .Z(N20) );
  GTECH_AND2 C50 ( .A(N14), .B(b_2), .Z(N19) );
  GTECH_AND2 C52 ( .A(N21), .B(N2), .Z(N22) );
  GTECH_AND2 C53 ( .A(b1[2]), .B(N15), .Z(N21) );
  GTECH_NOT I_7 ( .A(N29), .Z(b2[1]) );
  GTECH_OR2 C57 ( .A(N24), .B(N28), .Z(N29) );
  GTECH_AND2 C58 ( .A(N23), .B(b1[2]), .Z(N24) );
  GTECH_AND2 C59 ( .A(b2[2]), .B(b_4), .Z(N23) );
  GTECH_AND2 C60 ( .A(N27), .B(N14), .Z(N28) );
  GTECH_AND2 C61 ( .A(N25), .B(N26), .Z(N27) );
  GTECH_NOT I_8 ( .A(b2[2]), .Z(N25) );
  GTECH_NOT I_9 ( .A(b_4), .Z(N26) );
  GTECH_OR2 C65 ( .A(N31), .B(N33), .Z(b2[0]) );
  GTECH_AND2 C66 ( .A(N30), .B(b1[2]), .Z(N31) );
  GTECH_AND2 C67 ( .A(N25), .B(b_4), .Z(N30) );
  GTECH_AND2 C69 ( .A(N32), .B(N14), .Z(N33) );
  GTECH_AND2 C70 ( .A(b2[2]), .B(N26), .Z(N32) );
  GTECH_NOT I_10 ( .A(N40), .Z(b3[1]) );
  GTECH_OR2 C74 ( .A(N35), .B(N39), .Z(N40) );
  GTECH_AND2 C75 ( .A(N34), .B(b2[2]), .Z(N35) );
  GTECH_AND2 C76 ( .A(b3[2]), .B(b_6), .Z(N34) );
  GTECH_AND2 C77 ( .A(N38), .B(N25), .Z(N39) );
  GTECH_AND2 C78 ( .A(N36), .B(N37), .Z(N38) );
  GTECH_NOT I_11 ( .A(b3[2]), .Z(N36) );
  GTECH_NOT I_12 ( .A(b_6), .Z(N37) );
  GTECH_OR2 C82 ( .A(N42), .B(N44), .Z(b3[0]) );
  GTECH_AND2 C83 ( .A(N41), .B(b2[2]), .Z(N42) );
  GTECH_AND2 C84 ( .A(N36), .B(b_6), .Z(N41) );
  GTECH_AND2 C86 ( .A(N43), .B(N25), .Z(N44) );
  GTECH_AND2 C87 ( .A(b3[2]), .B(N37), .Z(N43) );
  GTECH_NOT I_13 ( .A(N51), .Z(b4[1]) );
  GTECH_OR2 C91 ( .A(N46), .B(N50), .Z(N51) );
  GTECH_AND2 C92 ( .A(N45), .B(b3[2]), .Z(N46) );
  GTECH_AND2 C93 ( .A(b4[2]), .B(b_8), .Z(N45) );
  GTECH_AND2 C94 ( .A(N49), .B(N36), .Z(N50) );
  GTECH_AND2 C95 ( .A(N47), .B(N48), .Z(N49) );
  GTECH_NOT I_14 ( .A(b4[2]), .Z(N47) );
  GTECH_NOT I_15 ( .A(b_8), .Z(N48) );
  GTECH_OR2 C99 ( .A(N53), .B(N55), .Z(b4[0]) );
  GTECH_AND2 C100 ( .A(N52), .B(b3[2]), .Z(N53) );
  GTECH_AND2 C101 ( .A(N47), .B(b_8), .Z(N52) );
  GTECH_AND2 C103 ( .A(N54), .B(N36), .Z(N55) );
  GTECH_AND2 C104 ( .A(b4[2]), .B(N48), .Z(N54) );
  GTECH_NOT I_16 ( .A(N62), .Z(b5[1]) );
  GTECH_OR2 C108 ( .A(N57), .B(N61), .Z(N62) );
  GTECH_AND2 C109 ( .A(N56), .B(b4[2]), .Z(N57) );
  GTECH_AND2 C110 ( .A(b5[2]), .B(b_10), .Z(N56) );
  GTECH_AND2 C111 ( .A(N60), .B(N47), .Z(N61) );
  GTECH_AND2 C112 ( .A(N58), .B(N59), .Z(N60) );
  GTECH_NOT I_17 ( .A(b5[2]), .Z(N58) );
  GTECH_NOT I_18 ( .A(b_10), .Z(N59) );
  GTECH_OR2 C116 ( .A(N64), .B(N66), .Z(b5[0]) );
  GTECH_AND2 C117 ( .A(N63), .B(b4[2]), .Z(N64) );
  GTECH_AND2 C118 ( .A(N58), .B(b_10), .Z(N63) );
  GTECH_AND2 C120 ( .A(N65), .B(N47), .Z(N66) );
  GTECH_AND2 C121 ( .A(b5[2]), .B(N59), .Z(N65) );
  GTECH_NOT I_19 ( .A(N73), .Z(b6[1]) );
  GTECH_OR2 C125 ( .A(N68), .B(N72), .Z(N73) );
  GTECH_AND2 C126 ( .A(N67), .B(b5[2]), .Z(N68) );
  GTECH_AND2 C127 ( .A(b6[2]), .B(b_12), .Z(N67) );
  GTECH_AND2 C128 ( .A(N71), .B(N58), .Z(N72) );
  GTECH_AND2 C129 ( .A(N69), .B(N70), .Z(N71) );
  GTECH_NOT I_20 ( .A(b6[2]), .Z(N69) );
  GTECH_NOT I_21 ( .A(b_12), .Z(N70) );
  GTECH_OR2 C133 ( .A(N75), .B(N77), .Z(b6[0]) );
  GTECH_AND2 C134 ( .A(N74), .B(b5[2]), .Z(N75) );
  GTECH_AND2 C135 ( .A(N69), .B(b_12), .Z(N74) );
  GTECH_AND2 C137 ( .A(N76), .B(N58), .Z(N77) );
  GTECH_AND2 C138 ( .A(b6[2]), .B(N70), .Z(N76) );
  GTECH_NOT I_22 ( .A(N84), .Z(b7[1]) );
  GTECH_OR2 C142 ( .A(N79), .B(N83), .Z(N84) );
  GTECH_AND2 C143 ( .A(N78), .B(b6[2]), .Z(N79) );
  GTECH_AND2 C144 ( .A(b7[2]), .B(b[14]), .Z(N78) );
  GTECH_AND2 C145 ( .A(N82), .B(N69), .Z(N83) );
  GTECH_AND2 C146 ( .A(N80), .B(N81), .Z(N82) );
  GTECH_NOT I_23 ( .A(b7[2]), .Z(N80) );
  GTECH_NOT I_24 ( .A(b[14]), .Z(N81) );
  GTECH_OR2 C150 ( .A(N86), .B(N88), .Z(b7[0]) );
  GTECH_AND2 C151 ( .A(N85), .B(b6[2]), .Z(N86) );
  GTECH_AND2 C152 ( .A(N80), .B(b[14]), .Z(N85) );
  GTECH_AND2 C154 ( .A(N87), .B(N69), .Z(N88) );
  GTECH_AND2 C155 ( .A(b7[2]), .B(N81), .Z(N87) );
endmodule


module dff_SIZE32 ( din, clk, q, se, si, so );
  input [31:0] din;
  output [31:0] q;
  input [31:0] si;
  output [31:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34;
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C42 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, 
        N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, 
        N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dp_mux2es_SIZE3 ( dout, in0, in1, sel );
  output [2:0] dout;
  input [2:0] in0;
  input [2:0] in1;
  input sel;
  wire   N0, N1, N2;

  SELECT_OP C13 ( .DATA1(in1), .DATA2(in0), .CONTROL1(N0), .CONTROL2(N1), .Z(
        dout) );
  GTECH_BUF B_0 ( .A(sel), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(sel), .Z(N2) );
endmodule


module dp_mux2es ( dout, in0, in1, sel );
  output [0:0] dout;
  input [0:0] in0;
  input [0:0] in1;
  input sel;
  wire   N0, N1, N2;

  SELECT_OP C11 ( .DATA1(in1[0]), .DATA2(in0[0]), .CONTROL1(N0), .CONTROL2(N1), 
        .Z(dout[0]) );
  GTECH_BUF B_0 ( .A(sel), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(sel), .Z(N2) );
endmodule


module dff_SIZE3 ( din, clk, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5;
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C13 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module mul_booth ( head, b_in, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, 
        b11, b12, b13, b14, b15, b16, clk, se, si, so, mul_step, tm_l );
  input [63:0] b_in;
  output [2:0] b0;
  output [2:0] b1;
  output [2:0] b2;
  output [2:0] b3;
  output [2:0] b4;
  output [2:0] b5;
  output [2:0] b6;
  output [2:0] b7;
  output [2:0] b8;
  output [2:0] b9;
  output [2:0] b10;
  output [2:0] b11;
  output [2:0] b12;
  output [2:0] b13;
  output [2:0] b14;
  output [2:0] b15;
  input head, clk, se, si, mul_step, tm_l;
  output b16, so;
  wire   clk_enb0, _1_net_, clk_enb1, _2_net_, _3_net_, _4_net_, _5_net_,
         _6_net_, _7_net_, _8_net_, _9_net_, _10_net_, _11_net_, _12_net_,
         _13_net_, _14_net_, _15_net_, _16_net_, _17_net_, _18_net_, b16_outmx,
         _20_net_, N0, net12126, net12127, net12128, net12129, net12130,
         net12131, net12132, net12133, net12134, net12135, net12136, net12137,
         net12138, net12139, net12140, net12141, net12142, net12143, net12144,
         net12145, net12146, net12147, net12148, net12149, net12150, net12151,
         net12152, net12153, net12154, net12155, net12156, net12157, net12158,
         net12159, net12160, net12161, net12162, net12163, net12164, net12165,
         net12166, net12167, net12168, net12169, net12170, net12171, net12172,
         net12173, net12174, net12175, net12176, net12177, net12178, net12179,
         net12180, net12181, net12182, net12183, net12184, net12185, net12186,
         net12187, net12188, net12189, net12190, net12191, net12192, net12193,
         net12194, net12195, net12196, net12197, net12198, net12199, net12200,
         net12201, net12202, net12203, net12204, net12205, net12206, net12207;
  wire   [2:0] b0_in0;
  wire   [2:0] b1_in0;
  wire   [2:0] b2_in0;
  wire   [2:0] b3_in0;
  wire   [2:0] b4_in0;
  wire   [2:0] b5_in0;
  wire   [2:0] b6_in0;
  wire   [2:0] b7_in0;
  wire   [2:0] b8_in0;
  wire   [2:0] b9_in0;
  wire   [2:0] b10_in0;
  wire   [2:0] b11_in0;
  wire   [2:0] b12_in0;
  wire   [2:0] b13_in0;
  wire   [2:0] b14_in0;
  wire   [2:0] b15_in0;
  wire   [63:31] b;
  wire   [2:0] b0_in1;
  wire   [2:0] b1_in1;
  wire   [2:0] b2_in1;
  wire   [2:0] b3_in1;
  wire   [2:0] b4_in1;
  wire   [2:0] b5_in1;
  wire   [2:0] b6_in1;
  wire   [2:0] b7_in1;
  wire   [2:0] b8_in1;
  wire   [2:0] b9_in1;
  wire   [2:0] b10_in1;
  wire   [2:0] b11_in1;
  wire   [2:0] b12_in1;
  wire   [2:0] b13_in1;
  wire   [2:0] b14_in1;
  wire   [2:0] b15_in1;
  wire   [2:0] b0_outmx;
  wire   [2:0] b1_outmx;
  wire   [2:0] b2_outmx;
  wire   [2:0] b3_outmx;
  wire   [2:0] b4_outmx;
  wire   [2:0] b5_outmx;
  wire   [2:0] b6_outmx;
  wire   [2:0] b7_outmx;
  wire   [2:0] b8_outmx;
  wire   [2:0] b9_outmx;
  wire   [2:0] b10_outmx;
  wire   [2:0] b11_outmx;
  wire   [2:0] b12_outmx;
  wire   [2:0] b13_outmx;
  wire   [2:0] b14_outmx;
  wire   [2:0] b15_outmx;

  mul_bodec encode0_a ( .x(1'b0), .b(b_in[15:0]), .b0(b0_in0), .b1(b1_in0), 
        .b2(b2_in0), .b3(b3_in0), .b4(b4_in0), .b5(b5_in0), .b6(b6_in0), .b7(
        b7_in0) );
  mul_bodec encode0_b ( .x(b_in[15]), .b(b_in[31:16]), .b0(b8_in0), .b1(b9_in0), .b2(b10_in0), .b3(b11_in0), .b4(b12_in0), .b5(b13_in0), .b6(b14_in0), .b7(
        b15_in0) );
  clken_buf ckbuf_0 ( .clk(clk_enb0), .rclk(clk), .enb_l(_1_net_), .tmb_l(tm_l) );
  clken_buf ckbuf_1 ( .clk(clk_enb1), .rclk(clk), .enb_l(_2_net_), .tmb_l(tm_l) );
  dff_SIZE1 hld_dff0 ( .din(b_in[31]), .clk(clk_enb1), .q(b[31]), .se(se), 
        .si(net12207) );
  dff_SIZE32 hld_dff ( .din(b_in[63:32]), .clk(clk_enb1), .q(b[63:32]), .se(se), .si({net12175, net12176, net12177, net12178, net12179, net12180, net12181, 
        net12182, net12183, net12184, net12185, net12186, net12187, net12188, 
        net12189, net12190, net12191, net12192, net12193, net12194, net12195, 
        net12196, net12197, net12198, net12199, net12200, net12201, net12202, 
        net12203, net12204, net12205, net12206}) );
  mul_bodec encode1_a ( .x(b[31]), .b(b[47:32]), .b0(b0_in1), .b1(b1_in1), 
        .b2(b2_in1), .b3(b3_in1), .b4(b4_in1), .b5(b5_in1), .b6(b6_in1), .b7(
        b7_in1) );
  mul_bodec encode1_b ( .x(b[47]), .b(b[63:48]), .b0(b8_in1), .b1(b9_in1), 
        .b2(b10_in1), .b3(b11_in1), .b4(b12_in1), .b5(b13_in1), .b6(b14_in1), 
        .b7(b15_in1) );
  dp_mux2es_SIZE3 out_mux0 ( .dout(b0_outmx), .in0(b0_in0), .in1(b0_in1), 
        .sel(_3_net_) );
  dp_mux2es_SIZE3 out_mux1 ( .dout(b1_outmx), .in0(b1_in0), .in1(b1_in1), 
        .sel(_4_net_) );
  dp_mux2es_SIZE3 out_mux2 ( .dout(b2_outmx), .in0(b2_in0), .in1(b2_in1), 
        .sel(_5_net_) );
  dp_mux2es_SIZE3 out_mux3 ( .dout(b3_outmx), .in0(b3_in0), .in1(b3_in1), 
        .sel(_6_net_) );
  dp_mux2es_SIZE3 out_mux4 ( .dout(b4_outmx), .in0(b4_in0), .in1(b4_in1), 
        .sel(_7_net_) );
  dp_mux2es_SIZE3 out_mux5 ( .dout(b5_outmx), .in0(b5_in0), .in1(b5_in1), 
        .sel(_8_net_) );
  dp_mux2es_SIZE3 out_mux6 ( .dout(b6_outmx), .in0(b6_in0), .in1(b6_in1), 
        .sel(_9_net_) );
  dp_mux2es_SIZE3 out_mux7 ( .dout(b7_outmx), .in0(b7_in0), .in1(b7_in1), 
        .sel(_10_net_) );
  dp_mux2es_SIZE3 out_mux8 ( .dout(b8_outmx), .in0(b8_in0), .in1(b8_in1), 
        .sel(_11_net_) );
  dp_mux2es_SIZE3 out_mux9 ( .dout(b9_outmx), .in0(b9_in0), .in1(b9_in1), 
        .sel(_12_net_) );
  dp_mux2es_SIZE3 out_mux10 ( .dout(b10_outmx), .in0(b10_in0), .in1(b10_in1), 
        .sel(_13_net_) );
  dp_mux2es_SIZE3 out_mux11 ( .dout(b11_outmx), .in0(b11_in0), .in1(b11_in1), 
        .sel(_14_net_) );
  dp_mux2es_SIZE3 out_mux12 ( .dout(b12_outmx), .in0(b12_in0), .in1(b12_in1), 
        .sel(_15_net_) );
  dp_mux2es_SIZE3 out_mux13 ( .dout(b13_outmx), .in0(b13_in0), .in1(b13_in1), 
        .sel(_16_net_) );
  dp_mux2es_SIZE3 out_mux14 ( .dout(b14_outmx), .in0(b14_in0), .in1(b14_in1), 
        .sel(_17_net_) );
  dp_mux2es_SIZE3 out_mux15 ( .dout(b15_outmx), .in0(b15_in0), .in1(b15_in1), 
        .sel(_18_net_) );
  dp_mux2es out_mux16 ( .dout(b16_outmx), .in0(1'b0), .in1(b[63]), .sel(
        _20_net_) );
  dff_SIZE3 out_dff0 ( .din(b0_outmx), .clk(clk_enb0), .q(b0), .se(se), .si({
        net12172, net12173, net12174}) );
  dff_SIZE3 out_dff1 ( .din(b1_outmx), .clk(clk_enb0), .q(b1), .se(se), .si({
        net12169, net12170, net12171}) );
  dff_SIZE3 out_dff2 ( .din(b2_outmx), .clk(clk_enb0), .q(b2), .se(se), .si({
        net12166, net12167, net12168}) );
  dff_SIZE3 out_dff3 ( .din(b3_outmx), .clk(clk_enb0), .q(b3), .se(se), .si({
        net12163, net12164, net12165}) );
  dff_SIZE3 out_dff4 ( .din(b4_outmx), .clk(clk_enb0), .q(b4), .se(se), .si({
        net12160, net12161, net12162}) );
  dff_SIZE3 out_dff5 ( .din(b5_outmx), .clk(clk_enb0), .q(b5), .se(se), .si({
        net12157, net12158, net12159}) );
  dff_SIZE3 out_dff6 ( .din(b6_outmx), .clk(clk_enb0), .q(b6), .se(se), .si({
        net12154, net12155, net12156}) );
  dff_SIZE3 out_dff7 ( .din(b7_outmx), .clk(clk_enb0), .q(b7), .se(se), .si({
        net12151, net12152, net12153}) );
  dff_SIZE3 out_dff8 ( .din(b8_outmx), .clk(clk_enb0), .q(b8), .se(se), .si({
        net12148, net12149, net12150}) );
  dff_SIZE3 out_dff9 ( .din(b9_outmx), .clk(clk_enb0), .q(b9), .se(se), .si({
        net12145, net12146, net12147}) );
  dff_SIZE3 out_dff10 ( .din(b10_outmx), .clk(clk_enb0), .q(b10), .se(se), 
        .si({net12142, net12143, net12144}) );
  dff_SIZE3 out_dff11 ( .din(b11_outmx), .clk(clk_enb0), .q(b11), .se(se), 
        .si({net12139, net12140, net12141}) );
  dff_SIZE3 out_dff12 ( .din(b12_outmx), .clk(clk_enb0), .q(b12), .se(se), 
        .si({net12136, net12137, net12138}) );
  dff_SIZE3 out_dff13 ( .din(b13_outmx), .clk(clk_enb0), .q(b13), .se(se), 
        .si({net12133, net12134, net12135}) );
  dff_SIZE3 out_dff14 ( .din(b14_outmx), .clk(clk_enb0), .q(b14), .se(se), 
        .si({net12130, net12131, net12132}) );
  dff_SIZE3 out_dff15 ( .din(b15_outmx), .clk(clk_enb0), .q(b15), .se(se), 
        .si({net12127, net12128, net12129}) );
  dff_SIZE1 out_dff16 ( .din(b16_outmx), .clk(clk_enb0), .q(b16), .se(se), 
        .si(net12126) );
  GTECH_NOT I_0 ( .A(mul_step), .Z(_1_net_) );
  GTECH_NOT I_1 ( .A(N0), .Z(_2_net_) );
  GTECH_AND2 C28 ( .A(head), .B(mul_step), .Z(N0) );
  GTECH_NOT I_2 ( .A(head), .Z(_3_net_) );
  GTECH_NOT I_3 ( .A(head), .Z(_4_net_) );
  GTECH_NOT I_4 ( .A(head), .Z(_5_net_) );
  GTECH_NOT I_5 ( .A(head), .Z(_6_net_) );
  GTECH_NOT I_6 ( .A(head), .Z(_7_net_) );
  GTECH_NOT I_7 ( .A(head), .Z(_8_net_) );
  GTECH_NOT I_8 ( .A(head), .Z(_9_net_) );
  GTECH_NOT I_9 ( .A(head), .Z(_10_net_) );
  GTECH_NOT I_10 ( .A(head), .Z(_11_net_) );
  GTECH_NOT I_11 ( .A(head), .Z(_12_net_) );
  GTECH_NOT I_12 ( .A(head), .Z(_13_net_) );
  GTECH_NOT I_13 ( .A(head), .Z(_14_net_) );
  GTECH_NOT I_14 ( .A(head), .Z(_15_net_) );
  GTECH_NOT I_15 ( .A(head), .Z(_16_net_) );
  GTECH_NOT I_16 ( .A(head), .Z(_17_net_) );
  GTECH_NOT I_17 ( .A(head), .Z(_18_net_) );
  GTECH_NOT I_18 ( .A(head), .Z(_20_net_) );
endmodule


module mul_negen ( n0, n1, b );
  input [2:0] b;
  output n0, n1;
  wire   N0, N1, N2;

  GTECH_AND2 C8 ( .A(N0), .B(N1), .Z(n0) );
  GTECH_AND2 C9 ( .A(b[2]), .B(b[1]), .Z(N0) );
  GTECH_NOT I_0 ( .A(b[0]), .Z(N1) );
  GTECH_AND2 C11 ( .A(N2), .B(b[0]), .Z(n1) );
  GTECH_AND2 C12 ( .A(b[2]), .B(b[1]), .Z(N2) );
endmodule


module mul_csa42 ( sum, carry, cout, a, b, c, d, cin );
  input a, b, c, d, cin;
  output sum, carry, cout;
  wire   x, y, z, N0, N1, N2, N3, N4, N5;

  GTECH_XOR2 C12 ( .A(a), .B(b), .Z(x) );
  GTECH_XOR2 C13 ( .A(c), .B(d), .Z(y) );
  GTECH_XOR2 C14 ( .A(x), .B(y), .Z(z) );
  GTECH_XOR2 C15 ( .A(z), .B(cin), .Z(sum) );
  GTECH_OR2 C16 ( .A(N1), .B(N2), .Z(carry) );
  GTECH_AND2 C17 ( .A(b), .B(N0), .Z(N1) );
  GTECH_NOT I_0 ( .A(z), .Z(N0) );
  GTECH_AND2 C19 ( .A(cin), .B(z), .Z(N2) );
  GTECH_OR2 C20 ( .A(N4), .B(N5), .Z(cout) );
  GTECH_AND2 C21 ( .A(d), .B(N3), .Z(N4) );
  GTECH_NOT I_1 ( .A(y), .Z(N3) );
  GTECH_AND2 C23 ( .A(a), .B(y), .Z(N5) );
endmodule


module mul_csa32 ( sum, cout, a, b, c );
  input a, b, c;
  output sum, cout;
  wire   x, y0, y1, y2, N0;

  GTECH_XOR2 C12 ( .A(a), .B(b), .Z(x) );
  GTECH_XOR2 C13 ( .A(c), .B(x), .Z(sum) );
  GTECH_AND2 C14 ( .A(a), .B(b), .Z(y0) );
  GTECH_AND2 C15 ( .A(a), .B(c), .Z(y1) );
  GTECH_AND2 C16 ( .A(b), .B(c), .Z(y2) );
  GTECH_OR2 C17 ( .A(N0), .B(y2), .Z(cout) );
  GTECH_OR2 C18 ( .A(y0), .B(y1), .Z(N0) );
endmodule


module mul_ha ( cout, sum, a, b );
  input a, b;
  output cout, sum;


  GTECH_XOR2 C8 ( .A(a), .B(b), .Z(sum) );
  GTECH_AND2 C9 ( .A(a), .B(b), .Z(cout) );
endmodule


module mul_ppgensign ( p_l, z, b, pm1_l );
  input [2:0] b;
  input pm1_l;
  output p_l, z;
  wire   N0, N1, N2, N3, N4;

  SELECT_OP C14 ( .DATA1(N2), .DATA2(N3), .CONTROL1(N0), .CONTROL2(N1), .Z(z)
         );
  GTECH_BUF B_0 ( .A(b[0]), .Z(N0) );
  GTECH_NOT I_0 ( .A(N4), .Z(p_l) );
  GTECH_AND2 C17 ( .A(b[1]), .B(b[2]), .Z(N4) );
  GTECH_NOT I_1 ( .A(b[0]), .Z(N1) );
  GTECH_NOT I_2 ( .A(pm1_l), .Z(N2) );
  GTECH_NOT I_3 ( .A(p_l), .Z(N3) );
endmodule


module mul_ppgen ( p_l, z, a, b, pm1_l );
  input [2:0] b;
  input a, pm1_l;
  output p_l, z;
  wire   N0, N1, N2, N3, N4, N5;

  SELECT_OP C14 ( .DATA1(N2), .DATA2(N3), .CONTROL1(N0), .CONTROL2(N1), .Z(z)
         );
  GTECH_BUF B_0 ( .A(b[0]), .Z(N0) );
  GTECH_NOT I_0 ( .A(N5), .Z(p_l) );
  GTECH_AND2 C17 ( .A(N4), .B(b[1]), .Z(N5) );
  GTECH_XOR2 C18 ( .A(a), .B(b[2]), .Z(N4) );
  GTECH_NOT I_1 ( .A(b[0]), .Z(N1) );
  GTECH_NOT I_2 ( .A(pm1_l), .Z(N2) );
  GTECH_NOT I_3 ( .A(p_l), .Z(N3) );
endmodule


module mul_ppgen3sign ( cout, sum, am1, am2, am3, am4, b0, b1, b2, bot, head, 
        p0m1_l, p1m1_l, p2m1_l );
  output [4:0] cout;
  output [5:0] sum;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am1, am2, am3, am4, bot, head, p0m1_l, p1m1_l, p2m1_l;
  wire   net075, net088, net0117, net37, net42, net47, p2_l_67, net073,
         p1_l_65, net38, net0118, p2_l_66, net078, p2_l_65, net8, p2_l_64,
         net15, p1_l_64, net43, net48, net35;

  mul_ppgensign p0_64_ ( .p_l(net088), .z(net47), .b(b0), .pm1_l(p0m1_l) );
  mul_ppgensign p2_68_ ( .p_l(net075), .z(net073), .b(b2), .pm1_l(p2_l_67) );
  mul_ppgensign p1_66_ ( .p_l(net0118), .z(net38), .b(b1), .pm1_l(p1_l_65) );
  mul_ha sc1_68_ ( .cout(cout[4]), .sum(sum[4]), .a(1'b1), .b(net073) );
  mul_ppgen p2_67_ ( .p_l(p2_l_67), .z(net078), .a(am1), .b(b2), .pm1_l(
        p2_l_66) );
  mul_ppgen p2_66_ ( .p_l(p2_l_66), .z(net8), .a(am2), .b(b2), .pm1_l(p2_l_65)
         );
  mul_ppgen p2_65_ ( .p_l(p2_l_65), .z(net15), .a(am3), .b(b2), .pm1_l(p2_l_64) );
  mul_ppgen p1_65_ ( .p_l(p1_l_65), .z(net43), .a(am1), .b(b1), .pm1_l(p1_l_64) );
  mul_ppgen p1_64_ ( .p_l(p1_l_64), .z(net48), .a(am2), .b(b1), .pm1_l(p1m1_l)
         );
  mul_ppgen p2_64_ ( .p_l(p2_l_64), .z(net35), .a(am4), .b(b2), .pm1_l(p2m1_l)
         );
  mul_csa32 sc1_67_ ( .sum(sum[3]), .cout(cout[3]), .a(net0118), .b(net0117), 
        .c(net078) );
  mul_csa32 sc1_66_ ( .sum(sum[2]), .cout(cout[2]), .a(net38), .b(net37), .c(
        net8) );
  mul_csa32 sc1_65_ ( .sum(sum[1]), .cout(cout[1]), .a(net43), .b(net42), .c(
        net15) );
  mul_csa32 sc1_64_ ( .sum(sum[0]), .cout(cout[0]), .a(net48), .b(net47), .c(
        net35) );
  GTECH_AND2 C10 ( .A(bot), .B(net075), .Z(sum[5]) );
  GTECH_AND2 C11 ( .A(head), .B(net088), .Z(net0117) );
  GTECH_NOT I_0 ( .A(net0117), .Z(net37) );
  GTECH_XOR2 C13 ( .A(head), .B(net088), .Z(net42) );
endmodule


module mul_ppgen3 ( cout, p0_l, p1_l, p2_l, sum, am2, am4, a, b0, b1, b2, 
        p0m1_l, p1m1_l, p2m1_l );
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input am2, am4, a, p0m1_l, p1m1_l, p2m1_l;
  output cout, p0_l, p1_l, p2_l, sum;
  wire   net046, net32, net043;

  mul_csa32 sc1 ( .sum(sum), .cout(cout), .a(net046), .b(net32), .c(net043) );
  mul_ppgen p2 ( .p_l(p2_l), .z(net043), .a(am4), .b(b2), .pm1_l(p2m1_l) );
  mul_ppgen p1 ( .p_l(p1_l), .z(net046), .a(am2), .b(b1), .pm1_l(p1m1_l) );
  mul_ppgen p0 ( .p_l(p0_l), .z(net32), .a(a), .b(b0), .pm1_l(p0m1_l) );
endmodule


module mul_ppgen3lsb4 ( cout, p0_l, p1_l, sum, a, b0, b1 );
  output [3:1] cout;
  output [3:0] sum;
  input [3:0] a;
  input [2:0] b0;
  input [2:0] b1;
  output p0_l, p1_l;
  wire   b0n_1, b0n_0, p0_0, b0n, b1n_1, b1n_0, p0_2, p1_2, p0_3, p1_3, p0_1,
         p0_l_2, p1_l_2, p0_l_1, p0_l_0, N0;

  mul_negen p0n ( .n0(b0n_0), .n1(b0n_1), .b(b0) );
  mul_negen p1n ( .n0(b1n_0), .n1(b1n_1), .b(b1) );
  mul_csa32 sc1_2_ ( .sum(sum[2]), .cout(cout[2]), .a(p0_2), .b(p1_2), .c(
        b1n_0) );
  mul_csa32 sc1_3_ ( .sum(sum[3]), .cout(cout[3]), .a(p0_3), .b(p1_3), .c(
        b1n_1) );
  mul_ha sc1_1_ ( .cout(cout[1]), .sum(sum[1]), .a(p0_1), .b(b0n) );
  mul_ppgen p0_3_ ( .p_l(p0_l), .z(p0_3), .a(a[3]), .b(b0), .pm1_l(p0_l_2) );
  mul_ppgen p1_3_ ( .p_l(p1_l), .z(p1_3), .a(a[1]), .b(b1), .pm1_l(p1_l_2) );
  mul_ppgen p0_2_ ( .p_l(p0_l_2), .z(p0_2), .a(a[2]), .b(b0), .pm1_l(p0_l_1)
         );
  mul_ppgen p0_1_ ( .p_l(p0_l_1), .z(p0_1), .a(a[1]), .b(b0), .pm1_l(p0_l_0)
         );
  mul_ppgen p0_0_ ( .p_l(p0_l_0), .z(p0_0), .a(a[0]), .b(b0), .pm1_l(1'b1) );
  mul_ppgen p1_2_ ( .p_l(p1_l_2), .z(p1_2), .a(a[0]), .b(b1), .pm1_l(1'b1) );
  GTECH_OR2 C8 ( .A(b0n_1), .B(N0), .Z(b0n) );
  GTECH_AND2 C9 ( .A(b0n_0), .B(p0_0), .Z(N0) );
  GTECH_XOR2 C10 ( .A(b0n_0), .B(p0_0), .Z(sum[0]) );
endmodule


module mul_ppgenrow3 ( cout, sum, a, b0, b1, b2, bot, head );
  output [68:1] cout;
  output [69:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input bot, head;

  wire   [63:4] p2_l;
  wire   [63:3] p1_l;
  wire   [63:3] p0_l;

  mul_ppgen3sign I2 ( .cout(cout[68:64]), .sum(sum[69:64]), .am1(a[63]), .am2(
        a[62]), .am3(a[61]), .am4(a[60]), .b0(b0), .b1(b1), .b2(b2), .bot(bot), 
        .head(head), .p0m1_l(p0_l[63]), .p1m1_l(p1_l[63]), .p2m1_l(p2_l[63])
         );
  mul_ppgen3 I1_63_ ( .cout(cout[63]), .p0_l(p0_l[63]), .p1_l(p1_l[63]), 
        .p2_l(p2_l[63]), .sum(sum[63]), .am2(a[61]), .am4(a[59]), .a(a[63]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[62]), .p1m1_l(p1_l[62]), 
        .p2m1_l(p2_l[62]) );
  mul_ppgen3 I1_62_ ( .cout(cout[62]), .p0_l(p0_l[62]), .p1_l(p1_l[62]), 
        .p2_l(p2_l[62]), .sum(sum[62]), .am2(a[60]), .am4(a[58]), .a(a[62]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[61]), .p1m1_l(p1_l[61]), 
        .p2m1_l(p2_l[61]) );
  mul_ppgen3 I1_61_ ( .cout(cout[61]), .p0_l(p0_l[61]), .p1_l(p1_l[61]), 
        .p2_l(p2_l[61]), .sum(sum[61]), .am2(a[59]), .am4(a[57]), .a(a[61]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[60]), .p1m1_l(p1_l[60]), 
        .p2m1_l(p2_l[60]) );
  mul_ppgen3 I1_60_ ( .cout(cout[60]), .p0_l(p0_l[60]), .p1_l(p1_l[60]), 
        .p2_l(p2_l[60]), .sum(sum[60]), .am2(a[58]), .am4(a[56]), .a(a[60]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[59]), .p1m1_l(p1_l[59]), 
        .p2m1_l(p2_l[59]) );
  mul_ppgen3 I1_59_ ( .cout(cout[59]), .p0_l(p0_l[59]), .p1_l(p1_l[59]), 
        .p2_l(p2_l[59]), .sum(sum[59]), .am2(a[57]), .am4(a[55]), .a(a[59]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[58]), .p1m1_l(p1_l[58]), 
        .p2m1_l(p2_l[58]) );
  mul_ppgen3 I1_58_ ( .cout(cout[58]), .p0_l(p0_l[58]), .p1_l(p1_l[58]), 
        .p2_l(p2_l[58]), .sum(sum[58]), .am2(a[56]), .am4(a[54]), .a(a[58]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[57]), .p1m1_l(p1_l[57]), 
        .p2m1_l(p2_l[57]) );
  mul_ppgen3 I1_57_ ( .cout(cout[57]), .p0_l(p0_l[57]), .p1_l(p1_l[57]), 
        .p2_l(p2_l[57]), .sum(sum[57]), .am2(a[55]), .am4(a[53]), .a(a[57]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[56]), .p1m1_l(p1_l[56]), 
        .p2m1_l(p2_l[56]) );
  mul_ppgen3 I1_56_ ( .cout(cout[56]), .p0_l(p0_l[56]), .p1_l(p1_l[56]), 
        .p2_l(p2_l[56]), .sum(sum[56]), .am2(a[54]), .am4(a[52]), .a(a[56]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[55]), .p1m1_l(p1_l[55]), 
        .p2m1_l(p2_l[55]) );
  mul_ppgen3 I1_55_ ( .cout(cout[55]), .p0_l(p0_l[55]), .p1_l(p1_l[55]), 
        .p2_l(p2_l[55]), .sum(sum[55]), .am2(a[53]), .am4(a[51]), .a(a[55]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[54]), .p1m1_l(p1_l[54]), 
        .p2m1_l(p2_l[54]) );
  mul_ppgen3 I1_54_ ( .cout(cout[54]), .p0_l(p0_l[54]), .p1_l(p1_l[54]), 
        .p2_l(p2_l[54]), .sum(sum[54]), .am2(a[52]), .am4(a[50]), .a(a[54]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[53]), .p1m1_l(p1_l[53]), 
        .p2m1_l(p2_l[53]) );
  mul_ppgen3 I1_53_ ( .cout(cout[53]), .p0_l(p0_l[53]), .p1_l(p1_l[53]), 
        .p2_l(p2_l[53]), .sum(sum[53]), .am2(a[51]), .am4(a[49]), .a(a[53]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[52]), .p1m1_l(p1_l[52]), 
        .p2m1_l(p2_l[52]) );
  mul_ppgen3 I1_52_ ( .cout(cout[52]), .p0_l(p0_l[52]), .p1_l(p1_l[52]), 
        .p2_l(p2_l[52]), .sum(sum[52]), .am2(a[50]), .am4(a[48]), .a(a[52]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[51]), .p1m1_l(p1_l[51]), 
        .p2m1_l(p2_l[51]) );
  mul_ppgen3 I1_51_ ( .cout(cout[51]), .p0_l(p0_l[51]), .p1_l(p1_l[51]), 
        .p2_l(p2_l[51]), .sum(sum[51]), .am2(a[49]), .am4(a[47]), .a(a[51]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[50]), .p1m1_l(p1_l[50]), 
        .p2m1_l(p2_l[50]) );
  mul_ppgen3 I1_50_ ( .cout(cout[50]), .p0_l(p0_l[50]), .p1_l(p1_l[50]), 
        .p2_l(p2_l[50]), .sum(sum[50]), .am2(a[48]), .am4(a[46]), .a(a[50]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[49]), .p1m1_l(p1_l[49]), 
        .p2m1_l(p2_l[49]) );
  mul_ppgen3 I1_49_ ( .cout(cout[49]), .p0_l(p0_l[49]), .p1_l(p1_l[49]), 
        .p2_l(p2_l[49]), .sum(sum[49]), .am2(a[47]), .am4(a[45]), .a(a[49]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[48]), .p1m1_l(p1_l[48]), 
        .p2m1_l(p2_l[48]) );
  mul_ppgen3 I1_48_ ( .cout(cout[48]), .p0_l(p0_l[48]), .p1_l(p1_l[48]), 
        .p2_l(p2_l[48]), .sum(sum[48]), .am2(a[46]), .am4(a[44]), .a(a[48]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[47]), .p1m1_l(p1_l[47]), 
        .p2m1_l(p2_l[47]) );
  mul_ppgen3 I1_47_ ( .cout(cout[47]), .p0_l(p0_l[47]), .p1_l(p1_l[47]), 
        .p2_l(p2_l[47]), .sum(sum[47]), .am2(a[45]), .am4(a[43]), .a(a[47]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[46]), .p1m1_l(p1_l[46]), 
        .p2m1_l(p2_l[46]) );
  mul_ppgen3 I1_46_ ( .cout(cout[46]), .p0_l(p0_l[46]), .p1_l(p1_l[46]), 
        .p2_l(p2_l[46]), .sum(sum[46]), .am2(a[44]), .am4(a[42]), .a(a[46]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[45]), .p1m1_l(p1_l[45]), 
        .p2m1_l(p2_l[45]) );
  mul_ppgen3 I1_45_ ( .cout(cout[45]), .p0_l(p0_l[45]), .p1_l(p1_l[45]), 
        .p2_l(p2_l[45]), .sum(sum[45]), .am2(a[43]), .am4(a[41]), .a(a[45]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[44]), .p1m1_l(p1_l[44]), 
        .p2m1_l(p2_l[44]) );
  mul_ppgen3 I1_44_ ( .cout(cout[44]), .p0_l(p0_l[44]), .p1_l(p1_l[44]), 
        .p2_l(p2_l[44]), .sum(sum[44]), .am2(a[42]), .am4(a[40]), .a(a[44]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[43]), .p1m1_l(p1_l[43]), 
        .p2m1_l(p2_l[43]) );
  mul_ppgen3 I1_43_ ( .cout(cout[43]), .p0_l(p0_l[43]), .p1_l(p1_l[43]), 
        .p2_l(p2_l[43]), .sum(sum[43]), .am2(a[41]), .am4(a[39]), .a(a[43]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[42]), .p1m1_l(p1_l[42]), 
        .p2m1_l(p2_l[42]) );
  mul_ppgen3 I1_42_ ( .cout(cout[42]), .p0_l(p0_l[42]), .p1_l(p1_l[42]), 
        .p2_l(p2_l[42]), .sum(sum[42]), .am2(a[40]), .am4(a[38]), .a(a[42]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[41]), .p1m1_l(p1_l[41]), 
        .p2m1_l(p2_l[41]) );
  mul_ppgen3 I1_41_ ( .cout(cout[41]), .p0_l(p0_l[41]), .p1_l(p1_l[41]), 
        .p2_l(p2_l[41]), .sum(sum[41]), .am2(a[39]), .am4(a[37]), .a(a[41]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[40]), .p1m1_l(p1_l[40]), 
        .p2m1_l(p2_l[40]) );
  mul_ppgen3 I1_40_ ( .cout(cout[40]), .p0_l(p0_l[40]), .p1_l(p1_l[40]), 
        .p2_l(p2_l[40]), .sum(sum[40]), .am2(a[38]), .am4(a[36]), .a(a[40]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[39]), .p1m1_l(p1_l[39]), 
        .p2m1_l(p2_l[39]) );
  mul_ppgen3 I1_39_ ( .cout(cout[39]), .p0_l(p0_l[39]), .p1_l(p1_l[39]), 
        .p2_l(p2_l[39]), .sum(sum[39]), .am2(a[37]), .am4(a[35]), .a(a[39]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[38]), .p1m1_l(p1_l[38]), 
        .p2m1_l(p2_l[38]) );
  mul_ppgen3 I1_38_ ( .cout(cout[38]), .p0_l(p0_l[38]), .p1_l(p1_l[38]), 
        .p2_l(p2_l[38]), .sum(sum[38]), .am2(a[36]), .am4(a[34]), .a(a[38]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[37]), .p1m1_l(p1_l[37]), 
        .p2m1_l(p2_l[37]) );
  mul_ppgen3 I1_37_ ( .cout(cout[37]), .p0_l(p0_l[37]), .p1_l(p1_l[37]), 
        .p2_l(p2_l[37]), .sum(sum[37]), .am2(a[35]), .am4(a[33]), .a(a[37]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[36]), .p1m1_l(p1_l[36]), 
        .p2m1_l(p2_l[36]) );
  mul_ppgen3 I1_36_ ( .cout(cout[36]), .p0_l(p0_l[36]), .p1_l(p1_l[36]), 
        .p2_l(p2_l[36]), .sum(sum[36]), .am2(a[34]), .am4(a[32]), .a(a[36]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[35]), .p1m1_l(p1_l[35]), 
        .p2m1_l(p2_l[35]) );
  mul_ppgen3 I1_35_ ( .cout(cout[35]), .p0_l(p0_l[35]), .p1_l(p1_l[35]), 
        .p2_l(p2_l[35]), .sum(sum[35]), .am2(a[33]), .am4(a[31]), .a(a[35]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[34]), .p1m1_l(p1_l[34]), 
        .p2m1_l(p2_l[34]) );
  mul_ppgen3 I1_34_ ( .cout(cout[34]), .p0_l(p0_l[34]), .p1_l(p1_l[34]), 
        .p2_l(p2_l[34]), .sum(sum[34]), .am2(a[32]), .am4(a[30]), .a(a[34]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[33]), .p1m1_l(p1_l[33]), 
        .p2m1_l(p2_l[33]) );
  mul_ppgen3 I1_33_ ( .cout(cout[33]), .p0_l(p0_l[33]), .p1_l(p1_l[33]), 
        .p2_l(p2_l[33]), .sum(sum[33]), .am2(a[31]), .am4(a[29]), .a(a[33]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[32]), .p1m1_l(p1_l[32]), 
        .p2m1_l(p2_l[32]) );
  mul_ppgen3 I1_32_ ( .cout(cout[32]), .p0_l(p0_l[32]), .p1_l(p1_l[32]), 
        .p2_l(p2_l[32]), .sum(sum[32]), .am2(a[30]), .am4(a[28]), .a(a[32]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[31]), .p1m1_l(p1_l[31]), 
        .p2m1_l(p2_l[31]) );
  mul_ppgen3 I1_31_ ( .cout(cout[31]), .p0_l(p0_l[31]), .p1_l(p1_l[31]), 
        .p2_l(p2_l[31]), .sum(sum[31]), .am2(a[29]), .am4(a[27]), .a(a[31]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[30]), .p1m1_l(p1_l[30]), 
        .p2m1_l(p2_l[30]) );
  mul_ppgen3 I1_30_ ( .cout(cout[30]), .p0_l(p0_l[30]), .p1_l(p1_l[30]), 
        .p2_l(p2_l[30]), .sum(sum[30]), .am2(a[28]), .am4(a[26]), .a(a[30]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[29]), .p1m1_l(p1_l[29]), 
        .p2m1_l(p2_l[29]) );
  mul_ppgen3 I1_29_ ( .cout(cout[29]), .p0_l(p0_l[29]), .p1_l(p1_l[29]), 
        .p2_l(p2_l[29]), .sum(sum[29]), .am2(a[27]), .am4(a[25]), .a(a[29]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[28]), .p1m1_l(p1_l[28]), 
        .p2m1_l(p2_l[28]) );
  mul_ppgen3 I1_28_ ( .cout(cout[28]), .p0_l(p0_l[28]), .p1_l(p1_l[28]), 
        .p2_l(p2_l[28]), .sum(sum[28]), .am2(a[26]), .am4(a[24]), .a(a[28]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[27]), .p1m1_l(p1_l[27]), 
        .p2m1_l(p2_l[27]) );
  mul_ppgen3 I1_27_ ( .cout(cout[27]), .p0_l(p0_l[27]), .p1_l(p1_l[27]), 
        .p2_l(p2_l[27]), .sum(sum[27]), .am2(a[25]), .am4(a[23]), .a(a[27]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[26]), .p1m1_l(p1_l[26]), 
        .p2m1_l(p2_l[26]) );
  mul_ppgen3 I1_26_ ( .cout(cout[26]), .p0_l(p0_l[26]), .p1_l(p1_l[26]), 
        .p2_l(p2_l[26]), .sum(sum[26]), .am2(a[24]), .am4(a[22]), .a(a[26]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[25]), .p1m1_l(p1_l[25]), 
        .p2m1_l(p2_l[25]) );
  mul_ppgen3 I1_25_ ( .cout(cout[25]), .p0_l(p0_l[25]), .p1_l(p1_l[25]), 
        .p2_l(p2_l[25]), .sum(sum[25]), .am2(a[23]), .am4(a[21]), .a(a[25]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[24]), .p1m1_l(p1_l[24]), 
        .p2m1_l(p2_l[24]) );
  mul_ppgen3 I1_24_ ( .cout(cout[24]), .p0_l(p0_l[24]), .p1_l(p1_l[24]), 
        .p2_l(p2_l[24]), .sum(sum[24]), .am2(a[22]), .am4(a[20]), .a(a[24]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[23]), .p1m1_l(p1_l[23]), 
        .p2m1_l(p2_l[23]) );
  mul_ppgen3 I1_23_ ( .cout(cout[23]), .p0_l(p0_l[23]), .p1_l(p1_l[23]), 
        .p2_l(p2_l[23]), .sum(sum[23]), .am2(a[21]), .am4(a[19]), .a(a[23]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[22]), .p1m1_l(p1_l[22]), 
        .p2m1_l(p2_l[22]) );
  mul_ppgen3 I1_22_ ( .cout(cout[22]), .p0_l(p0_l[22]), .p1_l(p1_l[22]), 
        .p2_l(p2_l[22]), .sum(sum[22]), .am2(a[20]), .am4(a[18]), .a(a[22]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[21]), .p1m1_l(p1_l[21]), 
        .p2m1_l(p2_l[21]) );
  mul_ppgen3 I1_21_ ( .cout(cout[21]), .p0_l(p0_l[21]), .p1_l(p1_l[21]), 
        .p2_l(p2_l[21]), .sum(sum[21]), .am2(a[19]), .am4(a[17]), .a(a[21]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[20]), .p1m1_l(p1_l[20]), 
        .p2m1_l(p2_l[20]) );
  mul_ppgen3 I1_20_ ( .cout(cout[20]), .p0_l(p0_l[20]), .p1_l(p1_l[20]), 
        .p2_l(p2_l[20]), .sum(sum[20]), .am2(a[18]), .am4(a[16]), .a(a[20]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[19]), .p1m1_l(p1_l[19]), 
        .p2m1_l(p2_l[19]) );
  mul_ppgen3 I1_19_ ( .cout(cout[19]), .p0_l(p0_l[19]), .p1_l(p1_l[19]), 
        .p2_l(p2_l[19]), .sum(sum[19]), .am2(a[17]), .am4(a[15]), .a(a[19]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[18]), .p1m1_l(p1_l[18]), 
        .p2m1_l(p2_l[18]) );
  mul_ppgen3 I1_18_ ( .cout(cout[18]), .p0_l(p0_l[18]), .p1_l(p1_l[18]), 
        .p2_l(p2_l[18]), .sum(sum[18]), .am2(a[16]), .am4(a[14]), .a(a[18]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[17]), .p1m1_l(p1_l[17]), 
        .p2m1_l(p2_l[17]) );
  mul_ppgen3 I1_17_ ( .cout(cout[17]), .p0_l(p0_l[17]), .p1_l(p1_l[17]), 
        .p2_l(p2_l[17]), .sum(sum[17]), .am2(a[15]), .am4(a[13]), .a(a[17]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[16]), .p1m1_l(p1_l[16]), 
        .p2m1_l(p2_l[16]) );
  mul_ppgen3 I1_16_ ( .cout(cout[16]), .p0_l(p0_l[16]), .p1_l(p1_l[16]), 
        .p2_l(p2_l[16]), .sum(sum[16]), .am2(a[14]), .am4(a[12]), .a(a[16]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[15]), .p1m1_l(p1_l[15]), 
        .p2m1_l(p2_l[15]) );
  mul_ppgen3 I1_15_ ( .cout(cout[15]), .p0_l(p0_l[15]), .p1_l(p1_l[15]), 
        .p2_l(p2_l[15]), .sum(sum[15]), .am2(a[13]), .am4(a[11]), .a(a[15]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[14]), .p1m1_l(p1_l[14]), 
        .p2m1_l(p2_l[14]) );
  mul_ppgen3 I1_14_ ( .cout(cout[14]), .p0_l(p0_l[14]), .p1_l(p1_l[14]), 
        .p2_l(p2_l[14]), .sum(sum[14]), .am2(a[12]), .am4(a[10]), .a(a[14]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[13]), .p1m1_l(p1_l[13]), 
        .p2m1_l(p2_l[13]) );
  mul_ppgen3 I1_13_ ( .cout(cout[13]), .p0_l(p0_l[13]), .p1_l(p1_l[13]), 
        .p2_l(p2_l[13]), .sum(sum[13]), .am2(a[11]), .am4(a[9]), .a(a[13]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[12]), .p1m1_l(p1_l[12]), 
        .p2m1_l(p2_l[12]) );
  mul_ppgen3 I1_12_ ( .cout(cout[12]), .p0_l(p0_l[12]), .p1_l(p1_l[12]), 
        .p2_l(p2_l[12]), .sum(sum[12]), .am2(a[10]), .am4(a[8]), .a(a[12]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[11]), .p1m1_l(p1_l[11]), 
        .p2m1_l(p2_l[11]) );
  mul_ppgen3 I1_11_ ( .cout(cout[11]), .p0_l(p0_l[11]), .p1_l(p1_l[11]), 
        .p2_l(p2_l[11]), .sum(sum[11]), .am2(a[9]), .am4(a[7]), .a(a[11]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[10]), .p1m1_l(p1_l[10]), 
        .p2m1_l(p2_l[10]) );
  mul_ppgen3 I1_10_ ( .cout(cout[10]), .p0_l(p0_l[10]), .p1_l(p1_l[10]), 
        .p2_l(p2_l[10]), .sum(sum[10]), .am2(a[8]), .am4(a[6]), .a(a[10]), 
        .b0(b0), .b1(b1), .b2(b2), .p0m1_l(p0_l[9]), .p1m1_l(p1_l[9]), 
        .p2m1_l(p2_l[9]) );
  mul_ppgen3 I1_9_ ( .cout(cout[9]), .p0_l(p0_l[9]), .p1_l(p1_l[9]), .p2_l(
        p2_l[9]), .sum(sum[9]), .am2(a[7]), .am4(a[5]), .a(a[9]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[8]), .p1m1_l(p1_l[8]), .p2m1_l(p2_l[8])
         );
  mul_ppgen3 I1_8_ ( .cout(cout[8]), .p0_l(p0_l[8]), .p1_l(p1_l[8]), .p2_l(
        p2_l[8]), .sum(sum[8]), .am2(a[6]), .am4(a[4]), .a(a[8]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[7]), .p1m1_l(p1_l[7]), .p2m1_l(p2_l[7])
         );
  mul_ppgen3 I1_7_ ( .cout(cout[7]), .p0_l(p0_l[7]), .p1_l(p1_l[7]), .p2_l(
        p2_l[7]), .sum(sum[7]), .am2(a[5]), .am4(a[3]), .a(a[7]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[6]), .p1m1_l(p1_l[6]), .p2m1_l(p2_l[6])
         );
  mul_ppgen3 I1_6_ ( .cout(cout[6]), .p0_l(p0_l[6]), .p1_l(p1_l[6]), .p2_l(
        p2_l[6]), .sum(sum[6]), .am2(a[4]), .am4(a[2]), .a(a[6]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[5]), .p1m1_l(p1_l[5]), .p2m1_l(p2_l[5])
         );
  mul_ppgen3 I1_5_ ( .cout(cout[5]), .p0_l(p0_l[5]), .p1_l(p1_l[5]), .p2_l(
        p2_l[5]), .sum(sum[5]), .am2(a[3]), .am4(a[1]), .a(a[5]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[4]), .p1m1_l(p1_l[4]), .p2m1_l(p2_l[4])
         );
  mul_ppgen3 I1_4_ ( .cout(cout[4]), .p0_l(p0_l[4]), .p1_l(p1_l[4]), .p2_l(
        p2_l[4]), .sum(sum[4]), .am2(a[2]), .am4(a[0]), .a(a[4]), .b0(b0), 
        .b1(b1), .b2(b2), .p0m1_l(p0_l[3]), .p1m1_l(p1_l[3]), .p2m1_l(1'b1) );
  mul_ppgen3lsb4 I0 ( .cout(cout[3:1]), .p0_l(p0_l[3]), .p1_l(p1_l[3]), .sum(
        sum[3:0]), .a(a[3:0]), .b0(b0), .b1(b1) );
endmodule


module mul_array1 ( cout, sum, a, b0, b1, b2, b3, b4, b5, b6, b7, b8, bot, 
        head );
  output [81:4] cout;
  output [81:0] sum;
  input [63:0] a;
  input [2:0] b0;
  input [2:0] b1;
  input [2:0] b2;
  input [2:0] b3;
  input [2:0] b4;
  input [2:0] b5;
  input [2:0] b6;
  input [2:0] b7;
  input [2:0] b8;
  input bot, head;

  wire   [1:0] b5n;
  wire   [1:0] b2n;
  wire   [76:10] s_2;
  wire   [75:11] co;
  wire   [70:2] c_1;
  wire   [76:10] c_2;
  wire   [69:0] s1;
  wire   [70:4] s_1;
  wire   [68:1] c1;
  wire   [68:1] c2;
  wire   [69:0] s2;
  wire   [68:1] c0;
  wire   [69:2] s0;

  mul_negen p1n ( .n0(b5n[0]), .n1(b5n[1]), .b(b5) );
  mul_negen p0n ( .n0(b2n[0]), .n1(b2n[1]), .b(b2) );
  mul_csa42 sc3_71_ ( .sum(sum[71]), .carry(cout[71]), .cout(co[71]), .a(
        c_1[70]), .b(c_2[70]), .c(s_2[71]), .d(s1[65]), .cin(co[70]) );
  mul_csa42 sc3_75_ ( .sum(sum[75]), .carry(cout[75]), .cout(co[75]), .a(1'b0), 
        .b(c_2[74]), .c(s_2[75]), .d(s1[69]), .cin(co[74]) );
  mul_csa42 sc3_74_ ( .sum(sum[74]), .carry(cout[74]), .cout(co[74]), .a(1'b0), 
        .b(c_2[73]), .c(s_2[74]), .d(s1[68]), .cin(co[73]) );
  mul_csa42 sc3_73_ ( .sum(sum[73]), .carry(cout[73]), .cout(co[73]), .a(1'b0), 
        .b(c_2[72]), .c(s_2[73]), .d(s1[67]), .cin(co[72]) );
  mul_csa42 sc3_72_ ( .sum(sum[72]), .carry(cout[72]), .cout(co[72]), .a(1'b0), 
        .b(c_2[71]), .c(s_2[72]), .d(s1[66]), .cin(co[71]) );
  mul_csa42 sc3_76_ ( .sum(sum[76]), .carry(cout[76]), .a(1'b0), .b(c_2[75]), 
        .c(s_2[76]), .d(1'b0), .cin(co[75]) );
  mul_csa42 sc3_70_ ( .sum(sum[70]), .carry(cout[70]), .cout(co[70]), .a(
        c_1[69]), .b(c_2[69]), .c(s_2[70]), .d(s_1[70]), .cin(co[69]) );
  mul_csa42 sc3_69_ ( .sum(sum[69]), .carry(cout[69]), .cout(co[69]), .a(
        c_1[68]), .b(c_2[68]), .c(s_2[69]), .d(s_1[69]), .cin(co[68]) );
  mul_csa42 sc3_68_ ( .sum(sum[68]), .carry(cout[68]), .cout(co[68]), .a(
        c_1[67]), .b(c_2[67]), .c(s_2[68]), .d(s_1[68]), .cin(co[67]) );
  mul_csa42 sc3_67_ ( .sum(sum[67]), .carry(cout[67]), .cout(co[67]), .a(
        c_1[66]), .b(c_2[66]), .c(s_2[67]), .d(s_1[67]), .cin(co[66]) );
  mul_csa42 sc3_66_ ( .sum(sum[66]), .carry(cout[66]), .cout(co[66]), .a(
        c_1[65]), .b(c_2[65]), .c(s_2[66]), .d(s_1[66]), .cin(co[65]) );
  mul_csa42 sc3_65_ ( .sum(sum[65]), .carry(cout[65]), .cout(co[65]), .a(
        c_1[64]), .b(c_2[64]), .c(s_2[65]), .d(s_1[65]), .cin(co[64]) );
  mul_csa42 sc3_64_ ( .sum(sum[64]), .carry(cout[64]), .cout(co[64]), .a(
        c_1[63]), .b(c_2[63]), .c(s_2[64]), .d(s_1[64]), .cin(co[63]) );
  mul_csa42 sc3_63_ ( .sum(sum[63]), .carry(cout[63]), .cout(co[63]), .a(
        c_1[62]), .b(c_2[62]), .c(s_2[63]), .d(s_1[63]), .cin(co[62]) );
  mul_csa42 sc3_62_ ( .sum(sum[62]), .carry(cout[62]), .cout(co[62]), .a(
        c_1[61]), .b(c_2[61]), .c(s_2[62]), .d(s_1[62]), .cin(co[61]) );
  mul_csa42 sc3_61_ ( .sum(sum[61]), .carry(cout[61]), .cout(co[61]), .a(
        c_1[60]), .b(c_2[60]), .c(s_2[61]), .d(s_1[61]), .cin(co[60]) );
  mul_csa42 sc3_60_ ( .sum(sum[60]), .carry(cout[60]), .cout(co[60]), .a(
        c_1[59]), .b(c_2[59]), .c(s_2[60]), .d(s_1[60]), .cin(co[59]) );
  mul_csa42 sc3_59_ ( .sum(sum[59]), .carry(cout[59]), .cout(co[59]), .a(
        c_1[58]), .b(c_2[58]), .c(s_2[59]), .d(s_1[59]), .cin(co[58]) );
  mul_csa42 sc3_58_ ( .sum(sum[58]), .carry(cout[58]), .cout(co[58]), .a(
        c_1[57]), .b(c_2[57]), .c(s_2[58]), .d(s_1[58]), .cin(co[57]) );
  mul_csa42 sc3_57_ ( .sum(sum[57]), .carry(cout[57]), .cout(co[57]), .a(
        c_1[56]), .b(c_2[56]), .c(s_2[57]), .d(s_1[57]), .cin(co[56]) );
  mul_csa42 sc3_56_ ( .sum(sum[56]), .carry(cout[56]), .cout(co[56]), .a(
        c_1[55]), .b(c_2[55]), .c(s_2[56]), .d(s_1[56]), .cin(co[55]) );
  mul_csa42 sc3_55_ ( .sum(sum[55]), .carry(cout[55]), .cout(co[55]), .a(
        c_1[54]), .b(c_2[54]), .c(s_2[55]), .d(s_1[55]), .cin(co[54]) );
  mul_csa42 sc3_54_ ( .sum(sum[54]), .carry(cout[54]), .cout(co[54]), .a(
        c_1[53]), .b(c_2[53]), .c(s_2[54]), .d(s_1[54]), .cin(co[53]) );
  mul_csa42 sc3_53_ ( .sum(sum[53]), .carry(cout[53]), .cout(co[53]), .a(
        c_1[52]), .b(c_2[52]), .c(s_2[53]), .d(s_1[53]), .cin(co[52]) );
  mul_csa42 sc3_52_ ( .sum(sum[52]), .carry(cout[52]), .cout(co[52]), .a(
        c_1[51]), .b(c_2[51]), .c(s_2[52]), .d(s_1[52]), .cin(co[51]) );
  mul_csa42 sc3_51_ ( .sum(sum[51]), .carry(cout[51]), .cout(co[51]), .a(
        c_1[50]), .b(c_2[50]), .c(s_2[51]), .d(s_1[51]), .cin(co[50]) );
  mul_csa42 sc3_50_ ( .sum(sum[50]), .carry(cout[50]), .cout(co[50]), .a(
        c_1[49]), .b(c_2[49]), .c(s_2[50]), .d(s_1[50]), .cin(co[49]) );
  mul_csa42 sc3_49_ ( .sum(sum[49]), .carry(cout[49]), .cout(co[49]), .a(
        c_1[48]), .b(c_2[48]), .c(s_2[49]), .d(s_1[49]), .cin(co[48]) );
  mul_csa42 sc3_48_ ( .sum(sum[48]), .carry(cout[48]), .cout(co[48]), .a(
        c_1[47]), .b(c_2[47]), .c(s_2[48]), .d(s_1[48]), .cin(co[47]) );
  mul_csa42 sc3_47_ ( .sum(sum[47]), .carry(cout[47]), .cout(co[47]), .a(
        c_1[46]), .b(c_2[46]), .c(s_2[47]), .d(s_1[47]), .cin(co[46]) );
  mul_csa42 sc3_46_ ( .sum(sum[46]), .carry(cout[46]), .cout(co[46]), .a(
        c_1[45]), .b(c_2[45]), .c(s_2[46]), .d(s_1[46]), .cin(co[45]) );
  mul_csa42 sc3_45_ ( .sum(sum[45]), .carry(cout[45]), .cout(co[45]), .a(
        c_1[44]), .b(c_2[44]), .c(s_2[45]), .d(s_1[45]), .cin(co[44]) );
  mul_csa42 sc3_44_ ( .sum(sum[44]), .carry(cout[44]), .cout(co[44]), .a(
        c_1[43]), .b(c_2[43]), .c(s_2[44]), .d(s_1[44]), .cin(co[43]) );
  mul_csa42 sc3_43_ ( .sum(sum[43]), .carry(cout[43]), .cout(co[43]), .a(
        c_1[42]), .b(c_2[42]), .c(s_2[43]), .d(s_1[43]), .cin(co[42]) );
  mul_csa42 sc3_42_ ( .sum(sum[42]), .carry(cout[42]), .cout(co[42]), .a(
        c_1[41]), .b(c_2[41]), .c(s_2[42]), .d(s_1[42]), .cin(co[41]) );
  mul_csa42 sc3_41_ ( .sum(sum[41]), .carry(cout[41]), .cout(co[41]), .a(
        c_1[40]), .b(c_2[40]), .c(s_2[41]), .d(s_1[41]), .cin(co[40]) );
  mul_csa42 sc3_40_ ( .sum(sum[40]), .carry(cout[40]), .cout(co[40]), .a(
        c_1[39]), .b(c_2[39]), .c(s_2[40]), .d(s_1[40]), .cin(co[39]) );
  mul_csa42 sc3_39_ ( .sum(sum[39]), .carry(cout[39]), .cout(co[39]), .a(
        c_1[38]), .b(c_2[38]), .c(s_2[39]), .d(s_1[39]), .cin(co[38]) );
  mul_csa42 sc3_38_ ( .sum(sum[38]), .carry(cout[38]), .cout(co[38]), .a(
        c_1[37]), .b(c_2[37]), .c(s_2[38]), .d(s_1[38]), .cin(co[37]) );
  mul_csa42 sc3_37_ ( .sum(sum[37]), .carry(cout[37]), .cout(co[37]), .a(
        c_1[36]), .b(c_2[36]), .c(s_2[37]), .d(s_1[37]), .cin(co[36]) );
  mul_csa42 sc3_36_ ( .sum(sum[36]), .carry(cout[36]), .cout(co[36]), .a(
        c_1[35]), .b(c_2[35]), .c(s_2[36]), .d(s_1[36]), .cin(co[35]) );
  mul_csa42 sc3_35_ ( .sum(sum[35]), .carry(cout[35]), .cout(co[35]), .a(
        c_1[34]), .b(c_2[34]), .c(s_2[35]), .d(s_1[35]), .cin(co[34]) );
  mul_csa42 sc3_34_ ( .sum(sum[34]), .carry(cout[34]), .cout(co[34]), .a(
        c_1[33]), .b(c_2[33]), .c(s_2[34]), .d(s_1[34]), .cin(co[33]) );
  mul_csa42 sc3_33_ ( .sum(sum[33]), .carry(cout[33]), .cout(co[33]), .a(
        c_1[32]), .b(c_2[32]), .c(s_2[33]), .d(s_1[33]), .cin(co[32]) );
  mul_csa42 sc3_32_ ( .sum(sum[32]), .carry(cout[32]), .cout(co[32]), .a(
        c_1[31]), .b(c_2[31]), .c(s_2[32]), .d(s_1[32]), .cin(co[31]) );
  mul_csa42 sc3_31_ ( .sum(sum[31]), .carry(cout[31]), .cout(co[31]), .a(
        c_1[30]), .b(c_2[30]), .c(s_2[31]), .d(s_1[31]), .cin(co[30]) );
  mul_csa42 sc3_30_ ( .sum(sum[30]), .carry(cout[30]), .cout(co[30]), .a(
        c_1[29]), .b(c_2[29]), .c(s_2[30]), .d(s_1[30]), .cin(co[29]) );
  mul_csa42 sc3_29_ ( .sum(sum[29]), .carry(cout[29]), .cout(co[29]), .a(
        c_1[28]), .b(c_2[28]), .c(s_2[29]), .d(s_1[29]), .cin(co[28]) );
  mul_csa42 sc3_28_ ( .sum(sum[28]), .carry(cout[28]), .cout(co[28]), .a(
        c_1[27]), .b(c_2[27]), .c(s_2[28]), .d(s_1[28]), .cin(co[27]) );
  mul_csa42 sc3_27_ ( .sum(sum[27]), .carry(cout[27]), .cout(co[27]), .a(
        c_1[26]), .b(c_2[26]), .c(s_2[27]), .d(s_1[27]), .cin(co[26]) );
  mul_csa42 sc3_26_ ( .sum(sum[26]), .carry(cout[26]), .cout(co[26]), .a(
        c_1[25]), .b(c_2[25]), .c(s_2[26]), .d(s_1[26]), .cin(co[25]) );
  mul_csa42 sc3_25_ ( .sum(sum[25]), .carry(cout[25]), .cout(co[25]), .a(
        c_1[24]), .b(c_2[24]), .c(s_2[25]), .d(s_1[25]), .cin(co[24]) );
  mul_csa42 sc3_24_ ( .sum(sum[24]), .carry(cout[24]), .cout(co[24]), .a(
        c_1[23]), .b(c_2[23]), .c(s_2[24]), .d(s_1[24]), .cin(co[23]) );
  mul_csa42 sc3_23_ ( .sum(sum[23]), .carry(cout[23]), .cout(co[23]), .a(
        c_1[22]), .b(c_2[22]), .c(s_2[23]), .d(s_1[23]), .cin(co[22]) );
  mul_csa42 sc3_22_ ( .sum(sum[22]), .carry(cout[22]), .cout(co[22]), .a(
        c_1[21]), .b(c_2[21]), .c(s_2[22]), .d(s_1[22]), .cin(co[21]) );
  mul_csa42 sc3_21_ ( .sum(sum[21]), .carry(cout[21]), .cout(co[21]), .a(
        c_1[20]), .b(c_2[20]), .c(s_2[21]), .d(s_1[21]), .cin(co[20]) );
  mul_csa42 sc3_20_ ( .sum(sum[20]), .carry(cout[20]), .cout(co[20]), .a(
        c_1[19]), .b(c_2[19]), .c(s_2[20]), .d(s_1[20]), .cin(co[19]) );
  mul_csa42 sc3_19_ ( .sum(sum[19]), .carry(cout[19]), .cout(co[19]), .a(
        c_1[18]), .b(c_2[18]), .c(s_2[19]), .d(s_1[19]), .cin(co[18]) );
  mul_csa42 sc3_18_ ( .sum(sum[18]), .carry(cout[18]), .cout(co[18]), .a(
        c_1[17]), .b(c_2[17]), .c(s_2[18]), .d(s_1[18]), .cin(co[17]) );
  mul_csa42 sc3_17_ ( .sum(sum[17]), .carry(cout[17]), .cout(co[17]), .a(
        c_1[16]), .b(c_2[16]), .c(s_2[17]), .d(s_1[17]), .cin(co[16]) );
  mul_csa42 sc3_16_ ( .sum(sum[16]), .carry(cout[16]), .cout(co[16]), .a(
        c_1[15]), .b(c_2[15]), .c(s_2[16]), .d(s_1[16]), .cin(co[15]) );
  mul_csa42 sc3_15_ ( .sum(sum[15]), .carry(cout[15]), .cout(co[15]), .a(
        c_1[14]), .b(c_2[14]), .c(s_2[15]), .d(s_1[15]), .cin(co[14]) );
  mul_csa42 sc3_14_ ( .sum(sum[14]), .carry(cout[14]), .cout(co[14]), .a(
        c_1[13]), .b(c_2[13]), .c(s_2[14]), .d(s_1[14]), .cin(co[13]) );
  mul_csa42 sc3_13_ ( .sum(sum[13]), .carry(cout[13]), .cout(co[13]), .a(
        c_1[12]), .b(c_2[12]), .c(s_2[13]), .d(s_1[13]), .cin(co[12]) );
  mul_csa42 sc3_12_ ( .sum(sum[12]), .carry(cout[12]), .cout(co[12]), .a(
        c_1[11]), .b(c_2[11]), .c(s_2[12]), .d(s_1[12]), .cin(co[11]) );
  mul_csa42 sc3_11_ ( .sum(sum[11]), .carry(cout[11]), .cout(co[11]), .a(
        c_1[10]), .b(c_2[10]), .c(s_2[11]), .d(s_1[11]), .cin(1'b0) );
  mul_csa32 sc2_2_70_ ( .sum(s_2[70]), .cout(c_2[70]), .a(s2[58]), .b(c2[57]), 
        .c(c1[63]) );
  mul_csa32 sc2_2_69_ ( .sum(s_2[69]), .cout(c_2[69]), .a(s2[57]), .b(c2[56]), 
        .c(c1[62]) );
  mul_csa32 sc2_2_68_ ( .sum(s_2[68]), .cout(c_2[68]), .a(s2[56]), .b(c2[55]), 
        .c(c1[61]) );
  mul_csa32 sc2_2_67_ ( .sum(s_2[67]), .cout(c_2[67]), .a(s2[55]), .b(c2[54]), 
        .c(c1[60]) );
  mul_csa32 sc2_2_66_ ( .sum(s_2[66]), .cout(c_2[66]), .a(s2[54]), .b(c2[53]), 
        .c(c1[59]) );
  mul_csa32 sc2_2_65_ ( .sum(s_2[65]), .cout(c_2[65]), .a(s2[53]), .b(c2[52]), 
        .c(c1[58]) );
  mul_csa32 sc2_2_64_ ( .sum(s_2[64]), .cout(c_2[64]), .a(s2[52]), .b(c2[51]), 
        .c(c1[57]) );
  mul_csa32 sc2_2_63_ ( .sum(s_2[63]), .cout(c_2[63]), .a(s2[51]), .b(c2[50]), 
        .c(c1[56]) );
  mul_csa32 sc2_2_62_ ( .sum(s_2[62]), .cout(c_2[62]), .a(s2[50]), .b(c2[49]), 
        .c(c1[55]) );
  mul_csa32 sc2_2_61_ ( .sum(s_2[61]), .cout(c_2[61]), .a(s2[49]), .b(c2[48]), 
        .c(c1[54]) );
  mul_csa32 sc2_2_60_ ( .sum(s_2[60]), .cout(c_2[60]), .a(s2[48]), .b(c2[47]), 
        .c(c1[53]) );
  mul_csa32 sc2_2_59_ ( .sum(s_2[59]), .cout(c_2[59]), .a(s2[47]), .b(c2[46]), 
        .c(c1[52]) );
  mul_csa32 sc2_2_58_ ( .sum(s_2[58]), .cout(c_2[58]), .a(s2[46]), .b(c2[45]), 
        .c(c1[51]) );
  mul_csa32 sc2_2_57_ ( .sum(s_2[57]), .cout(c_2[57]), .a(s2[45]), .b(c2[44]), 
        .c(c1[50]) );
  mul_csa32 sc2_2_56_ ( .sum(s_2[56]), .cout(c_2[56]), .a(s2[44]), .b(c2[43]), 
        .c(c1[49]) );
  mul_csa32 sc2_2_55_ ( .sum(s_2[55]), .cout(c_2[55]), .a(s2[43]), .b(c2[42]), 
        .c(c1[48]) );
  mul_csa32 sc2_2_54_ ( .sum(s_2[54]), .cout(c_2[54]), .a(s2[42]), .b(c2[41]), 
        .c(c1[47]) );
  mul_csa32 sc2_2_53_ ( .sum(s_2[53]), .cout(c_2[53]), .a(s2[41]), .b(c2[40]), 
        .c(c1[46]) );
  mul_csa32 sc2_2_52_ ( .sum(s_2[52]), .cout(c_2[52]), .a(s2[40]), .b(c2[39]), 
        .c(c1[45]) );
  mul_csa32 sc2_2_51_ ( .sum(s_2[51]), .cout(c_2[51]), .a(s2[39]), .b(c2[38]), 
        .c(c1[44]) );
  mul_csa32 sc2_2_50_ ( .sum(s_2[50]), .cout(c_2[50]), .a(s2[38]), .b(c2[37]), 
        .c(c1[43]) );
  mul_csa32 sc2_2_49_ ( .sum(s_2[49]), .cout(c_2[49]), .a(s2[37]), .b(c2[36]), 
        .c(c1[42]) );
  mul_csa32 sc2_2_48_ ( .sum(s_2[48]), .cout(c_2[48]), .a(s2[36]), .b(c2[35]), 
        .c(c1[41]) );
  mul_csa32 sc2_2_47_ ( .sum(s_2[47]), .cout(c_2[47]), .a(s2[35]), .b(c2[34]), 
        .c(c1[40]) );
  mul_csa32 sc2_2_46_ ( .sum(s_2[46]), .cout(c_2[46]), .a(s2[34]), .b(c2[33]), 
        .c(c1[39]) );
  mul_csa32 sc2_2_45_ ( .sum(s_2[45]), .cout(c_2[45]), .a(s2[33]), .b(c2[32]), 
        .c(c1[38]) );
  mul_csa32 sc2_2_44_ ( .sum(s_2[44]), .cout(c_2[44]), .a(s2[32]), .b(c2[31]), 
        .c(c1[37]) );
  mul_csa32 sc2_2_43_ ( .sum(s_2[43]), .cout(c_2[43]), .a(s2[31]), .b(c2[30]), 
        .c(c1[36]) );
  mul_csa32 sc2_2_42_ ( .sum(s_2[42]), .cout(c_2[42]), .a(s2[30]), .b(c2[29]), 
        .c(c1[35]) );
  mul_csa32 sc2_2_41_ ( .sum(s_2[41]), .cout(c_2[41]), .a(s2[29]), .b(c2[28]), 
        .c(c1[34]) );
  mul_csa32 sc2_2_40_ ( .sum(s_2[40]), .cout(c_2[40]), .a(s2[28]), .b(c2[27]), 
        .c(c1[33]) );
  mul_csa32 sc2_2_39_ ( .sum(s_2[39]), .cout(c_2[39]), .a(s2[27]), .b(c2[26]), 
        .c(c1[32]) );
  mul_csa32 sc2_2_38_ ( .sum(s_2[38]), .cout(c_2[38]), .a(s2[26]), .b(c2[25]), 
        .c(c1[31]) );
  mul_csa32 sc2_2_37_ ( .sum(s_2[37]), .cout(c_2[37]), .a(s2[25]), .b(c2[24]), 
        .c(c1[30]) );
  mul_csa32 sc2_2_36_ ( .sum(s_2[36]), .cout(c_2[36]), .a(s2[24]), .b(c2[23]), 
        .c(c1[29]) );
  mul_csa32 sc2_2_35_ ( .sum(s_2[35]), .cout(c_2[35]), .a(s2[23]), .b(c2[22]), 
        .c(c1[28]) );
  mul_csa32 sc2_2_34_ ( .sum(s_2[34]), .cout(c_2[34]), .a(s2[22]), .b(c2[21]), 
        .c(c1[27]) );
  mul_csa32 sc2_2_33_ ( .sum(s_2[33]), .cout(c_2[33]), .a(s2[21]), .b(c2[20]), 
        .c(c1[26]) );
  mul_csa32 sc2_2_32_ ( .sum(s_2[32]), .cout(c_2[32]), .a(s2[20]), .b(c2[19]), 
        .c(c1[25]) );
  mul_csa32 sc2_2_31_ ( .sum(s_2[31]), .cout(c_2[31]), .a(s2[19]), .b(c2[18]), 
        .c(c1[24]) );
  mul_csa32 sc2_2_30_ ( .sum(s_2[30]), .cout(c_2[30]), .a(s2[18]), .b(c2[17]), 
        .c(c1[23]) );
  mul_csa32 sc2_2_29_ ( .sum(s_2[29]), .cout(c_2[29]), .a(s2[17]), .b(c2[16]), 
        .c(c1[22]) );
  mul_csa32 sc2_2_28_ ( .sum(s_2[28]), .cout(c_2[28]), .a(s2[16]), .b(c2[15]), 
        .c(c1[21]) );
  mul_csa32 sc2_2_27_ ( .sum(s_2[27]), .cout(c_2[27]), .a(s2[15]), .b(c2[14]), 
        .c(c1[20]) );
  mul_csa32 sc2_2_26_ ( .sum(s_2[26]), .cout(c_2[26]), .a(s2[14]), .b(c2[13]), 
        .c(c1[19]) );
  mul_csa32 sc2_2_25_ ( .sum(s_2[25]), .cout(c_2[25]), .a(s2[13]), .b(c2[12]), 
        .c(c1[18]) );
  mul_csa32 sc2_2_24_ ( .sum(s_2[24]), .cout(c_2[24]), .a(s2[12]), .b(c2[11]), 
        .c(c1[17]) );
  mul_csa32 sc2_2_23_ ( .sum(s_2[23]), .cout(c_2[23]), .a(s2[11]), .b(c2[10]), 
        .c(c1[16]) );
  mul_csa32 sc2_2_22_ ( .sum(s_2[22]), .cout(c_2[22]), .a(s2[10]), .b(c2[9]), 
        .c(c1[15]) );
  mul_csa32 sc2_2_21_ ( .sum(s_2[21]), .cout(c_2[21]), .a(s2[9]), .b(c2[8]), 
        .c(c1[14]) );
  mul_csa32 sc2_2_20_ ( .sum(s_2[20]), .cout(c_2[20]), .a(s2[8]), .b(c2[7]), 
        .c(c1[13]) );
  mul_csa32 sc2_2_19_ ( .sum(s_2[19]), .cout(c_2[19]), .a(s2[7]), .b(c2[6]), 
        .c(c1[12]) );
  mul_csa32 sc2_2_18_ ( .sum(s_2[18]), .cout(c_2[18]), .a(s2[6]), .b(c2[5]), 
        .c(c1[11]) );
  mul_csa32 sc2_2_17_ ( .sum(s_2[17]), .cout(c_2[17]), .a(s2[5]), .b(c2[4]), 
        .c(c1[10]) );
  mul_csa32 sc2_2_16_ ( .sum(s_2[16]), .cout(c_2[16]), .a(s2[4]), .b(c2[3]), 
        .c(c1[9]) );
  mul_csa32 sc2_2_15_ ( .sum(s_2[15]), .cout(c_2[15]), .a(s2[3]), .b(c2[2]), 
        .c(c1[8]) );
  mul_csa32 sc2_2_14_ ( .sum(s_2[14]), .cout(c_2[14]), .a(s2[2]), .b(c2[1]), 
        .c(c1[7]) );
  mul_csa32 sc2_2_13_ ( .sum(s_2[13]), .cout(c_2[13]), .a(s2[1]), .b(s1[7]), 
        .c(c1[6]) );
  mul_csa32 sc2_2_12_ ( .sum(s_2[12]), .cout(c_2[12]), .a(s2[0]), .b(s1[6]), 
        .c(c1[5]) );
  mul_csa32 sc2_2_11_ ( .sum(s_2[11]), .cout(c_2[11]), .a(b5n[1]), .b(s1[5]), 
        .c(c1[4]) );
  mul_csa32 sc2_2_10_ ( .sum(s_2[10]), .cout(c_2[10]), .a(b5n[0]), .b(s1[4]), 
        .c(c1[3]) );
  mul_csa32 sc2_2_76_ ( .sum(s_2[76]), .cout(c_2[76]), .a(s2[64]), .b(c2[63]), 
        .c(1'b1) );
  mul_csa32 sc2_2_77_ ( .sum(sum[77]), .cout(cout[77]), .a(s2[65]), .b(c2[64]), 
        .c(c_2[76]) );
  mul_csa32 sc2_1_9_ ( .sum(s_1[9]), .cout(c_1[9]), .a(s0[9]), .b(c0[8]), .c(
        s1[3]) );
  mul_csa32 sc2_1_8_ ( .sum(s_1[8]), .cout(c_1[8]), .a(s0[8]), .b(c0[7]), .c(
        s1[2]) );
  mul_csa32 sc2_1_3_ ( .sum(sum[3]), .cout(c_1[3]), .a(s0[3]), .b(c0[2]), .c(
        c_1[2]) );
  mul_csa32 sc3_10_ ( .sum(sum[10]), .cout(cout[10]), .a(c_1[9]), .b(s_1[10]), 
        .c(s_2[10]) );
  mul_csa32 sc3_9_ ( .sum(sum[9]), .cout(cout[9]), .a(c_1[8]), .b(s_1[9]), .c(
        c1[2]) );
  mul_csa32 sc3_8_ ( .sum(sum[8]), .cout(cout[8]), .a(c_1[7]), .b(s_1[8]), .c(
        c1[1]) );
  mul_csa32 sc2_2_71_ ( .sum(s_2[71]), .cout(c_2[71]), .a(s2[59]), .b(c2[58]), 
        .c(c1[64]) );
  mul_csa32 sc2_2_75_ ( .sum(s_2[75]), .cout(c_2[75]), .a(s2[63]), .b(c2[62]), 
        .c(c1[68]) );
  mul_csa32 sc2_2_74_ ( .sum(s_2[74]), .cout(c_2[74]), .a(s2[62]), .b(c2[61]), 
        .c(c1[67]) );
  mul_csa32 sc2_2_73_ ( .sum(s_2[73]), .cout(c_2[73]), .a(s2[61]), .b(c2[60]), 
        .c(c1[66]) );
  mul_csa32 sc2_2_72_ ( .sum(s_2[72]), .cout(c_2[72]), .a(s2[60]), .b(c2[59]), 
        .c(c1[65]) );
  mul_csa32 sc2_1_69_ ( .sum(s_1[69]), .cout(c_1[69]), .a(s0[69]), .b(c0[68]), 
        .c(s1[63]) );
  mul_csa32 sc2_1_68_ ( .sum(s_1[68]), .cout(c_1[68]), .a(s0[68]), .b(c0[67]), 
        .c(s1[62]) );
  mul_csa32 sc2_1_67_ ( .sum(s_1[67]), .cout(c_1[67]), .a(s0[67]), .b(c0[66]), 
        .c(s1[61]) );
  mul_csa32 sc2_1_66_ ( .sum(s_1[66]), .cout(c_1[66]), .a(s0[66]), .b(c0[65]), 
        .c(s1[60]) );
  mul_csa32 sc2_1_65_ ( .sum(s_1[65]), .cout(c_1[65]), .a(s0[65]), .b(c0[64]), 
        .c(s1[59]) );
  mul_csa32 sc2_1_64_ ( .sum(s_1[64]), .cout(c_1[64]), .a(s0[64]), .b(c0[63]), 
        .c(s1[58]) );
  mul_csa32 sc2_1_63_ ( .sum(s_1[63]), .cout(c_1[63]), .a(s0[63]), .b(c0[62]), 
        .c(s1[57]) );
  mul_csa32 sc2_1_62_ ( .sum(s_1[62]), .cout(c_1[62]), .a(s0[62]), .b(c0[61]), 
        .c(s1[56]) );
  mul_csa32 sc2_1_61_ ( .sum(s_1[61]), .cout(c_1[61]), .a(s0[61]), .b(c0[60]), 
        .c(s1[55]) );
  mul_csa32 sc2_1_60_ ( .sum(s_1[60]), .cout(c_1[60]), .a(s0[60]), .b(c0[59]), 
        .c(s1[54]) );
  mul_csa32 sc2_1_59_ ( .sum(s_1[59]), .cout(c_1[59]), .a(s0[59]), .b(c0[58]), 
        .c(s1[53]) );
  mul_csa32 sc2_1_58_ ( .sum(s_1[58]), .cout(c_1[58]), .a(s0[58]), .b(c0[57]), 
        .c(s1[52]) );
  mul_csa32 sc2_1_57_ ( .sum(s_1[57]), .cout(c_1[57]), .a(s0[57]), .b(c0[56]), 
        .c(s1[51]) );
  mul_csa32 sc2_1_56_ ( .sum(s_1[56]), .cout(c_1[56]), .a(s0[56]), .b(c0[55]), 
        .c(s1[50]) );
  mul_csa32 sc2_1_55_ ( .sum(s_1[55]), .cout(c_1[55]), .a(s0[55]), .b(c0[54]), 
        .c(s1[49]) );
  mul_csa32 sc2_1_54_ ( .sum(s_1[54]), .cout(c_1[54]), .a(s0[54]), .b(c0[53]), 
        .c(s1[48]) );
  mul_csa32 sc2_1_53_ ( .sum(s_1[53]), .cout(c_1[53]), .a(s0[53]), .b(c0[52]), 
        .c(s1[47]) );
  mul_csa32 sc2_1_52_ ( .sum(s_1[52]), .cout(c_1[52]), .a(s0[52]), .b(c0[51]), 
        .c(s1[46]) );
  mul_csa32 sc2_1_51_ ( .sum(s_1[51]), .cout(c_1[51]), .a(s0[51]), .b(c0[50]), 
        .c(s1[45]) );
  mul_csa32 sc2_1_50_ ( .sum(s_1[50]), .cout(c_1[50]), .a(s0[50]), .b(c0[49]), 
        .c(s1[44]) );
  mul_csa32 sc2_1_49_ ( .sum(s_1[49]), .cout(c_1[49]), .a(s0[49]), .b(c0[48]), 
        .c(s1[43]) );
  mul_csa32 sc2_1_48_ ( .sum(s_1[48]), .cout(c_1[48]), .a(s0[48]), .b(c0[47]), 
        .c(s1[42]) );
  mul_csa32 sc2_1_47_ ( .sum(s_1[47]), .cout(c_1[47]), .a(s0[47]), .b(c0[46]), 
        .c(s1[41]) );
  mul_csa32 sc2_1_46_ ( .sum(s_1[46]), .cout(c_1[46]), .a(s0[46]), .b(c0[45]), 
        .c(s1[40]) );
  mul_csa32 sc2_1_45_ ( .sum(s_1[45]), .cout(c_1[45]), .a(s0[45]), .b(c0[44]), 
        .c(s1[39]) );
  mul_csa32 sc2_1_44_ ( .sum(s_1[44]), .cout(c_1[44]), .a(s0[44]), .b(c0[43]), 
        .c(s1[38]) );
  mul_csa32 sc2_1_43_ ( .sum(s_1[43]), .cout(c_1[43]), .a(s0[43]), .b(c0[42]), 
        .c(s1[37]) );
  mul_csa32 sc2_1_42_ ( .sum(s_1[42]), .cout(c_1[42]), .a(s0[42]), .b(c0[41]), 
        .c(s1[36]) );
  mul_csa32 sc2_1_41_ ( .sum(s_1[41]), .cout(c_1[41]), .a(s0[41]), .b(c0[40]), 
        .c(s1[35]) );
  mul_csa32 sc2_1_40_ ( .sum(s_1[40]), .cout(c_1[40]), .a(s0[40]), .b(c0[39]), 
        .c(s1[34]) );
  mul_csa32 sc2_1_39_ ( .sum(s_1[39]), .cout(c_1[39]), .a(s0[39]), .b(c0[38]), 
        .c(s1[33]) );
  mul_csa32 sc2_1_38_ ( .sum(s_1[38]), .cout(c_1[38]), .a(s0[38]), .b(c0[37]), 
        .c(s1[32]) );
  mul_csa32 sc2_1_37_ ( .sum(s_1[37]), .cout(c_1[37]), .a(s0[37]), .b(c0[36]), 
        .c(s1[31]) );
  mul_csa32 sc2_1_36_ ( .sum(s_1[36]), .cout(c_1[36]), .a(s0[36]), .b(c0[35]), 
        .c(s1[30]) );
  mul_csa32 sc2_1_35_ ( .sum(s_1[35]), .cout(c_1[35]), .a(s0[35]), .b(c0[34]), 
        .c(s1[29]) );
  mul_csa32 sc2_1_34_ ( .sum(s_1[34]), .cout(c_1[34]), .a(s0[34]), .b(c0[33]), 
        .c(s1[28]) );
  mul_csa32 sc2_1_33_ ( .sum(s_1[33]), .cout(c_1[33]), .a(s0[33]), .b(c0[32]), 
        .c(s1[27]) );
  mul_csa32 sc2_1_32_ ( .sum(s_1[32]), .cout(c_1[32]), .a(s0[32]), .b(c0[31]), 
        .c(s1[26]) );
  mul_csa32 sc2_1_31_ ( .sum(s_1[31]), .cout(c_1[31]), .a(s0[31]), .b(c0[30]), 
        .c(s1[25]) );
  mul_csa32 sc2_1_30_ ( .sum(s_1[30]), .cout(c_1[30]), .a(s0[30]), .b(c0[29]), 
        .c(s1[24]) );
  mul_csa32 sc2_1_29_ ( .sum(s_1[29]), .cout(c_1[29]), .a(s0[29]), .b(c0[28]), 
        .c(s1[23]) );
  mul_csa32 sc2_1_28_ ( .sum(s_1[28]), .cout(c_1[28]), .a(s0[28]), .b(c0[27]), 
        .c(s1[22]) );
  mul_csa32 sc2_1_27_ ( .sum(s_1[27]), .cout(c_1[27]), .a(s0[27]), .b(c0[26]), 
        .c(s1[21]) );
  mul_csa32 sc2_1_26_ ( .sum(s_1[26]), .cout(c_1[26]), .a(s0[26]), .b(c0[25]), 
        .c(s1[20]) );
  mul_csa32 sc2_1_25_ ( .sum(s_1[25]), .cout(c_1[25]), .a(s0[25]), .b(c0[24]), 
        .c(s1[19]) );
  mul_csa32 sc2_1_24_ ( .sum(s_1[24]), .cout(c_1[24]), .a(s0[24]), .b(c0[23]), 
        .c(s1[18]) );
  mul_csa32 sc2_1_23_ ( .sum(s_1[23]), .cout(c_1[23]), .a(s0[23]), .b(c0[22]), 
        .c(s1[17]) );
  mul_csa32 sc2_1_22_ ( .sum(s_1[22]), .cout(c_1[22]), .a(s0[22]), .b(c0[21]), 
        .c(s1[16]) );
  mul_csa32 sc2_1_21_ ( .sum(s_1[21]), .cout(c_1[21]), .a(s0[21]), .b(c0[20]), 
        .c(s1[15]) );
  mul_csa32 sc2_1_20_ ( .sum(s_1[20]), .cout(c_1[20]), .a(s0[20]), .b(c0[19]), 
        .c(s1[14]) );
  mul_csa32 sc2_1_19_ ( .sum(s_1[19]), .cout(c_1[19]), .a(s0[19]), .b(c0[18]), 
        .c(s1[13]) );
  mul_csa32 sc2_1_18_ ( .sum(s_1[18]), .cout(c_1[18]), .a(s0[18]), .b(c0[17]), 
        .c(s1[12]) );
  mul_csa32 sc2_1_17_ ( .sum(s_1[17]), .cout(c_1[17]), .a(s0[17]), .b(c0[16]), 
        .c(s1[11]) );
  mul_csa32 sc2_1_16_ ( .sum(s_1[16]), .cout(c_1[16]), .a(s0[16]), .b(c0[15]), 
        .c(s1[10]) );
  mul_csa32 sc2_1_15_ ( .sum(s_1[15]), .cout(c_1[15]), .a(s0[15]), .b(c0[14]), 
        .c(s1[9]) );
  mul_csa32 sc2_1_14_ ( .sum(s_1[14]), .cout(c_1[14]), .a(s0[14]), .b(c0[13]), 
        .c(s1[8]) );
  mul_csa32 sc2_1_7_ ( .sum(s_1[7]), .cout(c_1[7]), .a(s0[7]), .b(c0[6]), .c(
        s1[1]) );
  mul_csa32 sc2_1_6_ ( .sum(s_1[6]), .cout(c_1[6]), .a(s0[6]), .b(c0[5]), .c(
        s1[0]) );
  mul_csa32 sc2_1_5_ ( .sum(s_1[5]), .cout(c_1[5]), .a(s0[5]), .b(c0[4]), .c(
        b2n[1]) );
  mul_csa32 sc2_1_4_ ( .sum(s_1[4]), .cout(c_1[4]), .a(s0[4]), .b(c0[3]), .c(
        b2n[0]) );
  mul_ha sc2_1_10_ ( .cout(c_1[10]), .sum(s_1[10]), .a(s0[10]), .b(c0[9]) );
  mul_ha sc3_7_ ( .cout(cout[7]), .sum(sum[7]), .a(c_1[6]), .b(s_1[7]) );
  mul_ha sc3_6_ ( .cout(cout[6]), .sum(sum[6]), .a(c_1[5]), .b(s_1[6]) );
  mul_ha sc3_5_ ( .cout(cout[5]), .sum(sum[5]), .a(c_1[4]), .b(s_1[5]) );
  mul_ha sc3_4_ ( .cout(cout[4]), .sum(sum[4]), .a(c_1[3]), .b(s_1[4]) );
  mul_ha sc2_2_81_ ( .cout(cout[81]), .sum(sum[81]), .a(s2[69]), .b(c2[68]) );
  mul_ha sc2_2_80_ ( .cout(cout[80]), .sum(sum[80]), .a(s2[68]), .b(c2[67]) );
  mul_ha sc2_2_79_ ( .cout(cout[79]), .sum(sum[79]), .a(s2[67]), .b(c2[66]) );
  mul_ha sc2_2_78_ ( .cout(cout[78]), .sum(sum[78]), .a(s2[66]), .b(c2[65]) );
  mul_ha sc2_1_70_ ( .cout(c_1[70]), .sum(s_1[70]), .a(1'b1), .b(s1[64]) );
  mul_ha sc2_1_2_ ( .cout(c_1[2]), .sum(sum[2]), .a(s0[2]), .b(c0[1]) );
  mul_ha sc2_1_13_ ( .cout(c_1[13]), .sum(s_1[13]), .a(s0[13]), .b(c0[12]) );
  mul_ha sc2_1_12_ ( .cout(c_1[12]), .sum(s_1[12]), .a(s0[12]), .b(c0[11]) );
  mul_ha sc2_1_11_ ( .cout(c_1[11]), .sum(s_1[11]), .a(s0[11]), .b(c0[10]) );
  mul_ppgenrow3 I2 ( .cout(c2), .sum(s2), .a(a), .b0(b6), .b1(b7), .b2(b8), 
        .bot(bot), .head(1'b0) );
  mul_ppgenrow3 I1 ( .cout(c1), .sum(s1), .a(a), .b0(b3), .b1(b4), .b2(b5), 
        .bot(1'b1), .head(1'b0) );
  mul_ppgenrow3 I0 ( .cout(c0), .sum({s0, sum[1:0]}), .a(a), .b0(b0), .b1(b1), 
        .b2(b2), .bot(1'b1), .head(head) );
endmodule


module dff_SIZE78 ( din, clk, q, se, si, so );
  input [77:0] din;
  output [77:0] q;
  input [77:0] si;
  output [77:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80;
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C88 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE82 ( din, clk, q, se, si, so );
  input [81:0] din;
  output [81:0] q;
  input [81:0] si;
  output [81:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84;
  assign so[81] = q[81];
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C92 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module mul_mux2 ( z, d0, d1, s );
  input d0, d1, s;
  output z;
  wire   N0, N1, N2;

  SELECT_OP C11 ( .DATA1(d1), .DATA2(d0), .CONTROL1(N0), .CONTROL2(N1), .Z(z)
         );
  GTECH_BUF B_0 ( .A(s), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(s), .Z(N2) );
endmodule


module mul_array2 ( pcout, pcoutx2, psum, psumx2, a0c, a0s, a1c, a1s, areg, 
        bot, pc, ps, x2 );
  output [98:0] pcout;
  output [98:0] psum;
  input [81:4] a0c;
  input [81:0] a0s;
  input [81:4] a1c;
  input [81:0] a1s;
  input [96:0] areg;
  input [98:30] pc;
  input [98:31] ps;
  input bot, x2;
  output pcoutx2, psumx2;
  wire   ainx2, s1x2, c1x2;
  wire   [96:0] ain;
  wire   [67:20] co;
  wire   [81:15] c3;
  wire   [96:0] c2;
  wire   [96:0] s2;
  wire   [81:15] s3;
  wire   [82:0] s1;
  wire   [82:0] c1;

  mul_mux2 sh_82_ ( .z(ain[82]), .d0(areg[82]), .d1(areg[83]), .s(x2) );
  mul_mux2 sh_68_ ( .z(ain[68]), .d0(areg[68]), .d1(areg[69]), .s(x2) );
  mul_mux2 sh_67_ ( .z(ain[67]), .d0(areg[67]), .d1(areg[68]), .s(x2) );
  mul_mux2 sh_66_ ( .z(ain[66]), .d0(areg[66]), .d1(areg[67]), .s(x2) );
  mul_mux2 sh_65_ ( .z(ain[65]), .d0(areg[65]), .d1(areg[66]), .s(x2) );
  mul_mux2 sh_64_ ( .z(ain[64]), .d0(areg[64]), .d1(areg[65]), .s(x2) );
  mul_mux2 sh_63_ ( .z(ain[63]), .d0(areg[63]), .d1(areg[64]), .s(x2) );
  mul_mux2 sh_62_ ( .z(ain[62]), .d0(areg[62]), .d1(areg[63]), .s(x2) );
  mul_mux2 sh_61_ ( .z(ain[61]), .d0(areg[61]), .d1(areg[62]), .s(x2) );
  mul_mux2 sh_60_ ( .z(ain[60]), .d0(areg[60]), .d1(areg[61]), .s(x2) );
  mul_mux2 sh_59_ ( .z(ain[59]), .d0(areg[59]), .d1(areg[60]), .s(x2) );
  mul_mux2 sh_58_ ( .z(ain[58]), .d0(areg[58]), .d1(areg[59]), .s(x2) );
  mul_mux2 sh_57_ ( .z(ain[57]), .d0(areg[57]), .d1(areg[58]), .s(x2) );
  mul_mux2 sh_56_ ( .z(ain[56]), .d0(areg[56]), .d1(areg[57]), .s(x2) );
  mul_mux2 sh_55_ ( .z(ain[55]), .d0(areg[55]), .d1(areg[56]), .s(x2) );
  mul_mux2 sh_54_ ( .z(ain[54]), .d0(areg[54]), .d1(areg[55]), .s(x2) );
  mul_mux2 sh_53_ ( .z(ain[53]), .d0(areg[53]), .d1(areg[54]), .s(x2) );
  mul_mux2 sh_52_ ( .z(ain[52]), .d0(areg[52]), .d1(areg[53]), .s(x2) );
  mul_mux2 sh_51_ ( .z(ain[51]), .d0(areg[51]), .d1(areg[52]), .s(x2) );
  mul_mux2 sh_50_ ( .z(ain[50]), .d0(areg[50]), .d1(areg[51]), .s(x2) );
  mul_mux2 sh_49_ ( .z(ain[49]), .d0(areg[49]), .d1(areg[50]), .s(x2) );
  mul_mux2 sh_48_ ( .z(ain[48]), .d0(areg[48]), .d1(areg[49]), .s(x2) );
  mul_mux2 sh_47_ ( .z(ain[47]), .d0(areg[47]), .d1(areg[48]), .s(x2) );
  mul_mux2 sh_46_ ( .z(ain[46]), .d0(areg[46]), .d1(areg[47]), .s(x2) );
  mul_mux2 sh_45_ ( .z(ain[45]), .d0(areg[45]), .d1(areg[46]), .s(x2) );
  mul_mux2 sh_44_ ( .z(ain[44]), .d0(areg[44]), .d1(areg[45]), .s(x2) );
  mul_mux2 sh_43_ ( .z(ain[43]), .d0(areg[43]), .d1(areg[44]), .s(x2) );
  mul_mux2 sh_42_ ( .z(ain[42]), .d0(areg[42]), .d1(areg[43]), .s(x2) );
  mul_mux2 sh_41_ ( .z(ain[41]), .d0(areg[41]), .d1(areg[42]), .s(x2) );
  mul_mux2 sh_40_ ( .z(ain[40]), .d0(areg[40]), .d1(areg[41]), .s(x2) );
  mul_mux2 sh_39_ ( .z(ain[39]), .d0(areg[39]), .d1(areg[40]), .s(x2) );
  mul_mux2 sh_38_ ( .z(ain[38]), .d0(areg[38]), .d1(areg[39]), .s(x2) );
  mul_mux2 sh_37_ ( .z(ain[37]), .d0(areg[37]), .d1(areg[38]), .s(x2) );
  mul_mux2 sh_36_ ( .z(ain[36]), .d0(areg[36]), .d1(areg[37]), .s(x2) );
  mul_mux2 sh_35_ ( .z(ain[35]), .d0(areg[35]), .d1(areg[36]), .s(x2) );
  mul_mux2 sh_34_ ( .z(ain[34]), .d0(areg[34]), .d1(areg[35]), .s(x2) );
  mul_mux2 sh_33_ ( .z(ain[33]), .d0(areg[33]), .d1(areg[34]), .s(x2) );
  mul_mux2 sh_32_ ( .z(ain[32]), .d0(areg[32]), .d1(areg[33]), .s(x2) );
  mul_mux2 sh_31_ ( .z(ain[31]), .d0(areg[31]), .d1(areg[32]), .s(x2) );
  mul_mux2 sh_30_ ( .z(ain[30]), .d0(areg[30]), .d1(areg[31]), .s(x2) );
  mul_mux2 sh_29_ ( .z(ain[29]), .d0(areg[29]), .d1(areg[30]), .s(x2) );
  mul_mux2 sh_28_ ( .z(ain[28]), .d0(areg[28]), .d1(areg[29]), .s(x2) );
  mul_mux2 sh_27_ ( .z(ain[27]), .d0(areg[27]), .d1(areg[28]), .s(x2) );
  mul_mux2 sh_26_ ( .z(ain[26]), .d0(areg[26]), .d1(areg[27]), .s(x2) );
  mul_mux2 sh_25_ ( .z(ain[25]), .d0(areg[25]), .d1(areg[26]), .s(x2) );
  mul_mux2 sh_24_ ( .z(ain[24]), .d0(areg[24]), .d1(areg[25]), .s(x2) );
  mul_mux2 sh_23_ ( .z(ain[23]), .d0(areg[23]), .d1(areg[24]), .s(x2) );
  mul_mux2 sh_22_ ( .z(ain[22]), .d0(areg[22]), .d1(areg[23]), .s(x2) );
  mul_mux2 sh_21_ ( .z(ain[21]), .d0(areg[21]), .d1(areg[22]), .s(x2) );
  mul_mux2 sh_20_ ( .z(ain[20]), .d0(areg[20]), .d1(areg[21]), .s(x2) );
  mul_mux2 sh_96_ ( .z(ain[96]), .d0(areg[96]), .d1(1'b0), .s(x2) );
  mul_mux2 sh_95_ ( .z(ain[95]), .d0(areg[95]), .d1(areg[96]), .s(x2) );
  mul_mux2 sh_94_ ( .z(ain[94]), .d0(areg[94]), .d1(areg[95]), .s(x2) );
  mul_mux2 sh_93_ ( .z(ain[93]), .d0(areg[93]), .d1(areg[94]), .s(x2) );
  mul_mux2 sh_92_ ( .z(ain[92]), .d0(areg[92]), .d1(areg[93]), .s(x2) );
  mul_mux2 sh_91_ ( .z(ain[91]), .d0(areg[91]), .d1(areg[92]), .s(x2) );
  mul_mux2 sh_90_ ( .z(ain[90]), .d0(areg[90]), .d1(areg[91]), .s(x2) );
  mul_mux2 sh_89_ ( .z(ain[89]), .d0(areg[89]), .d1(areg[90]), .s(x2) );
  mul_mux2 sh_88_ ( .z(ain[88]), .d0(areg[88]), .d1(areg[89]), .s(x2) );
  mul_mux2 sh_87_ ( .z(ain[87]), .d0(areg[87]), .d1(areg[88]), .s(x2) );
  mul_mux2 sh_86_ ( .z(ain[86]), .d0(areg[86]), .d1(areg[87]), .s(x2) );
  mul_mux2 sh_85_ ( .z(ain[85]), .d0(areg[85]), .d1(areg[86]), .s(x2) );
  mul_mux2 sh_84_ ( .z(ain[84]), .d0(areg[84]), .d1(areg[85]), .s(x2) );
  mul_mux2 sh_0_ ( .z(ain[0]), .d0(areg[0]), .d1(areg[1]), .s(x2) );
  mul_mux2 sh_81_ ( .z(ain[81]), .d0(areg[81]), .d1(areg[82]), .s(x2) );
  mul_mux2 sh_80_ ( .z(ain[80]), .d0(areg[80]), .d1(areg[81]), .s(x2) );
  mul_mux2 sh_79_ ( .z(ain[79]), .d0(areg[79]), .d1(areg[80]), .s(x2) );
  mul_mux2 sh_78_ ( .z(ain[78]), .d0(areg[78]), .d1(areg[79]), .s(x2) );
  mul_mux2 sh_77_ ( .z(ain[77]), .d0(areg[77]), .d1(areg[78]), .s(x2) );
  mul_mux2 sh_76_ ( .z(ain[76]), .d0(areg[76]), .d1(areg[77]), .s(x2) );
  mul_mux2 sh_75_ ( .z(ain[75]), .d0(areg[75]), .d1(areg[76]), .s(x2) );
  mul_mux2 sh_74_ ( .z(ain[74]), .d0(areg[74]), .d1(areg[75]), .s(x2) );
  mul_mux2 sh_73_ ( .z(ain[73]), .d0(areg[73]), .d1(areg[74]), .s(x2) );
  mul_mux2 sh_72_ ( .z(ain[72]), .d0(areg[72]), .d1(areg[73]), .s(x2) );
  mul_mux2 sh_71_ ( .z(ain[71]), .d0(areg[71]), .d1(areg[72]), .s(x2) );
  mul_mux2 sh_70_ ( .z(ain[70]), .d0(areg[70]), .d1(areg[71]), .s(x2) );
  mul_mux2 sh_69_ ( .z(ain[69]), .d0(areg[69]), .d1(areg[70]), .s(x2) );
  mul_mux2 sh_19_ ( .z(ain[19]), .d0(areg[19]), .d1(areg[20]), .s(x2) );
  mul_mux2 sh_18_ ( .z(ain[18]), .d0(areg[18]), .d1(areg[19]), .s(x2) );
  mul_mux2 sh_17_ ( .z(ain[17]), .d0(areg[17]), .d1(areg[18]), .s(x2) );
  mul_mux2 sh_16_ ( .z(ain[16]), .d0(areg[16]), .d1(areg[17]), .s(x2) );
  mul_mux2 sh_15_ ( .z(ain[15]), .d0(areg[15]), .d1(areg[16]), .s(x2) );
  mul_mux2 sh_4_ ( .z(ain[4]), .d0(areg[4]), .d1(areg[5]), .s(x2) );
  mul_mux2 sh_3_ ( .z(ain[3]), .d0(areg[3]), .d1(areg[4]), .s(x2) );
  mul_mux2 sh_2_ ( .z(ain[2]), .d0(areg[2]), .d1(areg[3]), .s(x2) );
  mul_mux2 sh_1_ ( .z(ain[1]), .d0(areg[1]), .d1(areg[2]), .s(x2) );
  mul_mux2 shx2 ( .z(ainx2), .d0(1'b0), .d1(areg[0]), .s(x2) );
  mul_mux2 sh_83_ ( .z(ain[83]), .d0(areg[83]), .d1(areg[84]), .s(x2) );
  mul_mux2 sh_14_ ( .z(ain[14]), .d0(areg[14]), .d1(areg[15]), .s(x2) );
  mul_mux2 sh_13_ ( .z(ain[13]), .d0(areg[13]), .d1(areg[14]), .s(x2) );
  mul_mux2 sh_12_ ( .z(ain[12]), .d0(areg[12]), .d1(areg[13]), .s(x2) );
  mul_mux2 sh_11_ ( .z(ain[11]), .d0(areg[11]), .d1(areg[12]), .s(x2) );
  mul_mux2 sh_10_ ( .z(ain[10]), .d0(areg[10]), .d1(areg[11]), .s(x2) );
  mul_mux2 sh_9_ ( .z(ain[9]), .d0(areg[9]), .d1(areg[10]), .s(x2) );
  mul_mux2 sh_8_ ( .z(ain[8]), .d0(areg[8]), .d1(areg[9]), .s(x2) );
  mul_mux2 sh_7_ ( .z(ain[7]), .d0(areg[7]), .d1(areg[8]), .s(x2) );
  mul_mux2 sh_6_ ( .z(ain[6]), .d0(areg[6]), .d1(areg[7]), .s(x2) );
  mul_mux2 sh_5_ ( .z(ain[5]), .d0(areg[5]), .d1(areg[6]), .s(x2) );
  mul_csa42 sc3_68_ ( .sum(s3[68]), .carry(c3[68]), .a(1'b0), .b(s2[68]), .c(
        c2[67]), .d(1'b0), .cin(co[67]) );
  mul_csa42 sc3_67_ ( .sum(s3[67]), .carry(c3[67]), .cout(co[67]), .a(s1[67]), 
        .b(s2[67]), .c(c2[66]), .d(1'b0), .cin(co[66]) );
  mul_csa42 sc3_66_ ( .sum(s3[66]), .carry(c3[66]), .cout(co[66]), .a(s1[66]), 
        .b(s2[66]), .c(c2[65]), .d(c1[65]), .cin(co[65]) );
  mul_csa42 sc3_65_ ( .sum(s3[65]), .carry(c3[65]), .cout(co[65]), .a(s1[65]), 
        .b(s2[65]), .c(c2[64]), .d(c1[64]), .cin(co[64]) );
  mul_csa42 sc3_64_ ( .sum(s3[64]), .carry(c3[64]), .cout(co[64]), .a(s1[64]), 
        .b(s2[64]), .c(c2[63]), .d(c1[63]), .cin(co[63]) );
  mul_csa42 sc3_63_ ( .sum(s3[63]), .carry(c3[63]), .cout(co[63]), .a(s1[63]), 
        .b(s2[63]), .c(c2[62]), .d(c1[62]), .cin(co[62]) );
  mul_csa42 sc3_62_ ( .sum(s3[62]), .carry(c3[62]), .cout(co[62]), .a(s1[62]), 
        .b(s2[62]), .c(c2[61]), .d(c1[61]), .cin(co[61]) );
  mul_csa42 sc3_61_ ( .sum(s3[61]), .carry(c3[61]), .cout(co[61]), .a(s1[61]), 
        .b(s2[61]), .c(c2[60]), .d(c1[60]), .cin(co[60]) );
  mul_csa42 sc3_60_ ( .sum(s3[60]), .carry(c3[60]), .cout(co[60]), .a(s1[60]), 
        .b(s2[60]), .c(c2[59]), .d(c1[59]), .cin(co[59]) );
  mul_csa42 sc3_59_ ( .sum(s3[59]), .carry(c3[59]), .cout(co[59]), .a(s1[59]), 
        .b(s2[59]), .c(c2[58]), .d(c1[58]), .cin(co[58]) );
  mul_csa42 sc3_58_ ( .sum(s3[58]), .carry(c3[58]), .cout(co[58]), .a(s1[58]), 
        .b(s2[58]), .c(c2[57]), .d(c1[57]), .cin(co[57]) );
  mul_csa42 sc3_57_ ( .sum(s3[57]), .carry(c3[57]), .cout(co[57]), .a(s1[57]), 
        .b(s2[57]), .c(c2[56]), .d(c1[56]), .cin(co[56]) );
  mul_csa42 sc3_56_ ( .sum(s3[56]), .carry(c3[56]), .cout(co[56]), .a(s1[56]), 
        .b(s2[56]), .c(c2[55]), .d(c1[55]), .cin(co[55]) );
  mul_csa42 sc3_55_ ( .sum(s3[55]), .carry(c3[55]), .cout(co[55]), .a(s1[55]), 
        .b(s2[55]), .c(c2[54]), .d(c1[54]), .cin(co[54]) );
  mul_csa42 sc3_54_ ( .sum(s3[54]), .carry(c3[54]), .cout(co[54]), .a(s1[54]), 
        .b(s2[54]), .c(c2[53]), .d(c1[53]), .cin(co[53]) );
  mul_csa42 sc3_53_ ( .sum(s3[53]), .carry(c3[53]), .cout(co[53]), .a(s1[53]), 
        .b(s2[53]), .c(c2[52]), .d(c1[52]), .cin(co[52]) );
  mul_csa42 sc3_52_ ( .sum(s3[52]), .carry(c3[52]), .cout(co[52]), .a(s1[52]), 
        .b(s2[52]), .c(c2[51]), .d(c1[51]), .cin(co[51]) );
  mul_csa42 sc3_51_ ( .sum(s3[51]), .carry(c3[51]), .cout(co[51]), .a(s1[51]), 
        .b(s2[51]), .c(c2[50]), .d(c1[50]), .cin(co[50]) );
  mul_csa42 sc3_50_ ( .sum(s3[50]), .carry(c3[50]), .cout(co[50]), .a(s1[50]), 
        .b(s2[50]), .c(c2[49]), .d(c1[49]), .cin(co[49]) );
  mul_csa42 sc3_49_ ( .sum(s3[49]), .carry(c3[49]), .cout(co[49]), .a(s1[49]), 
        .b(s2[49]), .c(c2[48]), .d(c1[48]), .cin(co[48]) );
  mul_csa42 sc3_48_ ( .sum(s3[48]), .carry(c3[48]), .cout(co[48]), .a(s1[48]), 
        .b(s2[48]), .c(c2[47]), .d(c1[47]), .cin(co[47]) );
  mul_csa42 sc3_47_ ( .sum(s3[47]), .carry(c3[47]), .cout(co[47]), .a(s1[47]), 
        .b(s2[47]), .c(c2[46]), .d(c1[46]), .cin(co[46]) );
  mul_csa42 sc3_46_ ( .sum(s3[46]), .carry(c3[46]), .cout(co[46]), .a(s1[46]), 
        .b(s2[46]), .c(c2[45]), .d(c1[45]), .cin(co[45]) );
  mul_csa42 sc3_45_ ( .sum(s3[45]), .carry(c3[45]), .cout(co[45]), .a(s1[45]), 
        .b(s2[45]), .c(c2[44]), .d(c1[44]), .cin(co[44]) );
  mul_csa42 sc3_44_ ( .sum(s3[44]), .carry(c3[44]), .cout(co[44]), .a(s1[44]), 
        .b(s2[44]), .c(c2[43]), .d(c1[43]), .cin(co[43]) );
  mul_csa42 sc3_43_ ( .sum(s3[43]), .carry(c3[43]), .cout(co[43]), .a(s1[43]), 
        .b(s2[43]), .c(c2[42]), .d(c1[42]), .cin(co[42]) );
  mul_csa42 sc3_42_ ( .sum(s3[42]), .carry(c3[42]), .cout(co[42]), .a(s1[42]), 
        .b(s2[42]), .c(c2[41]), .d(c1[41]), .cin(co[41]) );
  mul_csa42 sc3_41_ ( .sum(s3[41]), .carry(c3[41]), .cout(co[41]), .a(s1[41]), 
        .b(s2[41]), .c(c2[40]), .d(c1[40]), .cin(co[40]) );
  mul_csa42 sc3_40_ ( .sum(s3[40]), .carry(c3[40]), .cout(co[40]), .a(s1[40]), 
        .b(s2[40]), .c(c2[39]), .d(c1[39]), .cin(co[39]) );
  mul_csa42 sc3_39_ ( .sum(s3[39]), .carry(c3[39]), .cout(co[39]), .a(s1[39]), 
        .b(s2[39]), .c(c2[38]), .d(c1[38]), .cin(co[38]) );
  mul_csa42 sc3_38_ ( .sum(s3[38]), .carry(c3[38]), .cout(co[38]), .a(s1[38]), 
        .b(s2[38]), .c(c2[37]), .d(c1[37]), .cin(co[37]) );
  mul_csa42 sc3_37_ ( .sum(s3[37]), .carry(c3[37]), .cout(co[37]), .a(s1[37]), 
        .b(s2[37]), .c(c2[36]), .d(c1[36]), .cin(co[36]) );
  mul_csa42 sc3_36_ ( .sum(s3[36]), .carry(c3[36]), .cout(co[36]), .a(s1[36]), 
        .b(s2[36]), .c(c2[35]), .d(c1[35]), .cin(co[35]) );
  mul_csa42 sc3_35_ ( .sum(s3[35]), .carry(c3[35]), .cout(co[35]), .a(s1[35]), 
        .b(s2[35]), .c(c2[34]), .d(c1[34]), .cin(co[34]) );
  mul_csa42 sc3_34_ ( .sum(s3[34]), .carry(c3[34]), .cout(co[34]), .a(s1[34]), 
        .b(s2[34]), .c(c2[33]), .d(c1[33]), .cin(co[33]) );
  mul_csa42 sc3_33_ ( .sum(s3[33]), .carry(c3[33]), .cout(co[33]), .a(s1[33]), 
        .b(s2[33]), .c(c2[32]), .d(c1[32]), .cin(co[32]) );
  mul_csa42 sc3_32_ ( .sum(s3[32]), .carry(c3[32]), .cout(co[32]), .a(s1[32]), 
        .b(s2[32]), .c(c2[31]), .d(c1[31]), .cin(co[31]) );
  mul_csa42 sc3_31_ ( .sum(s3[31]), .carry(c3[31]), .cout(co[31]), .a(s1[31]), 
        .b(s2[31]), .c(c2[30]), .d(c1[30]), .cin(co[30]) );
  mul_csa42 sc3_30_ ( .sum(s3[30]), .carry(c3[30]), .cout(co[30]), .a(s1[30]), 
        .b(s2[30]), .c(c2[29]), .d(c1[29]), .cin(co[29]) );
  mul_csa42 sc3_29_ ( .sum(s3[29]), .carry(c3[29]), .cout(co[29]), .a(s1[29]), 
        .b(s2[29]), .c(c2[28]), .d(c1[28]), .cin(co[28]) );
  mul_csa42 sc3_28_ ( .sum(s3[28]), .carry(c3[28]), .cout(co[28]), .a(s1[28]), 
        .b(s2[28]), .c(c2[27]), .d(c1[27]), .cin(co[27]) );
  mul_csa42 sc3_27_ ( .sum(s3[27]), .carry(c3[27]), .cout(co[27]), .a(s1[27]), 
        .b(s2[27]), .c(c2[26]), .d(c1[26]), .cin(co[26]) );
  mul_csa42 sc3_26_ ( .sum(s3[26]), .carry(c3[26]), .cout(co[26]), .a(s1[26]), 
        .b(s2[26]), .c(c2[25]), .d(c1[25]), .cin(co[25]) );
  mul_csa42 sc3_25_ ( .sum(s3[25]), .carry(c3[25]), .cout(co[25]), .a(s1[25]), 
        .b(s2[25]), .c(c2[24]), .d(c1[24]), .cin(co[24]) );
  mul_csa42 sc3_24_ ( .sum(s3[24]), .carry(c3[24]), .cout(co[24]), .a(s1[24]), 
        .b(s2[24]), .c(c2[23]), .d(c1[23]), .cin(co[23]) );
  mul_csa42 sc3_23_ ( .sum(s3[23]), .carry(c3[23]), .cout(co[23]), .a(s1[23]), 
        .b(s2[23]), .c(c2[22]), .d(c1[22]), .cin(co[22]) );
  mul_csa42 sc3_22_ ( .sum(s3[22]), .carry(c3[22]), .cout(co[22]), .a(s1[22]), 
        .b(s2[22]), .c(c2[21]), .d(c1[21]), .cin(co[21]) );
  mul_csa42 sc3_21_ ( .sum(s3[21]), .carry(c3[21]), .cout(co[21]), .a(s1[21]), 
        .b(s2[21]), .c(c2[20]), .d(c1[20]), .cin(co[20]) );
  mul_csa42 sc3_20_ ( .sum(s3[20]), .carry(c3[20]), .cout(co[20]), .a(s1[20]), 
        .b(s2[20]), .c(c2[19]), .d(c1[19]), .cin(1'b0) );
  mul_csa32 sc4_82_ ( .sum(psum[82]), .cout(pcout[82]), .a(ain[82]), .b(s2[82]), .c(c3[81]) );
  mul_csa32 sc4_68_ ( .sum(psum[68]), .cout(pcout[68]), .a(ain[68]), .b(s3[68]), .c(c3[67]) );
  mul_csa32 sc4_67_ ( .sum(psum[67]), .cout(pcout[67]), .a(ain[67]), .b(s3[67]), .c(c3[66]) );
  mul_csa32 sc4_66_ ( .sum(psum[66]), .cout(pcout[66]), .a(ain[66]), .b(s3[66]), .c(c3[65]) );
  mul_csa32 sc4_65_ ( .sum(psum[65]), .cout(pcout[65]), .a(ain[65]), .b(s3[65]), .c(c3[64]) );
  mul_csa32 sc4_64_ ( .sum(psum[64]), .cout(pcout[64]), .a(ain[64]), .b(s3[64]), .c(c3[63]) );
  mul_csa32 sc4_63_ ( .sum(psum[63]), .cout(pcout[63]), .a(ain[63]), .b(s3[63]), .c(c3[62]) );
  mul_csa32 sc4_62_ ( .sum(psum[62]), .cout(pcout[62]), .a(ain[62]), .b(s3[62]), .c(c3[61]) );
  mul_csa32 sc4_61_ ( .sum(psum[61]), .cout(pcout[61]), .a(ain[61]), .b(s3[61]), .c(c3[60]) );
  mul_csa32 sc4_60_ ( .sum(psum[60]), .cout(pcout[60]), .a(ain[60]), .b(s3[60]), .c(c3[59]) );
  mul_csa32 sc4_59_ ( .sum(psum[59]), .cout(pcout[59]), .a(ain[59]), .b(s3[59]), .c(c3[58]) );
  mul_csa32 sc4_58_ ( .sum(psum[58]), .cout(pcout[58]), .a(ain[58]), .b(s3[58]), .c(c3[57]) );
  mul_csa32 sc4_57_ ( .sum(psum[57]), .cout(pcout[57]), .a(ain[57]), .b(s3[57]), .c(c3[56]) );
  mul_csa32 sc4_56_ ( .sum(psum[56]), .cout(pcout[56]), .a(ain[56]), .b(s3[56]), .c(c3[55]) );
  mul_csa32 sc4_55_ ( .sum(psum[55]), .cout(pcout[55]), .a(ain[55]), .b(s3[55]), .c(c3[54]) );
  mul_csa32 sc4_54_ ( .sum(psum[54]), .cout(pcout[54]), .a(ain[54]), .b(s3[54]), .c(c3[53]) );
  mul_csa32 sc4_53_ ( .sum(psum[53]), .cout(pcout[53]), .a(ain[53]), .b(s3[53]), .c(c3[52]) );
  mul_csa32 sc4_52_ ( .sum(psum[52]), .cout(pcout[52]), .a(ain[52]), .b(s3[52]), .c(c3[51]) );
  mul_csa32 sc4_51_ ( .sum(psum[51]), .cout(pcout[51]), .a(ain[51]), .b(s3[51]), .c(c3[50]) );
  mul_csa32 sc4_50_ ( .sum(psum[50]), .cout(pcout[50]), .a(ain[50]), .b(s3[50]), .c(c3[49]) );
  mul_csa32 sc4_49_ ( .sum(psum[49]), .cout(pcout[49]), .a(ain[49]), .b(s3[49]), .c(c3[48]) );
  mul_csa32 sc4_48_ ( .sum(psum[48]), .cout(pcout[48]), .a(ain[48]), .b(s3[48]), .c(c3[47]) );
  mul_csa32 sc4_47_ ( .sum(psum[47]), .cout(pcout[47]), .a(ain[47]), .b(s3[47]), .c(c3[46]) );
  mul_csa32 sc4_46_ ( .sum(psum[46]), .cout(pcout[46]), .a(ain[46]), .b(s3[46]), .c(c3[45]) );
  mul_csa32 sc4_45_ ( .sum(psum[45]), .cout(pcout[45]), .a(ain[45]), .b(s3[45]), .c(c3[44]) );
  mul_csa32 sc4_44_ ( .sum(psum[44]), .cout(pcout[44]), .a(ain[44]), .b(s3[44]), .c(c3[43]) );
  mul_csa32 sc4_43_ ( .sum(psum[43]), .cout(pcout[43]), .a(ain[43]), .b(s3[43]), .c(c3[42]) );
  mul_csa32 sc4_42_ ( .sum(psum[42]), .cout(pcout[42]), .a(ain[42]), .b(s3[42]), .c(c3[41]) );
  mul_csa32 sc4_41_ ( .sum(psum[41]), .cout(pcout[41]), .a(ain[41]), .b(s3[41]), .c(c3[40]) );
  mul_csa32 sc4_40_ ( .sum(psum[40]), .cout(pcout[40]), .a(ain[40]), .b(s3[40]), .c(c3[39]) );
  mul_csa32 sc4_39_ ( .sum(psum[39]), .cout(pcout[39]), .a(ain[39]), .b(s3[39]), .c(c3[38]) );
  mul_csa32 sc4_38_ ( .sum(psum[38]), .cout(pcout[38]), .a(ain[38]), .b(s3[38]), .c(c3[37]) );
  mul_csa32 sc4_37_ ( .sum(psum[37]), .cout(pcout[37]), .a(ain[37]), .b(s3[37]), .c(c3[36]) );
  mul_csa32 sc4_36_ ( .sum(psum[36]), .cout(pcout[36]), .a(ain[36]), .b(s3[36]), .c(c3[35]) );
  mul_csa32 sc4_35_ ( .sum(psum[35]), .cout(pcout[35]), .a(ain[35]), .b(s3[35]), .c(c3[34]) );
  mul_csa32 sc4_34_ ( .sum(psum[34]), .cout(pcout[34]), .a(ain[34]), .b(s3[34]), .c(c3[33]) );
  mul_csa32 sc4_33_ ( .sum(psum[33]), .cout(pcout[33]), .a(ain[33]), .b(s3[33]), .c(c3[32]) );
  mul_csa32 sc4_32_ ( .sum(psum[32]), .cout(pcout[32]), .a(ain[32]), .b(s3[32]), .c(c3[31]) );
  mul_csa32 sc4_31_ ( .sum(psum[31]), .cout(pcout[31]), .a(ain[31]), .b(s3[31]), .c(c3[30]) );
  mul_csa32 sc4_30_ ( .sum(psum[30]), .cout(pcout[30]), .a(ain[30]), .b(s3[30]), .c(c3[29]) );
  mul_csa32 sc4_29_ ( .sum(psum[29]), .cout(pcout[29]), .a(ain[29]), .b(s3[29]), .c(c3[28]) );
  mul_csa32 sc4_28_ ( .sum(psum[28]), .cout(pcout[28]), .a(ain[28]), .b(s3[28]), .c(c3[27]) );
  mul_csa32 sc4_27_ ( .sum(psum[27]), .cout(pcout[27]), .a(ain[27]), .b(s3[27]), .c(c3[26]) );
  mul_csa32 sc4_26_ ( .sum(psum[26]), .cout(pcout[26]), .a(ain[26]), .b(s3[26]), .c(c3[25]) );
  mul_csa32 sc4_25_ ( .sum(psum[25]), .cout(pcout[25]), .a(ain[25]), .b(s3[25]), .c(c3[24]) );
  mul_csa32 sc4_24_ ( .sum(psum[24]), .cout(pcout[24]), .a(ain[24]), .b(s3[24]), .c(c3[23]) );
  mul_csa32 sc4_23_ ( .sum(psum[23]), .cout(pcout[23]), .a(ain[23]), .b(s3[23]), .c(c3[22]) );
  mul_csa32 sc4_22_ ( .sum(psum[22]), .cout(pcout[22]), .a(ain[22]), .b(s3[22]), .c(c3[21]) );
  mul_csa32 sc4_21_ ( .sum(psum[21]), .cout(pcout[21]), .a(ain[21]), .b(s3[21]), .c(c3[20]) );
  mul_csa32 sc4_20_ ( .sum(psum[20]), .cout(pcout[20]), .a(ain[20]), .b(s3[20]), .c(c3[19]) );
  mul_csa32 sc4_96_ ( .sum(psum[96]), .cout(pcout[96]), .a(ain[96]), .b(s2[96]), .c(c2[95]) );
  mul_csa32 sc4_95_ ( .sum(psum[95]), .cout(pcout[95]), .a(ain[95]), .b(s2[95]), .c(c2[94]) );
  mul_csa32 sc4_94_ ( .sum(psum[94]), .cout(pcout[94]), .a(ain[94]), .b(s2[94]), .c(c2[93]) );
  mul_csa32 sc4_93_ ( .sum(psum[93]), .cout(pcout[93]), .a(ain[93]), .b(s2[93]), .c(c2[92]) );
  mul_csa32 sc4_92_ ( .sum(psum[92]), .cout(pcout[92]), .a(ain[92]), .b(s2[92]), .c(c2[91]) );
  mul_csa32 sc4_91_ ( .sum(psum[91]), .cout(pcout[91]), .a(ain[91]), .b(s2[91]), .c(c2[90]) );
  mul_csa32 sc4_90_ ( .sum(psum[90]), .cout(pcout[90]), .a(ain[90]), .b(s2[90]), .c(c2[89]) );
  mul_csa32 sc4_89_ ( .sum(psum[89]), .cout(pcout[89]), .a(ain[89]), .b(s2[89]), .c(c2[88]) );
  mul_csa32 sc4_88_ ( .sum(psum[88]), .cout(pcout[88]), .a(ain[88]), .b(s2[88]), .c(c2[87]) );
  mul_csa32 sc4_87_ ( .sum(psum[87]), .cout(pcout[87]), .a(ain[87]), .b(s2[87]), .c(c2[86]) );
  mul_csa32 sc4_86_ ( .sum(psum[86]), .cout(pcout[86]), .a(ain[86]), .b(s2[86]), .c(c2[85]) );
  mul_csa32 sc4_85_ ( .sum(psum[85]), .cout(pcout[85]), .a(ain[85]), .b(s2[85]), .c(c2[84]) );
  mul_csa32 sc4_84_ ( .sum(psum[84]), .cout(pcout[84]), .a(ain[84]), .b(s2[84]), .c(c2[83]) );
  mul_csa32 sc4_81_ ( .sum(psum[81]), .cout(pcout[81]), .a(ain[81]), .b(s3[81]), .c(c3[80]) );
  mul_csa32 sc4_80_ ( .sum(psum[80]), .cout(pcout[80]), .a(ain[80]), .b(s3[80]), .c(c3[79]) );
  mul_csa32 sc4_79_ ( .sum(psum[79]), .cout(pcout[79]), .a(ain[79]), .b(s3[79]), .c(c3[78]) );
  mul_csa32 sc4_78_ ( .sum(psum[78]), .cout(pcout[78]), .a(ain[78]), .b(s3[78]), .c(c3[77]) );
  mul_csa32 sc4_77_ ( .sum(psum[77]), .cout(pcout[77]), .a(ain[77]), .b(s3[77]), .c(c3[76]) );
  mul_csa32 sc4_76_ ( .sum(psum[76]), .cout(pcout[76]), .a(ain[76]), .b(s3[76]), .c(c3[75]) );
  mul_csa32 sc4_75_ ( .sum(psum[75]), .cout(pcout[75]), .a(ain[75]), .b(s3[75]), .c(c3[74]) );
  mul_csa32 sc4_74_ ( .sum(psum[74]), .cout(pcout[74]), .a(ain[74]), .b(s3[74]), .c(c3[73]) );
  mul_csa32 sc4_73_ ( .sum(psum[73]), .cout(pcout[73]), .a(ain[73]), .b(s3[73]), .c(c3[72]) );
  mul_csa32 sc4_72_ ( .sum(psum[72]), .cout(pcout[72]), .a(ain[72]), .b(s3[72]), .c(c3[71]) );
  mul_csa32 sc4_71_ ( .sum(psum[71]), .cout(pcout[71]), .a(ain[71]), .b(s3[71]), .c(c3[70]) );
  mul_csa32 sc4_70_ ( .sum(psum[70]), .cout(pcout[70]), .a(ain[70]), .b(s3[70]), .c(c3[69]) );
  mul_csa32 sc4_69_ ( .sum(psum[69]), .cout(pcout[69]), .a(ain[69]), .b(s3[69]), .c(c3[68]) );
  mul_csa32 acc_4_ ( .sum(psum[4]), .cout(pcout[4]), .a(ain[4]), .b(s2[4]), 
        .c(c2[3]) );
  mul_csa32 acc_3_ ( .sum(psum[3]), .cout(pcout[3]), .a(ain[3]), .b(s2[3]), 
        .c(c2[2]) );
  mul_csa32 acc_2_ ( .sum(psum[2]), .cout(pcout[2]), .a(ain[2]), .b(s2[2]), 
        .c(c2[1]) );
  mul_csa32 acc_1_ ( .sum(psum[1]), .cout(pcout[1]), .a(ain[1]), .b(s2[1]), 
        .c(c2[0]) );
  mul_csa32 sc3_97_ ( .sum(psum[97]), .cout(pcout[97]), .a(a1s[81]), .b(
        a1c[80]), .c(c2[96]) );
  mul_csa32 sc1_19_ ( .sum(s1[19]), .cout(c1[19]), .a(ps[51]), .b(pc[50]), .c(
        a1s[3]) );
  mul_csa32 sc1_18_ ( .sum(s1[18]), .cout(c1[18]), .a(ps[50]), .b(pc[49]), .c(
        a1s[2]) );
  mul_csa32 sc1_17_ ( .sum(s1[17]), .cout(c1[17]), .a(ps[49]), .b(pc[48]), .c(
        a1s[1]) );
  mul_csa32 sc1_16_ ( .sum(s1[16]), .cout(c1[16]), .a(ps[48]), .b(pc[47]), .c(
        a1s[0]) );
  mul_csa32 sc1_15_ ( .sum(s1[15]), .cout(c1[15]), .a(ps[47]), .b(pc[46]), .c(
        1'b0) );
  mul_csa32 sc4_83_ ( .sum(psum[83]), .cout(pcout[83]), .a(ain[83]), .b(s2[83]), .c(c2[82]) );
  mul_csa32 sc2_83_ ( .sum(s2[83]), .cout(c2[83]), .a(a1s[67]), .b(a1c[66]), 
        .c(c1[82]) );
  mul_csa32 sc2_19_ ( .sum(s2[19]), .cout(c2[19]), .a(s1[19]), .b(a0s[19]), 
        .c(a0c[18]) );
  mul_csa32 sc2_18_ ( .sum(s2[18]), .cout(c2[18]), .a(s1[18]), .b(a0s[18]), 
        .c(a0c[17]) );
  mul_csa32 sc2_17_ ( .sum(s2[17]), .cout(c2[17]), .a(s1[17]), .b(a0s[17]), 
        .c(a0c[16]) );
  mul_csa32 sc2_16_ ( .sum(s2[16]), .cout(c2[16]), .a(s1[16]), .b(a0s[16]), 
        .c(a0c[15]) );
  mul_csa32 sc2_15_ ( .sum(s2[15]), .cout(c2[15]), .a(s1[15]), .b(a0s[15]), 
        .c(a0c[14]) );
  mul_csa32 sc1_81_ ( .sum(s1[81]), .cout(c1[81]), .a(a1s[65]), .b(a1c[64]), 
        .c(a0s[81]) );
  mul_csa32 sc1_80_ ( .sum(s1[80]), .cout(c1[80]), .a(a1s[64]), .b(a1c[63]), 
        .c(a0s[80]) );
  mul_csa32 sc1_79_ ( .sum(s1[79]), .cout(c1[79]), .a(a1s[63]), .b(a1c[62]), 
        .c(a0s[79]) );
  mul_csa32 sc1_78_ ( .sum(s1[78]), .cout(c1[78]), .a(a1s[62]), .b(a1c[61]), 
        .c(a0s[78]) );
  mul_csa32 sc1_77_ ( .sum(s1[77]), .cout(c1[77]), .a(a1s[61]), .b(a1c[60]), 
        .c(a0s[77]) );
  mul_csa32 sc1_76_ ( .sum(s1[76]), .cout(c1[76]), .a(a1s[60]), .b(a1c[59]), 
        .c(a0s[76]) );
  mul_csa32 sc1_75_ ( .sum(s1[75]), .cout(c1[75]), .a(a1s[59]), .b(a1c[58]), 
        .c(a0s[75]) );
  mul_csa32 sc1_74_ ( .sum(s1[74]), .cout(c1[74]), .a(a1s[58]), .b(a1c[57]), 
        .c(a0s[74]) );
  mul_csa32 sc1_73_ ( .sum(s1[73]), .cout(c1[73]), .a(a1s[57]), .b(a1c[56]), 
        .c(a0s[73]) );
  mul_csa32 sc1_72_ ( .sum(s1[72]), .cout(c1[72]), .a(a1s[56]), .b(a1c[55]), 
        .c(a0s[72]) );
  mul_csa32 sc1_71_ ( .sum(s1[71]), .cout(c1[71]), .a(a1s[55]), .b(a1c[54]), 
        .c(a0s[71]) );
  mul_csa32 sc1_70_ ( .sum(s1[70]), .cout(c1[70]), .a(a1s[54]), .b(a1c[53]), 
        .c(a0s[70]) );
  mul_csa32 sc1_69_ ( .sum(s1[69]), .cout(c1[69]), .a(a1s[53]), .b(a1c[52]), 
        .c(a0s[69]) );
  mul_csa32 sc1_68_ ( .sum(s1[68]), .cout(c1[68]), .a(a1s[52]), .b(a1c[51]), 
        .c(a0s[68]) );
  mul_csa32 sc3_19_ ( .sum(s3[19]), .cout(c3[19]), .a(s2[19]), .b(c1[18]), .c(
        c2[18]) );
  mul_csa32 sc3_18_ ( .sum(s3[18]), .cout(c3[18]), .a(s2[18]), .b(c1[17]), .c(
        c2[17]) );
  mul_csa32 sc3_17_ ( .sum(s3[17]), .cout(c3[17]), .a(s2[17]), .b(c1[16]), .c(
        c2[16]) );
  mul_csa32 sc3_16_ ( .sum(s3[16]), .cout(c3[16]), .a(s2[16]), .b(c1[15]), .c(
        c2[15]) );
  mul_csa32 sc3_15_ ( .sum(s3[15]), .cout(c3[15]), .a(s2[15]), .b(c1[14]), .c(
        c2[14]) );
  mul_csa32 sc1_82_ ( .sum(s1[82]), .cout(c1[82]), .a(a1s[66]), .b(a1c[65]), 
        .c(a0c[81]) );
  mul_csa32 acc_14_ ( .sum(psum[14]), .cout(pcout[14]), .a(ain[14]), .b(s2[14]), .c(c2[13]) );
  mul_csa32 acc_13_ ( .sum(psum[13]), .cout(pcout[13]), .a(ain[13]), .b(s2[13]), .c(c2[12]) );
  mul_csa32 acc_12_ ( .sum(psum[12]), .cout(pcout[12]), .a(ain[12]), .b(s2[12]), .c(c2[11]) );
  mul_csa32 acc_11_ ( .sum(psum[11]), .cout(pcout[11]), .a(ain[11]), .b(s2[11]), .c(c2[10]) );
  mul_csa32 acc_10_ ( .sum(psum[10]), .cout(pcout[10]), .a(ain[10]), .b(s2[10]), .c(c2[9]) );
  mul_csa32 acc_9_ ( .sum(psum[9]), .cout(pcout[9]), .a(ain[9]), .b(s2[9]), 
        .c(c2[8]) );
  mul_csa32 acc_8_ ( .sum(psum[8]), .cout(pcout[8]), .a(ain[8]), .b(s2[8]), 
        .c(c2[7]) );
  mul_csa32 acc_7_ ( .sum(psum[7]), .cout(pcout[7]), .a(ain[7]), .b(s2[7]), 
        .c(c2[6]) );
  mul_csa32 acc_6_ ( .sum(psum[6]), .cout(pcout[6]), .a(ain[6]), .b(s2[6]), 
        .c(c2[5]) );
  mul_csa32 acc_5_ ( .sum(psum[5]), .cout(pcout[5]), .a(ain[5]), .b(s2[5]), 
        .c(c2[4]) );
  mul_csa32 sc2_67_ ( .sum(s2[67]), .cout(c2[67]), .a(a0s[67]), .b(c1[66]), 
        .c(a0c[66]) );
  mul_csa32 sc1_14_ ( .sum(s1[14]), .cout(c1[14]), .a(ps[46]), .b(pc[45]), .c(
        a0s[14]) );
  mul_csa32 sc1_13_ ( .sum(s1[13]), .cout(c1[13]), .a(ps[45]), .b(pc[44]), .c(
        a0s[13]) );
  mul_csa32 sc1_12_ ( .sum(s1[12]), .cout(c1[12]), .a(ps[44]), .b(pc[43]), .c(
        a0s[12]) );
  mul_csa32 sc1_11_ ( .sum(s1[11]), .cout(c1[11]), .a(ps[43]), .b(pc[42]), .c(
        a0s[11]) );
  mul_csa32 sc1_10_ ( .sum(s1[10]), .cout(c1[10]), .a(ps[42]), .b(pc[41]), .c(
        a0s[10]) );
  mul_csa32 sc1_9_ ( .sum(s1[9]), .cout(c1[9]), .a(ps[41]), .b(pc[40]), .c(
        a0s[9]) );
  mul_csa32 sc1_8_ ( .sum(s1[8]), .cout(c1[8]), .a(ps[40]), .b(pc[39]), .c(
        a0s[8]) );
  mul_csa32 sc1_7_ ( .sum(s1[7]), .cout(c1[7]), .a(ps[39]), .b(pc[38]), .c(
        a0s[7]) );
  mul_csa32 sc1_6_ ( .sum(s1[6]), .cout(c1[6]), .a(ps[38]), .b(pc[37]), .c(
        a0s[6]) );
  mul_csa32 sc1_5_ ( .sum(s1[5]), .cout(c1[5]), .a(ps[37]), .b(pc[36]), .c(
        a0s[5]) );
  mul_csa32 sc2_14_ ( .sum(s2[14]), .cout(c2[14]), .a(s1[14]), .b(c1[13]), .c(
        a0c[13]) );
  mul_csa32 sc2_13_ ( .sum(s2[13]), .cout(c2[13]), .a(s1[13]), .b(c1[12]), .c(
        a0c[12]) );
  mul_csa32 sc2_12_ ( .sum(s2[12]), .cout(c2[12]), .a(s1[12]), .b(c1[11]), .c(
        a0c[11]) );
  mul_csa32 sc2_11_ ( .sum(s2[11]), .cout(c2[11]), .a(s1[11]), .b(c1[10]), .c(
        a0c[10]) );
  mul_csa32 sc2_10_ ( .sum(s2[10]), .cout(c2[10]), .a(s1[10]), .b(c1[9]), .c(
        a0c[9]) );
  mul_csa32 sc2_9_ ( .sum(s2[9]), .cout(c2[9]), .a(s1[9]), .b(c1[8]), .c(
        a0c[8]) );
  mul_csa32 sc2_8_ ( .sum(s2[8]), .cout(c2[8]), .a(s1[8]), .b(c1[7]), .c(
        a0c[7]) );
  mul_csa32 sc2_7_ ( .sum(s2[7]), .cout(c2[7]), .a(s1[7]), .b(c1[6]), .c(
        a0c[6]) );
  mul_csa32 sc2_6_ ( .sum(s2[6]), .cout(c2[6]), .a(s1[6]), .b(c1[5]), .c(
        a0c[5]) );
  mul_csa32 sc2_5_ ( .sum(s2[5]), .cout(c2[5]), .a(s1[5]), .b(c1[4]), .c(
        a0c[4]) );
  mul_csa32 sc2_82_ ( .sum(s2[82]), .cout(c2[82]), .a(s1[82]), .b(c1[81]), .c(
        c2[81]) );
  mul_csa32 sc1_4_ ( .sum(s1[4]), .cout(c1[4]), .a(ps[36]), .b(pc[35]), .c(
        a0s[4]) );
  mul_csa32 sc1_3_ ( .sum(s1[3]), .cout(c1[3]), .a(ps[35]), .b(pc[34]), .c(
        a0s[3]) );
  mul_csa32 sc1_2_ ( .sum(s1[2]), .cout(c1[2]), .a(ps[34]), .b(pc[33]), .c(
        a0s[2]) );
  mul_csa32 sc1_1_ ( .sum(s1[1]), .cout(c1[1]), .a(ps[33]), .b(pc[32]), .c(
        a0s[1]) );
  mul_csa32 sc2_66_ ( .sum(s2[66]), .cout(c2[66]), .a(a1c[49]), .b(a0s[66]), 
        .c(a0c[65]) );
  mul_csa32 sc2_65_ ( .sum(s2[65]), .cout(c2[65]), .a(a1c[48]), .b(a0s[65]), 
        .c(a0c[64]) );
  mul_csa32 sc2_64_ ( .sum(s2[64]), .cout(c2[64]), .a(a1c[47]), .b(a0s[64]), 
        .c(a0c[63]) );
  mul_csa32 sc2_63_ ( .sum(s2[63]), .cout(c2[63]), .a(a1c[46]), .b(a0s[63]), 
        .c(a0c[62]) );
  mul_csa32 sc2_62_ ( .sum(s2[62]), .cout(c2[62]), .a(a1c[45]), .b(a0s[62]), 
        .c(a0c[61]) );
  mul_csa32 sc2_61_ ( .sum(s2[61]), .cout(c2[61]), .a(a1c[44]), .b(a0s[61]), 
        .c(a0c[60]) );
  mul_csa32 sc2_60_ ( .sum(s2[60]), .cout(c2[60]), .a(a1c[43]), .b(a0s[60]), 
        .c(a0c[59]) );
  mul_csa32 sc2_59_ ( .sum(s2[59]), .cout(c2[59]), .a(a1c[42]), .b(a0s[59]), 
        .c(a0c[58]) );
  mul_csa32 sc2_58_ ( .sum(s2[58]), .cout(c2[58]), .a(a1c[41]), .b(a0s[58]), 
        .c(a0c[57]) );
  mul_csa32 sc2_57_ ( .sum(s2[57]), .cout(c2[57]), .a(a1c[40]), .b(a0s[57]), 
        .c(a0c[56]) );
  mul_csa32 sc2_56_ ( .sum(s2[56]), .cout(c2[56]), .a(a1c[39]), .b(a0s[56]), 
        .c(a0c[55]) );
  mul_csa32 sc2_55_ ( .sum(s2[55]), .cout(c2[55]), .a(a1c[38]), .b(a0s[55]), 
        .c(a0c[54]) );
  mul_csa32 sc2_54_ ( .sum(s2[54]), .cout(c2[54]), .a(a1c[37]), .b(a0s[54]), 
        .c(a0c[53]) );
  mul_csa32 sc2_53_ ( .sum(s2[53]), .cout(c2[53]), .a(a1c[36]), .b(a0s[53]), 
        .c(a0c[52]) );
  mul_csa32 sc2_52_ ( .sum(s2[52]), .cout(c2[52]), .a(a1c[35]), .b(a0s[52]), 
        .c(a0c[51]) );
  mul_csa32 sc2_51_ ( .sum(s2[51]), .cout(c2[51]), .a(a1c[34]), .b(a0s[51]), 
        .c(a0c[50]) );
  mul_csa32 sc2_50_ ( .sum(s2[50]), .cout(c2[50]), .a(a1c[33]), .b(a0s[50]), 
        .c(a0c[49]) );
  mul_csa32 sc2_49_ ( .sum(s2[49]), .cout(c2[49]), .a(a1c[32]), .b(a0s[49]), 
        .c(a0c[48]) );
  mul_csa32 sc2_48_ ( .sum(s2[48]), .cout(c2[48]), .a(a1c[31]), .b(a0s[48]), 
        .c(a0c[47]) );
  mul_csa32 sc2_47_ ( .sum(s2[47]), .cout(c2[47]), .a(a1c[30]), .b(a0s[47]), 
        .c(a0c[46]) );
  mul_csa32 sc2_46_ ( .sum(s2[46]), .cout(c2[46]), .a(a1c[29]), .b(a0s[46]), 
        .c(a0c[45]) );
  mul_csa32 sc2_45_ ( .sum(s2[45]), .cout(c2[45]), .a(a1c[28]), .b(a0s[45]), 
        .c(a0c[44]) );
  mul_csa32 sc2_44_ ( .sum(s2[44]), .cout(c2[44]), .a(a1c[27]), .b(a0s[44]), 
        .c(a0c[43]) );
  mul_csa32 sc2_43_ ( .sum(s2[43]), .cout(c2[43]), .a(a1c[26]), .b(a0s[43]), 
        .c(a0c[42]) );
  mul_csa32 sc2_42_ ( .sum(s2[42]), .cout(c2[42]), .a(a1c[25]), .b(a0s[42]), 
        .c(a0c[41]) );
  mul_csa32 sc2_41_ ( .sum(s2[41]), .cout(c2[41]), .a(a1c[24]), .b(a0s[41]), 
        .c(a0c[40]) );
  mul_csa32 sc2_40_ ( .sum(s2[40]), .cout(c2[40]), .a(a1c[23]), .b(a0s[40]), 
        .c(a0c[39]) );
  mul_csa32 sc2_39_ ( .sum(s2[39]), .cout(c2[39]), .a(a1c[22]), .b(a0s[39]), 
        .c(a0c[38]) );
  mul_csa32 sc2_38_ ( .sum(s2[38]), .cout(c2[38]), .a(a1c[21]), .b(a0s[38]), 
        .c(a0c[37]) );
  mul_csa32 sc2_37_ ( .sum(s2[37]), .cout(c2[37]), .a(a1c[20]), .b(a0s[37]), 
        .c(a0c[36]) );
  mul_csa32 sc2_36_ ( .sum(s2[36]), .cout(c2[36]), .a(a1c[19]), .b(a0s[36]), 
        .c(a0c[35]) );
  mul_csa32 sc2_35_ ( .sum(s2[35]), .cout(c2[35]), .a(a1c[18]), .b(a0s[35]), 
        .c(a0c[34]) );
  mul_csa32 sc2_34_ ( .sum(s2[34]), .cout(c2[34]), .a(a1c[17]), .b(a0s[34]), 
        .c(a0c[33]) );
  mul_csa32 sc2_33_ ( .sum(s2[33]), .cout(c2[33]), .a(a1c[16]), .b(a0s[33]), 
        .c(a0c[32]) );
  mul_csa32 sc2_32_ ( .sum(s2[32]), .cout(c2[32]), .a(a1c[15]), .b(a0s[32]), 
        .c(a0c[31]) );
  mul_csa32 sc2_31_ ( .sum(s2[31]), .cout(c2[31]), .a(a1c[14]), .b(a0s[31]), 
        .c(a0c[30]) );
  mul_csa32 sc2_30_ ( .sum(s2[30]), .cout(c2[30]), .a(a1c[13]), .b(a0s[30]), 
        .c(a0c[29]) );
  mul_csa32 sc2_29_ ( .sum(s2[29]), .cout(c2[29]), .a(a1c[12]), .b(a0s[29]), 
        .c(a0c[28]) );
  mul_csa32 sc2_28_ ( .sum(s2[28]), .cout(c2[28]), .a(a1c[11]), .b(a0s[28]), 
        .c(a0c[27]) );
  mul_csa32 sc2_27_ ( .sum(s2[27]), .cout(c2[27]), .a(a1c[10]), .b(a0s[27]), 
        .c(a0c[26]) );
  mul_csa32 sc2_26_ ( .sum(s2[26]), .cout(c2[26]), .a(a1c[9]), .b(a0s[26]), 
        .c(a0c[25]) );
  mul_csa32 sc2_25_ ( .sum(s2[25]), .cout(c2[25]), .a(a1c[8]), .b(a0s[25]), 
        .c(a0c[24]) );
  mul_csa32 sc2_24_ ( .sum(s2[24]), .cout(c2[24]), .a(a1c[7]), .b(a0s[24]), 
        .c(a0c[23]) );
  mul_csa32 sc2_23_ ( .sum(s2[23]), .cout(c2[23]), .a(a1c[6]), .b(a0s[23]), 
        .c(a0c[22]) );
  mul_csa32 sc2_22_ ( .sum(s2[22]), .cout(c2[22]), .a(a1c[5]), .b(a0s[22]), 
        .c(a0c[21]) );
  mul_csa32 sc2_21_ ( .sum(s2[21]), .cout(c2[21]), .a(a1c[4]), .b(a0s[21]), 
        .c(a0c[20]) );
  mul_csa32 sc2_20_ ( .sum(s2[20]), .cout(c2[20]), .a(1'b0), .b(a0s[20]), .c(
        a0c[19]) );
  mul_csa32 sc1_66_ ( .sum(s1[66]), .cout(c1[66]), .a(ps[98]), .b(pc[97]), .c(
        a1s[50]) );
  mul_csa32 sc1_65_ ( .sum(s1[65]), .cout(c1[65]), .a(ps[97]), .b(pc[96]), .c(
        a1s[49]) );
  mul_csa32 sc1_64_ ( .sum(s1[64]), .cout(c1[64]), .a(ps[96]), .b(pc[95]), .c(
        a1s[48]) );
  mul_csa32 sc1_63_ ( .sum(s1[63]), .cout(c1[63]), .a(ps[95]), .b(pc[94]), .c(
        a1s[47]) );
  mul_csa32 sc1_62_ ( .sum(s1[62]), .cout(c1[62]), .a(ps[94]), .b(pc[93]), .c(
        a1s[46]) );
  mul_csa32 sc1_61_ ( .sum(s1[61]), .cout(c1[61]), .a(ps[93]), .b(pc[92]), .c(
        a1s[45]) );
  mul_csa32 sc1_60_ ( .sum(s1[60]), .cout(c1[60]), .a(ps[92]), .b(pc[91]), .c(
        a1s[44]) );
  mul_csa32 sc1_59_ ( .sum(s1[59]), .cout(c1[59]), .a(ps[91]), .b(pc[90]), .c(
        a1s[43]) );
  mul_csa32 sc1_58_ ( .sum(s1[58]), .cout(c1[58]), .a(ps[90]), .b(pc[89]), .c(
        a1s[42]) );
  mul_csa32 sc1_57_ ( .sum(s1[57]), .cout(c1[57]), .a(ps[89]), .b(pc[88]), .c(
        a1s[41]) );
  mul_csa32 sc1_56_ ( .sum(s1[56]), .cout(c1[56]), .a(ps[88]), .b(pc[87]), .c(
        a1s[40]) );
  mul_csa32 sc1_55_ ( .sum(s1[55]), .cout(c1[55]), .a(ps[87]), .b(pc[86]), .c(
        a1s[39]) );
  mul_csa32 sc1_54_ ( .sum(s1[54]), .cout(c1[54]), .a(ps[86]), .b(pc[85]), .c(
        a1s[38]) );
  mul_csa32 sc1_53_ ( .sum(s1[53]), .cout(c1[53]), .a(ps[85]), .b(pc[84]), .c(
        a1s[37]) );
  mul_csa32 sc1_52_ ( .sum(s1[52]), .cout(c1[52]), .a(ps[84]), .b(pc[83]), .c(
        a1s[36]) );
  mul_csa32 sc1_51_ ( .sum(s1[51]), .cout(c1[51]), .a(ps[83]), .b(pc[82]), .c(
        a1s[35]) );
  mul_csa32 sc1_50_ ( .sum(s1[50]), .cout(c1[50]), .a(ps[82]), .b(pc[81]), .c(
        a1s[34]) );
  mul_csa32 sc1_49_ ( .sum(s1[49]), .cout(c1[49]), .a(ps[81]), .b(pc[80]), .c(
        a1s[33]) );
  mul_csa32 sc1_48_ ( .sum(s1[48]), .cout(c1[48]), .a(ps[80]), .b(pc[79]), .c(
        a1s[32]) );
  mul_csa32 sc1_47_ ( .sum(s1[47]), .cout(c1[47]), .a(ps[79]), .b(pc[78]), .c(
        a1s[31]) );
  mul_csa32 sc1_46_ ( .sum(s1[46]), .cout(c1[46]), .a(ps[78]), .b(pc[77]), .c(
        a1s[30]) );
  mul_csa32 sc1_45_ ( .sum(s1[45]), .cout(c1[45]), .a(ps[77]), .b(pc[76]), .c(
        a1s[29]) );
  mul_csa32 sc1_44_ ( .sum(s1[44]), .cout(c1[44]), .a(ps[76]), .b(pc[75]), .c(
        a1s[28]) );
  mul_csa32 sc1_43_ ( .sum(s1[43]), .cout(c1[43]), .a(ps[75]), .b(pc[74]), .c(
        a1s[27]) );
  mul_csa32 sc1_42_ ( .sum(s1[42]), .cout(c1[42]), .a(ps[74]), .b(pc[73]), .c(
        a1s[26]) );
  mul_csa32 sc1_41_ ( .sum(s1[41]), .cout(c1[41]), .a(ps[73]), .b(pc[72]), .c(
        a1s[25]) );
  mul_csa32 sc1_40_ ( .sum(s1[40]), .cout(c1[40]), .a(ps[72]), .b(pc[71]), .c(
        a1s[24]) );
  mul_csa32 sc1_39_ ( .sum(s1[39]), .cout(c1[39]), .a(ps[71]), .b(pc[70]), .c(
        a1s[23]) );
  mul_csa32 sc1_38_ ( .sum(s1[38]), .cout(c1[38]), .a(ps[70]), .b(pc[69]), .c(
        a1s[22]) );
  mul_csa32 sc1_37_ ( .sum(s1[37]), .cout(c1[37]), .a(ps[69]), .b(pc[68]), .c(
        a1s[21]) );
  mul_csa32 sc1_36_ ( .sum(s1[36]), .cout(c1[36]), .a(ps[68]), .b(pc[67]), .c(
        a1s[20]) );
  mul_csa32 sc1_35_ ( .sum(s1[35]), .cout(c1[35]), .a(ps[67]), .b(pc[66]), .c(
        a1s[19]) );
  mul_csa32 sc1_34_ ( .sum(s1[34]), .cout(c1[34]), .a(ps[66]), .b(pc[65]), .c(
        a1s[18]) );
  mul_csa32 sc1_33_ ( .sum(s1[33]), .cout(c1[33]), .a(ps[65]), .b(pc[64]), .c(
        a1s[17]) );
  mul_csa32 sc1_32_ ( .sum(s1[32]), .cout(c1[32]), .a(ps[64]), .b(pc[63]), .c(
        a1s[16]) );
  mul_csa32 sc1_31_ ( .sum(s1[31]), .cout(c1[31]), .a(ps[63]), .b(pc[62]), .c(
        a1s[15]) );
  mul_csa32 sc1_30_ ( .sum(s1[30]), .cout(c1[30]), .a(ps[62]), .b(pc[61]), .c(
        a1s[14]) );
  mul_csa32 sc1_29_ ( .sum(s1[29]), .cout(c1[29]), .a(ps[61]), .b(pc[60]), .c(
        a1s[13]) );
  mul_csa32 sc1_28_ ( .sum(s1[28]), .cout(c1[28]), .a(ps[60]), .b(pc[59]), .c(
        a1s[12]) );
  mul_csa32 sc1_27_ ( .sum(s1[27]), .cout(c1[27]), .a(ps[59]), .b(pc[58]), .c(
        a1s[11]) );
  mul_csa32 sc1_26_ ( .sum(s1[26]), .cout(c1[26]), .a(ps[58]), .b(pc[57]), .c(
        a1s[10]) );
  mul_csa32 sc1_25_ ( .sum(s1[25]), .cout(c1[25]), .a(ps[57]), .b(pc[56]), .c(
        a1s[9]) );
  mul_csa32 sc1_24_ ( .sum(s1[24]), .cout(c1[24]), .a(ps[56]), .b(pc[55]), .c(
        a1s[8]) );
  mul_csa32 sc1_23_ ( .sum(s1[23]), .cout(c1[23]), .a(ps[55]), .b(pc[54]), .c(
        a1s[7]) );
  mul_csa32 sc1_22_ ( .sum(s1[22]), .cout(c1[22]), .a(ps[54]), .b(pc[53]), .c(
        a1s[6]) );
  mul_csa32 sc1_21_ ( .sum(s1[21]), .cout(c1[21]), .a(ps[53]), .b(pc[52]), .c(
        a1s[5]) );
  mul_csa32 sc1_20_ ( .sum(s1[20]), .cout(c1[20]), .a(ps[52]), .b(pc[51]), .c(
        a1s[4]) );
  mul_csa32 sc2_81_ ( .sum(s2[81]), .cout(c2[81]), .a(s1[81]), .b(c1[80]), .c(
        a0c[80]) );
  mul_csa32 sc2_80_ ( .sum(s2[80]), .cout(c2[80]), .a(s1[80]), .b(c1[79]), .c(
        a0c[79]) );
  mul_csa32 sc2_79_ ( .sum(s2[79]), .cout(c2[79]), .a(s1[79]), .b(c1[78]), .c(
        a0c[78]) );
  mul_csa32 sc2_78_ ( .sum(s2[78]), .cout(c2[78]), .a(s1[78]), .b(c1[77]), .c(
        a0c[77]) );
  mul_csa32 sc2_77_ ( .sum(s2[77]), .cout(c2[77]), .a(s1[77]), .b(c1[76]), .c(
        a0c[76]) );
  mul_csa32 sc2_76_ ( .sum(s2[76]), .cout(c2[76]), .a(s1[76]), .b(c1[75]), .c(
        a0c[75]) );
  mul_csa32 sc2_75_ ( .sum(s2[75]), .cout(c2[75]), .a(s1[75]), .b(c1[74]), .c(
        a0c[74]) );
  mul_csa32 sc2_74_ ( .sum(s2[74]), .cout(c2[74]), .a(s1[74]), .b(c1[73]), .c(
        a0c[73]) );
  mul_csa32 sc2_73_ ( .sum(s2[73]), .cout(c2[73]), .a(s1[73]), .b(c1[72]), .c(
        a0c[72]) );
  mul_csa32 sc2_72_ ( .sum(s2[72]), .cout(c2[72]), .a(s1[72]), .b(c1[71]), .c(
        a0c[71]) );
  mul_csa32 sc2_71_ ( .sum(s2[71]), .cout(c2[71]), .a(s1[71]), .b(c1[70]), .c(
        a0c[70]) );
  mul_csa32 sc2_70_ ( .sum(s2[70]), .cout(c2[70]), .a(s1[70]), .b(c1[69]), .c(
        a0c[69]) );
  mul_csa32 sc2_69_ ( .sum(s2[69]), .cout(c2[69]), .a(s1[69]), .b(c1[68]), .c(
        a0c[68]) );
  mul_csa32 sc2_68_ ( .sum(s2[68]), .cout(c2[68]), .a(s1[68]), .b(c1[67]), .c(
        a0c[67]) );
  mul_csa32 acc_19_ ( .sum(psum[19]), .cout(pcout[19]), .a(ain[19]), .b(s3[19]), .c(c3[18]) );
  mul_csa32 acc_18_ ( .sum(psum[18]), .cout(pcout[18]), .a(ain[18]), .b(s3[18]), .c(c3[17]) );
  mul_csa32 acc_17_ ( .sum(psum[17]), .cout(pcout[17]), .a(ain[17]), .b(s3[17]), .c(c3[16]) );
  mul_csa32 acc_16_ ( .sum(psum[16]), .cout(pcout[16]), .a(ain[16]), .b(s3[16]), .c(c3[15]) );
  mul_csa32 acc_15_ ( .sum(psum[15]), .cout(pcout[15]), .a(ain[15]), .b(s3[15]), .c(1'b0) );
  mul_csa32 sc1_0_ ( .sum(s1[0]), .cout(c1[0]), .a(ps[32]), .b(pc[31]), .c(
        a0s[0]) );
  mul_csa32 sc1_67_ ( .sum(s1[67]), .cout(c1[67]), .a(a1s[51]), .b(pc[98]), 
        .c(a1c[50]) );
  mul_ha acc_0_ ( .cout(pcout[0]), .sum(psum[0]), .a(ain[0]), .b(s2[0]) );
  mul_ha sc3_98_ ( .cout(pcout[98]), .sum(psum[98]), .a(bot), .b(a1c[81]) );
  mul_ha sc2_96_ ( .cout(c2[96]), .sum(s2[96]), .a(a1s[80]), .b(a1c[79]) );
  mul_ha sc2_95_ ( .cout(c2[95]), .sum(s2[95]), .a(a1s[79]), .b(a1c[78]) );
  mul_ha sc2_94_ ( .cout(c2[94]), .sum(s2[94]), .a(a1s[78]), .b(a1c[77]) );
  mul_ha sc2_93_ ( .cout(c2[93]), .sum(s2[93]), .a(a1s[77]), .b(a1c[76]) );
  mul_ha sc2_92_ ( .cout(c2[92]), .sum(s2[92]), .a(a1s[76]), .b(a1c[75]) );
  mul_ha sc2_91_ ( .cout(c2[91]), .sum(s2[91]), .a(a1s[75]), .b(a1c[74]) );
  mul_ha sc2_90_ ( .cout(c2[90]), .sum(s2[90]), .a(a1s[74]), .b(a1c[73]) );
  mul_ha sc2_89_ ( .cout(c2[89]), .sum(s2[89]), .a(a1s[73]), .b(a1c[72]) );
  mul_ha sc2_88_ ( .cout(c2[88]), .sum(s2[88]), .a(a1s[72]), .b(a1c[71]) );
  mul_ha sc2_87_ ( .cout(c2[87]), .sum(s2[87]), .a(a1s[71]), .b(a1c[70]) );
  mul_ha sc2_86_ ( .cout(c2[86]), .sum(s2[86]), .a(a1s[70]), .b(a1c[69]) );
  mul_ha sc2_85_ ( .cout(c2[85]), .sum(s2[85]), .a(a1s[69]), .b(a1c[68]) );
  mul_ha sc2_84_ ( .cout(c2[84]), .sum(s2[84]), .a(a1s[68]), .b(a1c[67]) );
  mul_ha sc3_81_ ( .cout(c3[81]), .sum(s3[81]), .a(s2[81]), .b(c2[80]) );
  mul_ha sc3_80_ ( .cout(c3[80]), .sum(s3[80]), .a(s2[80]), .b(c2[79]) );
  mul_ha sc3_79_ ( .cout(c3[79]), .sum(s3[79]), .a(s2[79]), .b(c2[78]) );
  mul_ha sc3_78_ ( .cout(c3[78]), .sum(s3[78]), .a(s2[78]), .b(c2[77]) );
  mul_ha sc3_77_ ( .cout(c3[77]), .sum(s3[77]), .a(s2[77]), .b(c2[76]) );
  mul_ha sc3_76_ ( .cout(c3[76]), .sum(s3[76]), .a(s2[76]), .b(c2[75]) );
  mul_ha sc3_75_ ( .cout(c3[75]), .sum(s3[75]), .a(s2[75]), .b(c2[74]) );
  mul_ha sc3_74_ ( .cout(c3[74]), .sum(s3[74]), .a(s2[74]), .b(c2[73]) );
  mul_ha sc3_73_ ( .cout(c3[73]), .sum(s3[73]), .a(s2[73]), .b(c2[72]) );
  mul_ha sc3_72_ ( .cout(c3[72]), .sum(s3[72]), .a(s2[72]), .b(c2[71]) );
  mul_ha sc3_71_ ( .cout(c3[71]), .sum(s3[71]), .a(s2[71]), .b(c2[70]) );
  mul_ha sc3_70_ ( .cout(c3[70]), .sum(s3[70]), .a(s2[70]), .b(c2[69]) );
  mul_ha sc3_69_ ( .cout(c3[69]), .sum(s3[69]), .a(s2[69]), .b(c2[68]) );
  mul_ha accx2 ( .cout(pcoutx2), .sum(psumx2), .a(ainx2), .b(s1x2) );
  mul_ha sc2_4_ ( .cout(c2[4]), .sum(s2[4]), .a(s1[4]), .b(c1[3]) );
  mul_ha sc2_3_ ( .cout(c2[3]), .sum(s2[3]), .a(s1[3]), .b(c1[2]) );
  mul_ha sc2_2_ ( .cout(c2[2]), .sum(s2[2]), .a(s1[2]), .b(c1[1]) );
  mul_ha sc2_1_ ( .cout(c2[1]), .sum(s2[1]), .a(s1[1]), .b(c1[0]) );
  mul_ha sc2_0_ ( .cout(c2[0]), .sum(s2[0]), .a(s1[0]), .b(c1x2) );
  mul_ha sc1x2 ( .cout(c1x2), .sum(s1x2), .a(ps[31]), .b(pc[30]) );
endmodule


module dp_mux2es_SIZE97 ( dout, in0, in1, sel );
  output [96:0] dout;
  input [96:0] in0;
  input [96:0] in1;
  input sel;
  wire   N0, N1, N2;

  SELECT_OP C107 ( .DATA1(in1), .DATA2(in0), .CONTROL1(N0), .CONTROL2(N1), .Z(
        dout) );
  GTECH_BUF B_0 ( .A(sel), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(sel), .Z(N2) );
endmodule


module dff_SIZE97 ( din, clk, q, se, si, so );
  input [96:0] din;
  output [96:0] q;
  input [96:0] si;
  output [96:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99;
  assign so[96] = q[96];
  assign so[95] = q[95];
  assign so[94] = q[94];
  assign so[93] = q[93];
  assign so[92] = q[92];
  assign so[91] = q[91];
  assign so[90] = q[90];
  assign so[89] = q[89];
  assign so[88] = q[88];
  assign so[87] = q[87];
  assign so[86] = q[86];
  assign so[85] = q[85];
  assign so[84] = q[84];
  assign so[83] = q[83];
  assign so[82] = q[82];
  assign so[81] = q[81];
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(N99), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(N98), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(N97), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(N96), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(N95), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(N94), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(N93), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(N92), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(N91), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(N90), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(N89), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(N88), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(N87), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(N86), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(N85), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C107 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, 
        N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dp_mux2es_SIZE98 ( dout, in0, in1, sel );
  output [97:0] dout;
  input [97:0] in0;
  input [97:0] in1;
  input sel;
  wire   N0, N1, N2;

  SELECT_OP C108 ( .DATA1(in1), .DATA2(in0), .CONTROL1(N0), .CONTROL2(N1), .Z(
        dout) );
  GTECH_BUF B_0 ( .A(sel), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(sel), .Z(N2) );
endmodule


module dff_SIZE98 ( din, clk, q, se, si, so );
  input [97:0] din;
  output [97:0] q;
  input [97:0] si;
  output [97:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100;
  assign so[97] = q[97];
  assign so[96] = q[96];
  assign so[95] = q[95];
  assign so[94] = q[94];
  assign so[93] = q[93];
  assign so[92] = q[92];
  assign so[91] = q[91];
  assign so[90] = q[90];
  assign so[89] = q[89];
  assign so[88] = q[88];
  assign so[87] = q[87];
  assign so[86] = q[86];
  assign so[85] = q[85];
  assign so[84] = q[84];
  assign so[83] = q[83];
  assign so[82] = q[82];
  assign so[81] = q[81];
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[97]  ( .clear(1'b0), .preset(1'b0), .next_state(N100), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(N99), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(N98), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(N97), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(N96), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(N95), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(N94), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(N93), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(N92), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(N91), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(N90), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(N89), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(N88), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(N87), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(N86), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(N85), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C108 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, 
        N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE68 ( din, clk, q, se, si, so );
  input [67:0] din;
  output [67:0] q;
  input [67:0] si;
  output [67:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70;
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C78 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE69 ( din, clk, q, se, si, so );
  input [68:0] din;
  output [68:0] q;
  input [68:0] si;
  output [68:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71;
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C79 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE104 ( din, clk, q, se, si, so );
  input [103:0] din;
  output [103:0] q;
  input [103:0] si;
  output [103:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106;
  assign so[103] = q[103];
  assign so[102] = q[102];
  assign so[101] = q[101];
  assign so[100] = q[100];
  assign so[99] = q[99];
  assign so[98] = q[98];
  assign so[97] = q[97];
  assign so[96] = q[96];
  assign so[95] = q[95];
  assign so[94] = q[94];
  assign so[93] = q[93];
  assign so[92] = q[92];
  assign so[91] = q[91];
  assign so[90] = q[90];
  assign so[89] = q[89];
  assign so[88] = q[88];
  assign so[87] = q[87];
  assign so[86] = q[86];
  assign so[85] = q[85];
  assign so[84] = q[84];
  assign so[83] = q[83];
  assign so[82] = q[82];
  assign so[81] = q[81];
  assign so[80] = q[80];
  assign so[79] = q[79];
  assign so[78] = q[78];
  assign so[77] = q[77];
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[103]  ( .clear(1'b0), .preset(1'b0), .next_state(N106), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[103]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[102]  ( .clear(1'b0), .preset(1'b0), .next_state(N105), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[102]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[101]  ( .clear(1'b0), .preset(1'b0), .next_state(N104), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[101]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[100]  ( .clear(1'b0), .preset(1'b0), .next_state(N103), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[100]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[99]  ( .clear(1'b0), .preset(1'b0), .next_state(N102), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[98]  ( .clear(1'b0), .preset(1'b0), .next_state(N101), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[97]  ( .clear(1'b0), .preset(1'b0), .next_state(N100), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[96]  ( .clear(1'b0), .preset(1'b0), .next_state(N99), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[95]  ( .clear(1'b0), .preset(1'b0), .next_state(N98), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[94]  ( .clear(1'b0), .preset(1'b0), .next_state(N97), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[93]  ( .clear(1'b0), .preset(1'b0), .next_state(N96), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[92]  ( .clear(1'b0), .preset(1'b0), .next_state(N95), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[91]  ( .clear(1'b0), .preset(1'b0), .next_state(N94), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[90]  ( .clear(1'b0), .preset(1'b0), .next_state(N93), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[89]  ( .clear(1'b0), .preset(1'b0), .next_state(N92), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[88]  ( .clear(1'b0), .preset(1'b0), .next_state(N91), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[87]  ( .clear(1'b0), .preset(1'b0), .next_state(N90), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[86]  ( .clear(1'b0), .preset(1'b0), .next_state(N89), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[85]  ( .clear(1'b0), .preset(1'b0), .next_state(N88), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[84]  ( .clear(1'b0), .preset(1'b0), .next_state(N87), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[83]  ( .clear(1'b0), .preset(1'b0), .next_state(N86), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[82]  ( .clear(1'b0), .preset(1'b0), .next_state(N85), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[81]  ( .clear(1'b0), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[80]  ( .clear(1'b0), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[79]  ( .clear(1'b0), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[78]  ( .clear(1'b0), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[77]  ( .clear(1'b0), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C114 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, 
        N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module mul64 ( rs1_l, rs2, valid, areg, accreg, x2, out, rclk, si, so, se, 
        mul_rst_l, mul_step );
  input [63:0] rs1_l;
  input [63:0] rs2;
  input [96:0] areg;
  input [135:129] accreg;
  output [135:0] out;
  input valid, x2, rclk, si, se, mul_rst_l, mul_step;
  output so;
  wire   rst, tm_l, clk_enb0, _0_net_, cyc1, cyc2, cyc3, x2_c1, x2_c2, x2_c3,
         x2_c2c3, clk_enb1, _1_net_, b16, pcoutx2, psumx2, add_co31, add_cin,
         addin_cin, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13,
         N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, add_co96, N66,
         net12994, net12995, net12996, net12997, net12998, net12999, net13000,
         net13001, net13002, net13003, net13004, net13005, net13006, net13007,
         net13008, net13009, net13010, net13011, net13012, net13013, net13014,
         net13015, net13016, net13017, net13018, net13019, net13020, net13021,
         net13022, net13023, net13024, net13025, net13026, net13027, net13028,
         net13029, net13030, net13031, net13032, net13033, net13034, net13035,
         net13036, net13037, net13038, net13039, net13040, net13041, net13042,
         net13043, net13044, net13045, net13046, net13047, net13048, net13049,
         net13050, net13051, net13052, net13053, net13054, net13055, net13056,
         net13057, net13058, net13059, net13060, net13061, net13062, net13063,
         net13064, net13065, net13066, net13067, net13068, net13069, net13070,
         net13071, net13072, net13073, net13074, net13075, net13076, net13077,
         net13078, net13079, net13080, net13081, net13082, net13083, net13084,
         net13085, net13086, net13087, net13088, net13089, net13090, net13091,
         net13092, net13093, net13094, net13095, net13096, net13097, net13098,
         net13099, net13100, net13101, net13102, net13103, net13104, net13105,
         net13106, net13107, net13108, net13109, net13110, net13111, net13112,
         net13113, net13114, net13115, net13116, net13117, net13118, net13119,
         net13120, net13121, net13122, net13123, net13124, net13125, net13126,
         net13127, net13128, net13129, net13130, net13131, net13132, net13133,
         net13134, net13135, net13136, net13137, net13138, net13139, net13140,
         net13141, net13142, net13143, net13144, net13145, net13146, net13147,
         net13148, net13149, net13150, net13151, net13152, net13153, net13154,
         net13155, net13156, net13157, net13158, net13159, net13160, net13161,
         net13162, net13163, net13164, net13165, net13166, net13167, net13168,
         net13169, net13170, net13171, net13172, net13173, net13174, net13175,
         net13176, net13177, net13178, net13179, net13180, net13181, net13182,
         net13183, net13184, net13185, net13186, net13187, net13188, net13189,
         net13190, net13191, net13192, net13193, net13194, net13195, net13196,
         net13197, net13198, net13199, net13200, net13201, net13202, net13203,
         net13204, net13205, net13206, net13207, net13208, net13209, net13210,
         net13211, net13212, net13213, net13214, net13215, net13216, net13217,
         net13218, net13219, net13220, net13221, net13222, net13223, net13224,
         net13225, net13226, net13227, net13228, net13229, net13230, net13231,
         net13232, net13233, net13234, net13235, net13236, net13237, net13238,
         net13239, net13240, net13241, net13242, net13243, net13244, net13245,
         net13246, net13247, net13248, net13249, net13250, net13251, net13252,
         net13253, net13254, net13255, net13256, net13257, net13258, net13259,
         net13260, net13261, net13262, net13263, net13264, net13265, net13266,
         net13267, net13268, net13269, net13270, net13271, net13272, net13273,
         net13274, net13275, net13276, net13277, net13278, net13279, net13280,
         net13281, net13282, net13283, net13284, net13285, net13286, net13287,
         net13288, net13289, net13290, net13291, net13292, net13293, net13294,
         net13295, net13296, net13297, net13298, net13299, net13300, net13301,
         net13302, net13303, net13304, net13305, net13306, net13307, net13308,
         net13309, net13310, net13311, net13312, net13313, net13314, net13315,
         net13316, net13317, net13318, net13319, net13320, net13321, net13322,
         net13323, net13324, net13325, net13326, net13327, net13328, net13329,
         net13330, net13331, net13332, net13333, net13334, net13335, net13336,
         net13337, net13338, net13339, net13340, net13341, net13342, net13343,
         net13344, net13345, net13346, net13347, net13348, net13349, net13350,
         net13351, net13352, net13353, net13354, net13355, net13356, net13357,
         net13358, net13359, net13360, net13361, net13362, net13363, net13364,
         net13365, net13366, net13367, net13368, net13369, net13370, net13371,
         net13372, net13373, net13374, net13375, net13376, net13377, net13378,
         net13379, net13380, net13381, net13382, net13383, net13384, net13385,
         net13386, net13387, net13388, net13389, net13390, net13391, net13392,
         net13393, net13394, net13395, net13396, net13397, net13398, net13399,
         net13400, net13401, net13402, net13403, net13404, net13405, net13406,
         net13407, net13408, net13409, net13410, net13411, net13412, net13413,
         net13414, net13415, net13416, net13417, net13418, net13419, net13420,
         net13421, net13422, net13423, net13424, net13425, net13426, net13427,
         net13428, net13429, net13430, net13431, net13432, net13433, net13434,
         net13435, net13436, net13437, net13438, net13439, net13440, net13441,
         net13442, net13443, net13444, net13445, net13446, net13447, net13448,
         net13449, net13450, net13451, net13452, net13453, net13454, net13455,
         net13456, net13457, net13458, net13459, net13460, net13461, net13462,
         net13463, net13464, net13465, net13466, net13467, net13468, net13469,
         net13470, net13471, net13472, net13473, net13474, net13475, net13476,
         net13477, net13478, net13479, net13480, net13481, net13482, net13483,
         net13484, net13485, net13486, net13487, net13488, net13489, net13490,
         net13491, net13492, net13493, net13494, net13495, net13496, net13497,
         net13498, net13499, net13500, net13501, net13502, net13503, net13504,
         net13505, net13506, net13507, net13508, net13509, net13510, net13511,
         net13512, net13513, net13514, net13515, net13516, net13517, net13518,
         net13519, net13520, net13521, net13522, net13523, net13524, net13525,
         net13526, net13527, net13528, net13529, net13530, net13531, net13532,
         net13533, net13534, net13535, net13536, net13537, net13538, net13539,
         net13540, net13541, net13542, net13543, net13544, net13545, net13546,
         net13547, net13548, net13549, net13550, net13551, net13552, net13553,
         net13554, net13555, net13556, net13557, net13558, net13559, net13560,
         net13561, net13562, net13563, net13564, net13565, net13566, net13567,
         net13568, net13569, net13570, net13571, net13572, net13573, net13574,
         net13575, net13576, net13577, net13578, net13579, net13580, net13581,
         net13582, net13583, net13584, net13585, net13586, net13587, net13588,
         net13589, net13590, net13591, net13592, net13593, net13594, net13595,
         net13596, net13597, net13598, net13599, net13600, net13601, net13602,
         net13603, net13604, net13605, net13606, net13607, net13608, net13609,
         net13610, net13611, net13612, net13613, net13614, net13615, net13616,
         net13617, net13618, net13619, net13620, net13621, net13622, net13623,
         net13624, net13625, net13626, net13627, net13628, net13629, net13630,
         net13631, net13632, net13633, net13634, net13635, net13636, net13637,
         net13638, net13639, net13640, net13641, net13642, net13643, net13644,
         net13645, net13646, net13647, net13648, net13649, net13650, net13651,
         net13652, net13653, net13654, net13655, net13656, net13657, net13658,
         net13659, net13660, net13661, net13662, net13663, net13664, net13665,
         net13666, net13667, net13668, net13669, net13670, net13671, net13672,
         net13673, net13674, net13675, net13676, net13677, net13678, net13679,
         net13680, net13681, net13682, net13683, net13684, net13685, net13686,
         net13687, net13688, net13689, net13690, net13691, net13692, net13693,
         net13694, net13695, net13696, net13697, net13698, net13699, net13700,
         net13701, net13702, net13703, net13704, net13705, net13706, net13707,
         net13708, net13709, net13710, net13711, net13712, net13713, net13714,
         net13715, net13716, net13717, net13718, net13719, net13720, net13721,
         net13722, net13723, net13724, net13725, net13726, net13727, net13728,
         net13729, net13730, net13731, net13732, net13733, net13734, net13735,
         net13736, net13737, net13738, net13739, net13740, net13741, net13742,
         net13743, net13744, net13745, net13746, net13747, net13748, net13749,
         net13750, net13751, net13752, net13753, net13754, net13755, net13756,
         net13757, net13758, net13759, net13760, net13761, net13762, net13763,
         net13764, net13765, net13766, net13767, net13768, net13769, net13770,
         net13771, net13772, net13773, net13774, net13775, net13776, net13777,
         net13778, net13779, net13780, net13781, net13782, net13783, net13784,
         net13785, net13786, net13787, net13788, net13789, net13790, net13791,
         net13792, net13793, net13794, net13795, net13796, net13797, net13798,
         net13799, net13800, net13801, net13802, net13803, net13804, net13805,
         net13806, net13807, net13808, net13809, net13810, net13811, net13812,
         net13813, net13814, net13815, net13816, net13817, net13818, net13819,
         net13820, net13821, net13822, net13823, net13824, net13825, net13826,
         net13827, net13828, net13829, net13830, net13831, net13832, net13833,
         net13834, net13835, net13836, net13837, net13838, net13839, net13840,
         net13841, net13842, net13843, net13844, net13845, net13846, net13847,
         net13848, net13849, net13850, net13851, net13852, net13853, net13854;
  wire   [63:0] op1_l;
  wire   [63:0] op1;
  wire   [2:0] b0;
  wire   [2:0] b1;
  wire   [2:0] b2;
  wire   [2:0] b3;
  wire   [2:0] b4;
  wire   [2:0] b5;
  wire   [2:0] b6;
  wire   [2:0] b7;
  wire   [2:0] b8;
  wire   [2:0] b9;
  wire   [2:0] b10;
  wire   [2:0] b11;
  wire   [2:0] b12;
  wire   [2:0] b13;
  wire   [2:0] b14;
  wire   [2:0] b15;
  wire   [81:4] a0cout;
  wire   [81:0] a0sum;
  wire   [81:4] a0c;
  wire   [81:0] a0s;
  wire   [81:4] a1cout;
  wire   [81:0] a1sum;
  wire   [81:4] a1c;
  wire   [81:0] a1s;
  wire   [98:0] pcout;
  wire   [98:0] psum;
  wire   [98:30] pc;
  wire   [98:31] ps;
  wire   [96:0] ary2_cout;
  wire   [96:0] addin_cout;
  wire   [97:0] ary2_sum;
  wire   [97:0] addin_sum;
  wire   [98:31] psum_in;
  wire   [98:30] pcout_in;
  wire   [103:0] addout;

  clken_buf ckbuf_0 ( .clk(clk_enb0), .rclk(rclk), .enb_l(_0_net_), .tmb_l(
        tm_l) );
  dffr_SIZE1 cyc1_dff ( .din(valid), .clk(clk_enb0), .rst(rst), .q(cyc1), .se(
        se), .si(net13854) );
  dffr_SIZE1 cyc2_dff ( .din(cyc1), .clk(clk_enb0), .rst(rst), .q(cyc2), .se(
        se), .si(net13853) );
  dffr_SIZE1 cyc3_dff ( .din(cyc2), .clk(clk_enb0), .rst(rst), .q(cyc3), .se(
        se), .si(net13852) );
  dffr_SIZE1 x2c1_dff ( .din(x2), .clk(clk_enb0), .rst(rst), .q(x2_c1), .se(se), .si(net13851) );
  dffr_SIZE1 x2c2_dff ( .din(x2_c1), .clk(clk_enb0), .rst(rst), .q(x2_c2), 
        .se(se), .si(net13850) );
  dffr_SIZE1 x2c3_dff ( .din(x2_c2), .clk(clk_enb0), .rst(rst), .q(x2_c3), 
        .se(se), .si(net13849) );
  clken_buf ckbuf_1 ( .clk(clk_enb1), .rclk(rclk), .enb_l(_1_net_), .tmb_l(
        tm_l) );
  dff_SIZE64 ffrs1 ( .din(rs1_l), .clk(clk_enb1), .q(op1_l), .se(se), .si({
        net13785, net13786, net13787, net13788, net13789, net13790, net13791, 
        net13792, net13793, net13794, net13795, net13796, net13797, net13798, 
        net13799, net13800, net13801, net13802, net13803, net13804, net13805, 
        net13806, net13807, net13808, net13809, net13810, net13811, net13812, 
        net13813, net13814, net13815, net13816, net13817, net13818, net13819, 
        net13820, net13821, net13822, net13823, net13824, net13825, net13826, 
        net13827, net13828, net13829, net13830, net13831, net13832, net13833, 
        net13834, net13835, net13836, net13837, net13838, net13839, net13840, 
        net13841, net13842, net13843, net13844, net13845, net13846, net13847, 
        net13848}) );
  mul_booth booth ( .head(valid), .b_in(rs2), .b0(b0), .b1(b1), .b2(b2), .b3(
        b3), .b4(b4), .b5(b5), .b6(b6), .b7(b7), .b8(b8), .b9(b9), .b10(b10), 
        .b11(b11), .b12(b12), .b13(b13), .b14(b14), .b15(b15), .b16(b16), 
        .clk(rclk), .se(se), .si(net13784), .mul_step(mul_step), .tm_l(tm_l)
         );
  mul_array1 ary1_a0 ( .cout(a0cout), .sum(a0sum), .a(op1), .b0(b0), .b1(b1), 
        .b2(b2), .b3(b3), .b4(b4), .b5(b5), .b6(b6), .b7(b7), .b8({1'b0, 1'b0, 
        1'b0}), .bot(1'b0), .head(cyc1) );
  dff_SIZE78 a0cot_dff ( .din(a0cout), .clk(clk_enb0), .q(a0c), .se(se), .si({
        net13706, net13707, net13708, net13709, net13710, net13711, net13712, 
        net13713, net13714, net13715, net13716, net13717, net13718, net13719, 
        net13720, net13721, net13722, net13723, net13724, net13725, net13726, 
        net13727, net13728, net13729, net13730, net13731, net13732, net13733, 
        net13734, net13735, net13736, net13737, net13738, net13739, net13740, 
        net13741, net13742, net13743, net13744, net13745, net13746, net13747, 
        net13748, net13749, net13750, net13751, net13752, net13753, net13754, 
        net13755, net13756, net13757, net13758, net13759, net13760, net13761, 
        net13762, net13763, net13764, net13765, net13766, net13767, net13768, 
        net13769, net13770, net13771, net13772, net13773, net13774, net13775, 
        net13776, net13777, net13778, net13779, net13780, net13781, net13782, 
        net13783}) );
  dff_SIZE82 a0sum_dff ( .din(a0sum), .clk(clk_enb0), .q(a0s), .se(se), .si({
        net13624, net13625, net13626, net13627, net13628, net13629, net13630, 
        net13631, net13632, net13633, net13634, net13635, net13636, net13637, 
        net13638, net13639, net13640, net13641, net13642, net13643, net13644, 
        net13645, net13646, net13647, net13648, net13649, net13650, net13651, 
        net13652, net13653, net13654, net13655, net13656, net13657, net13658, 
        net13659, net13660, net13661, net13662, net13663, net13664, net13665, 
        net13666, net13667, net13668, net13669, net13670, net13671, net13672, 
        net13673, net13674, net13675, net13676, net13677, net13678, net13679, 
        net13680, net13681, net13682, net13683, net13684, net13685, net13686, 
        net13687, net13688, net13689, net13690, net13691, net13692, net13693, 
        net13694, net13695, net13696, net13697, net13698, net13699, net13700, 
        net13701, net13702, net13703, net13704, net13705}) );
  mul_array1 ary1_a1 ( .cout(a1cout), .sum(a1sum), .a(op1), .b0(b8), .b1(b9), 
        .b2(b10), .b3(b11), .b4(b12), .b5(b13), .b6(b14), .b7(b15), .b8({1'b0, 
        b16, 1'b0}), .bot(cyc2), .head(1'b0) );
  dff_SIZE78 a1cot_dff ( .din(a1cout), .clk(clk_enb0), .q(a1c), .se(se), .si({
        net13546, net13547, net13548, net13549, net13550, net13551, net13552, 
        net13553, net13554, net13555, net13556, net13557, net13558, net13559, 
        net13560, net13561, net13562, net13563, net13564, net13565, net13566, 
        net13567, net13568, net13569, net13570, net13571, net13572, net13573, 
        net13574, net13575, net13576, net13577, net13578, net13579, net13580, 
        net13581, net13582, net13583, net13584, net13585, net13586, net13587, 
        net13588, net13589, net13590, net13591, net13592, net13593, net13594, 
        net13595, net13596, net13597, net13598, net13599, net13600, net13601, 
        net13602, net13603, net13604, net13605, net13606, net13607, net13608, 
        net13609, net13610, net13611, net13612, net13613, net13614, net13615, 
        net13616, net13617, net13618, net13619, net13620, net13621, net13622, 
        net13623}) );
  dff_SIZE82 a1sum_dff ( .din(a1sum), .clk(clk_enb0), .q(a1s), .se(se), .si({
        net13464, net13465, net13466, net13467, net13468, net13469, net13470, 
        net13471, net13472, net13473, net13474, net13475, net13476, net13477, 
        net13478, net13479, net13480, net13481, net13482, net13483, net13484, 
        net13485, net13486, net13487, net13488, net13489, net13490, net13491, 
        net13492, net13493, net13494, net13495, net13496, net13497, net13498, 
        net13499, net13500, net13501, net13502, net13503, net13504, net13505, 
        net13506, net13507, net13508, net13509, net13510, net13511, net13512, 
        net13513, net13514, net13515, net13516, net13517, net13518, net13519, 
        net13520, net13521, net13522, net13523, net13524, net13525, net13526, 
        net13527, net13528, net13529, net13530, net13531, net13532, net13533, 
        net13534, net13535, net13536, net13537, net13538, net13539, net13540, 
        net13541, net13542, net13543, net13544, net13545}) );
  mul_array2 array2 ( .pcout(pcout), .pcoutx2(pcoutx2), .psum(psum), .psumx2(
        psumx2), .a0c(a0c), .a0s(a0s), .a1c(a1c), .a1s(a1s), .areg(areg), 
        .bot(cyc3), .pc(pc), .ps(ps), .x2(x2_c2c3) );
  dp_mux2es_SIZE97 ary2_cmux ( .dout(ary2_cout), .in0(pcout[96:0]), .in1({
        pcout[95:0], pcoutx2}), .sel(x2_c2c3) );
  dff_SIZE97 a2cot_dff ( .din(ary2_cout), .clk(clk_enb0), .q(addin_cout), .se(
        se), .si({net13367, net13368, net13369, net13370, net13371, net13372, 
        net13373, net13374, net13375, net13376, net13377, net13378, net13379, 
        net13380, net13381, net13382, net13383, net13384, net13385, net13386, 
        net13387, net13388, net13389, net13390, net13391, net13392, net13393, 
        net13394, net13395, net13396, net13397, net13398, net13399, net13400, 
        net13401, net13402, net13403, net13404, net13405, net13406, net13407, 
        net13408, net13409, net13410, net13411, net13412, net13413, net13414, 
        net13415, net13416, net13417, net13418, net13419, net13420, net13421, 
        net13422, net13423, net13424, net13425, net13426, net13427, net13428, 
        net13429, net13430, net13431, net13432, net13433, net13434, net13435, 
        net13436, net13437, net13438, net13439, net13440, net13441, net13442, 
        net13443, net13444, net13445, net13446, net13447, net13448, net13449, 
        net13450, net13451, net13452, net13453, net13454, net13455, net13456, 
        net13457, net13458, net13459, net13460, net13461, net13462, net13463})
         );
  dp_mux2es_SIZE98 ary2_smux ( .dout(ary2_sum), .in0(psum[97:0]), .in1({
        psum[96:0], psumx2}), .sel(x2_c2c3) );
  dff_SIZE98 a2sum_dff ( .din(ary2_sum), .clk(clk_enb0), .q(addin_sum), .se(se), .si({net13269, net13270, net13271, net13272, net13273, net13274, net13275, 
        net13276, net13277, net13278, net13279, net13280, net13281, net13282, 
        net13283, net13284, net13285, net13286, net13287, net13288, net13289, 
        net13290, net13291, net13292, net13293, net13294, net13295, net13296, 
        net13297, net13298, net13299, net13300, net13301, net13302, net13303, 
        net13304, net13305, net13306, net13307, net13308, net13309, net13310, 
        net13311, net13312, net13313, net13314, net13315, net13316, net13317, 
        net13318, net13319, net13320, net13321, net13322, net13323, net13324, 
        net13325, net13326, net13327, net13328, net13329, net13330, net13331, 
        net13332, net13333, net13334, net13335, net13336, net13337, net13338, 
        net13339, net13340, net13341, net13342, net13343, net13344, net13345, 
        net13346, net13347, net13348, net13349, net13350, net13351, net13352, 
        net13353, net13354, net13355, net13356, net13357, net13358, net13359, 
        net13360, net13361, net13362, net13363, net13364, net13365, net13366})
         );
  dff_SIZE68 psum_dff ( .din(psum_in), .clk(clk_enb0), .q(ps), .se(se), .si({
        net13201, net13202, net13203, net13204, net13205, net13206, net13207, 
        net13208, net13209, net13210, net13211, net13212, net13213, net13214, 
        net13215, net13216, net13217, net13218, net13219, net13220, net13221, 
        net13222, net13223, net13224, net13225, net13226, net13227, net13228, 
        net13229, net13230, net13231, net13232, net13233, net13234, net13235, 
        net13236, net13237, net13238, net13239, net13240, net13241, net13242, 
        net13243, net13244, net13245, net13246, net13247, net13248, net13249, 
        net13250, net13251, net13252, net13253, net13254, net13255, net13256, 
        net13257, net13258, net13259, net13260, net13261, net13262, net13263, 
        net13264, net13265, net13266, net13267, net13268}) );
  dff_SIZE69 pcout_dff ( .din(pcout_in), .clk(clk_enb0), .q(pc), .se(se), .si(
        {net13132, net13133, net13134, net13135, net13136, net13137, net13138, 
        net13139, net13140, net13141, net13142, net13143, net13144, net13145, 
        net13146, net13147, net13148, net13149, net13150, net13151, net13152, 
        net13153, net13154, net13155, net13156, net13157, net13158, net13159, 
        net13160, net13161, net13162, net13163, net13164, net13165, net13166, 
        net13167, net13168, net13169, net13170, net13171, net13172, net13173, 
        net13174, net13175, net13176, net13177, net13178, net13179, net13180, 
        net13181, net13182, net13183, net13184, net13185, net13186, net13187, 
        net13188, net13189, net13190, net13191, net13192, net13193, net13194, 
        net13195, net13196, net13197, net13198, net13199, net13200}) );
  dff_SIZE1 co31_dff ( .din(add_cin), .clk(clk_enb0), .q(addin_cin), .se(se), 
        .si(net13131) );
  dff_SIZE104 out_dff ( .din(addout), .clk(clk_enb0), .q(out[135:32]), .se(se), 
        .si({net13027, net13028, net13029, net13030, net13031, net13032, 
        net13033, net13034, net13035, net13036, net13037, net13038, net13039, 
        net13040, net13041, net13042, net13043, net13044, net13045, net13046, 
        net13047, net13048, net13049, net13050, net13051, net13052, net13053, 
        net13054, net13055, net13056, net13057, net13058, net13059, net13060, 
        net13061, net13062, net13063, net13064, net13065, net13066, net13067, 
        net13068, net13069, net13070, net13071, net13072, net13073, net13074, 
        net13075, net13076, net13077, net13078, net13079, net13080, net13081, 
        net13082, net13083, net13084, net13085, net13086, net13087, net13088, 
        net13089, net13090, net13091, net13092, net13093, net13094, net13095, 
        net13096, net13097, net13098, net13099, net13100, net13101, net13102, 
        net13103, net13104, net13105, net13106, net13107, net13108, net13109, 
        net13110, net13111, net13112, net13113, net13114, net13115, net13116, 
        net13117, net13118, net13119, net13120, net13121, net13122, net13123, 
        net13124, net13125, net13126, net13127, net13128, net13129, net13130})
         );
  dff_SIZE32 pip_dff ( .din(out[63:32]), .clk(clk_enb0), .q(out[31:0]), .se(se), .si({net12995, net12996, net12997, net12998, net12999, net13000, net13001, 
        net13002, net13003, net13004, net13005, net13006, net13007, net13008, 
        net13009, net13010, net13011, net13012, net13013, net13014, net13015, 
        net13016, net13017, net13018, net13019, net13020, net13021, net13022, 
        net13023, net13024, net13025, net13026}) );
  ADD_UNS_OP add_293 ( .A(addin_sum[97:32]), .B(addin_cout[96:31]), .Z({N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, 
        N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, 
        N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, 
        N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  ADD_UNS_OP add_289 ( .A(addin_sum[31:0]), .B({addin_cout[30:0], addin_cin}), 
        .Z({add_co31, addout[31:0]}) );
  ADD_UNS_OP add_293_2 ( .A({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), .B(
        add_co31), .Z({add_co96, addout[96:32]}) );
  ADD_UNS_OP add_297 ( .A(accreg), .B(add_co96), .Z(addout[103:97]) );
  GTECH_NOT I_0 ( .A(mul_rst_l), .Z(rst) );
  GTECH_NOT I_1 ( .A(se), .Z(tm_l) );
  GTECH_NOT I_2 ( .A(mul_step), .Z(_0_net_) );
  GTECH_OR2 C217 ( .A(x2_c2), .B(x2_c3), .Z(x2_c2c3) );
  GTECH_NOT I_3 ( .A(N66), .Z(_1_net_) );
  GTECH_AND2 C219 ( .A(valid), .B(mul_step), .Z(N66) );
  GTECH_NOT I_4 ( .A(op1_l[63]), .Z(op1[63]) );
  GTECH_NOT I_5 ( .A(op1_l[62]), .Z(op1[62]) );
  GTECH_NOT I_6 ( .A(op1_l[61]), .Z(op1[61]) );
  GTECH_NOT I_7 ( .A(op1_l[60]), .Z(op1[60]) );
  GTECH_NOT I_8 ( .A(op1_l[59]), .Z(op1[59]) );
  GTECH_NOT I_9 ( .A(op1_l[58]), .Z(op1[58]) );
  GTECH_NOT I_10 ( .A(op1_l[57]), .Z(op1[57]) );
  GTECH_NOT I_11 ( .A(op1_l[56]), .Z(op1[56]) );
  GTECH_NOT I_12 ( .A(op1_l[55]), .Z(op1[55]) );
  GTECH_NOT I_13 ( .A(op1_l[54]), .Z(op1[54]) );
  GTECH_NOT I_14 ( .A(op1_l[53]), .Z(op1[53]) );
  GTECH_NOT I_15 ( .A(op1_l[52]), .Z(op1[52]) );
  GTECH_NOT I_16 ( .A(op1_l[51]), .Z(op1[51]) );
  GTECH_NOT I_17 ( .A(op1_l[50]), .Z(op1[50]) );
  GTECH_NOT I_18 ( .A(op1_l[49]), .Z(op1[49]) );
  GTECH_NOT I_19 ( .A(op1_l[48]), .Z(op1[48]) );
  GTECH_NOT I_20 ( .A(op1_l[47]), .Z(op1[47]) );
  GTECH_NOT I_21 ( .A(op1_l[46]), .Z(op1[46]) );
  GTECH_NOT I_22 ( .A(op1_l[45]), .Z(op1[45]) );
  GTECH_NOT I_23 ( .A(op1_l[44]), .Z(op1[44]) );
  GTECH_NOT I_24 ( .A(op1_l[43]), .Z(op1[43]) );
  GTECH_NOT I_25 ( .A(op1_l[42]), .Z(op1[42]) );
  GTECH_NOT I_26 ( .A(op1_l[41]), .Z(op1[41]) );
  GTECH_NOT I_27 ( .A(op1_l[40]), .Z(op1[40]) );
  GTECH_NOT I_28 ( .A(op1_l[39]), .Z(op1[39]) );
  GTECH_NOT I_29 ( .A(op1_l[38]), .Z(op1[38]) );
  GTECH_NOT I_30 ( .A(op1_l[37]), .Z(op1[37]) );
  GTECH_NOT I_31 ( .A(op1_l[36]), .Z(op1[36]) );
  GTECH_NOT I_32 ( .A(op1_l[35]), .Z(op1[35]) );
  GTECH_NOT I_33 ( .A(op1_l[34]), .Z(op1[34]) );
  GTECH_NOT I_34 ( .A(op1_l[33]), .Z(op1[33]) );
  GTECH_NOT I_35 ( .A(op1_l[32]), .Z(op1[32]) );
  GTECH_NOT I_36 ( .A(op1_l[31]), .Z(op1[31]) );
  GTECH_NOT I_37 ( .A(op1_l[30]), .Z(op1[30]) );
  GTECH_NOT I_38 ( .A(op1_l[29]), .Z(op1[29]) );
  GTECH_NOT I_39 ( .A(op1_l[28]), .Z(op1[28]) );
  GTECH_NOT I_40 ( .A(op1_l[27]), .Z(op1[27]) );
  GTECH_NOT I_41 ( .A(op1_l[26]), .Z(op1[26]) );
  GTECH_NOT I_42 ( .A(op1_l[25]), .Z(op1[25]) );
  GTECH_NOT I_43 ( .A(op1_l[24]), .Z(op1[24]) );
  GTECH_NOT I_44 ( .A(op1_l[23]), .Z(op1[23]) );
  GTECH_NOT I_45 ( .A(op1_l[22]), .Z(op1[22]) );
  GTECH_NOT I_46 ( .A(op1_l[21]), .Z(op1[21]) );
  GTECH_NOT I_47 ( .A(op1_l[20]), .Z(op1[20]) );
  GTECH_NOT I_48 ( .A(op1_l[19]), .Z(op1[19]) );
  GTECH_NOT I_49 ( .A(op1_l[18]), .Z(op1[18]) );
  GTECH_NOT I_50 ( .A(op1_l[17]), .Z(op1[17]) );
  GTECH_NOT I_51 ( .A(op1_l[16]), .Z(op1[16]) );
  GTECH_NOT I_52 ( .A(op1_l[15]), .Z(op1[15]) );
  GTECH_NOT I_53 ( .A(op1_l[14]), .Z(op1[14]) );
  GTECH_NOT I_54 ( .A(op1_l[13]), .Z(op1[13]) );
  GTECH_NOT I_55 ( .A(op1_l[12]), .Z(op1[12]) );
  GTECH_NOT I_56 ( .A(op1_l[11]), .Z(op1[11]) );
  GTECH_NOT I_57 ( .A(op1_l[10]), .Z(op1[10]) );
  GTECH_NOT I_58 ( .A(op1_l[9]), .Z(op1[9]) );
  GTECH_NOT I_59 ( .A(op1_l[8]), .Z(op1[8]) );
  GTECH_NOT I_60 ( .A(op1_l[7]), .Z(op1[7]) );
  GTECH_NOT I_61 ( .A(op1_l[6]), .Z(op1[6]) );
  GTECH_NOT I_62 ( .A(op1_l[5]), .Z(op1[5]) );
  GTECH_NOT I_63 ( .A(op1_l[4]), .Z(op1[4]) );
  GTECH_NOT I_64 ( .A(op1_l[3]), .Z(op1[3]) );
  GTECH_NOT I_65 ( .A(op1_l[2]), .Z(op1[2]) );
  GTECH_NOT I_66 ( .A(op1_l[1]), .Z(op1[1]) );
  GTECH_NOT I_67 ( .A(op1_l[0]), .Z(op1[0]) );
  GTECH_AND2 C284 ( .A(psum[98]), .B(cyc2), .Z(psum_in[98]) );
  GTECH_AND2 C285 ( .A(psum[97]), .B(cyc2), .Z(psum_in[97]) );
  GTECH_AND2 C286 ( .A(psum[96]), .B(cyc2), .Z(psum_in[96]) );
  GTECH_AND2 C287 ( .A(psum[95]), .B(cyc2), .Z(psum_in[95]) );
  GTECH_AND2 C288 ( .A(psum[94]), .B(cyc2), .Z(psum_in[94]) );
  GTECH_AND2 C289 ( .A(psum[93]), .B(cyc2), .Z(psum_in[93]) );
  GTECH_AND2 C290 ( .A(psum[92]), .B(cyc2), .Z(psum_in[92]) );
  GTECH_AND2 C291 ( .A(psum[91]), .B(cyc2), .Z(psum_in[91]) );
  GTECH_AND2 C292 ( .A(psum[90]), .B(cyc2), .Z(psum_in[90]) );
  GTECH_AND2 C293 ( .A(psum[89]), .B(cyc2), .Z(psum_in[89]) );
  GTECH_AND2 C294 ( .A(psum[88]), .B(cyc2), .Z(psum_in[88]) );
  GTECH_AND2 C295 ( .A(psum[87]), .B(cyc2), .Z(psum_in[87]) );
  GTECH_AND2 C296 ( .A(psum[86]), .B(cyc2), .Z(psum_in[86]) );
  GTECH_AND2 C297 ( .A(psum[85]), .B(cyc2), .Z(psum_in[85]) );
  GTECH_AND2 C298 ( .A(psum[84]), .B(cyc2), .Z(psum_in[84]) );
  GTECH_AND2 C299 ( .A(psum[83]), .B(cyc2), .Z(psum_in[83]) );
  GTECH_AND2 C300 ( .A(psum[82]), .B(cyc2), .Z(psum_in[82]) );
  GTECH_AND2 C301 ( .A(psum[81]), .B(cyc2), .Z(psum_in[81]) );
  GTECH_AND2 C302 ( .A(psum[80]), .B(cyc2), .Z(psum_in[80]) );
  GTECH_AND2 C303 ( .A(psum[79]), .B(cyc2), .Z(psum_in[79]) );
  GTECH_AND2 C304 ( .A(psum[78]), .B(cyc2), .Z(psum_in[78]) );
  GTECH_AND2 C305 ( .A(psum[77]), .B(cyc2), .Z(psum_in[77]) );
  GTECH_AND2 C306 ( .A(psum[76]), .B(cyc2), .Z(psum_in[76]) );
  GTECH_AND2 C307 ( .A(psum[75]), .B(cyc2), .Z(psum_in[75]) );
  GTECH_AND2 C308 ( .A(psum[74]), .B(cyc2), .Z(psum_in[74]) );
  GTECH_AND2 C309 ( .A(psum[73]), .B(cyc2), .Z(psum_in[73]) );
  GTECH_AND2 C310 ( .A(psum[72]), .B(cyc2), .Z(psum_in[72]) );
  GTECH_AND2 C311 ( .A(psum[71]), .B(cyc2), .Z(psum_in[71]) );
  GTECH_AND2 C312 ( .A(psum[70]), .B(cyc2), .Z(psum_in[70]) );
  GTECH_AND2 C313 ( .A(psum[69]), .B(cyc2), .Z(psum_in[69]) );
  GTECH_AND2 C314 ( .A(psum[68]), .B(cyc2), .Z(psum_in[68]) );
  GTECH_AND2 C315 ( .A(psum[67]), .B(cyc2), .Z(psum_in[67]) );
  GTECH_AND2 C316 ( .A(psum[66]), .B(cyc2), .Z(psum_in[66]) );
  GTECH_AND2 C317 ( .A(psum[65]), .B(cyc2), .Z(psum_in[65]) );
  GTECH_AND2 C318 ( .A(psum[64]), .B(cyc2), .Z(psum_in[64]) );
  GTECH_AND2 C319 ( .A(psum[63]), .B(cyc2), .Z(psum_in[63]) );
  GTECH_AND2 C320 ( .A(psum[62]), .B(cyc2), .Z(psum_in[62]) );
  GTECH_AND2 C321 ( .A(psum[61]), .B(cyc2), .Z(psum_in[61]) );
  GTECH_AND2 C322 ( .A(psum[60]), .B(cyc2), .Z(psum_in[60]) );
  GTECH_AND2 C323 ( .A(psum[59]), .B(cyc2), .Z(psum_in[59]) );
  GTECH_AND2 C324 ( .A(psum[58]), .B(cyc2), .Z(psum_in[58]) );
  GTECH_AND2 C325 ( .A(psum[57]), .B(cyc2), .Z(psum_in[57]) );
  GTECH_AND2 C326 ( .A(psum[56]), .B(cyc2), .Z(psum_in[56]) );
  GTECH_AND2 C327 ( .A(psum[55]), .B(cyc2), .Z(psum_in[55]) );
  GTECH_AND2 C328 ( .A(psum[54]), .B(cyc2), .Z(psum_in[54]) );
  GTECH_AND2 C329 ( .A(psum[53]), .B(cyc2), .Z(psum_in[53]) );
  GTECH_AND2 C330 ( .A(psum[52]), .B(cyc2), .Z(psum_in[52]) );
  GTECH_AND2 C331 ( .A(psum[51]), .B(cyc2), .Z(psum_in[51]) );
  GTECH_AND2 C332 ( .A(psum[50]), .B(cyc2), .Z(psum_in[50]) );
  GTECH_AND2 C333 ( .A(psum[49]), .B(cyc2), .Z(psum_in[49]) );
  GTECH_AND2 C334 ( .A(psum[48]), .B(cyc2), .Z(psum_in[48]) );
  GTECH_AND2 C335 ( .A(psum[47]), .B(cyc2), .Z(psum_in[47]) );
  GTECH_AND2 C336 ( .A(psum[46]), .B(cyc2), .Z(psum_in[46]) );
  GTECH_AND2 C337 ( .A(psum[45]), .B(cyc2), .Z(psum_in[45]) );
  GTECH_AND2 C338 ( .A(psum[44]), .B(cyc2), .Z(psum_in[44]) );
  GTECH_AND2 C339 ( .A(psum[43]), .B(cyc2), .Z(psum_in[43]) );
  GTECH_AND2 C340 ( .A(psum[42]), .B(cyc2), .Z(psum_in[42]) );
  GTECH_AND2 C341 ( .A(psum[41]), .B(cyc2), .Z(psum_in[41]) );
  GTECH_AND2 C342 ( .A(psum[40]), .B(cyc2), .Z(psum_in[40]) );
  GTECH_AND2 C343 ( .A(psum[39]), .B(cyc2), .Z(psum_in[39]) );
  GTECH_AND2 C344 ( .A(psum[38]), .B(cyc2), .Z(psum_in[38]) );
  GTECH_AND2 C345 ( .A(psum[37]), .B(cyc2), .Z(psum_in[37]) );
  GTECH_AND2 C346 ( .A(psum[36]), .B(cyc2), .Z(psum_in[36]) );
  GTECH_AND2 C347 ( .A(psum[35]), .B(cyc2), .Z(psum_in[35]) );
  GTECH_AND2 C348 ( .A(psum[34]), .B(cyc2), .Z(psum_in[34]) );
  GTECH_AND2 C349 ( .A(psum[33]), .B(cyc2), .Z(psum_in[33]) );
  GTECH_AND2 C350 ( .A(psum[32]), .B(cyc2), .Z(psum_in[32]) );
  GTECH_AND2 C351 ( .A(psum[31]), .B(x2_c2), .Z(psum_in[31]) );
  GTECH_AND2 C352 ( .A(pcout[98]), .B(cyc2), .Z(pcout_in[98]) );
  GTECH_AND2 C353 ( .A(pcout[97]), .B(cyc2), .Z(pcout_in[97]) );
  GTECH_AND2 C354 ( .A(pcout[96]), .B(cyc2), .Z(pcout_in[96]) );
  GTECH_AND2 C355 ( .A(pcout[95]), .B(cyc2), .Z(pcout_in[95]) );
  GTECH_AND2 C356 ( .A(pcout[94]), .B(cyc2), .Z(pcout_in[94]) );
  GTECH_AND2 C357 ( .A(pcout[93]), .B(cyc2), .Z(pcout_in[93]) );
  GTECH_AND2 C358 ( .A(pcout[92]), .B(cyc2), .Z(pcout_in[92]) );
  GTECH_AND2 C359 ( .A(pcout[91]), .B(cyc2), .Z(pcout_in[91]) );
  GTECH_AND2 C360 ( .A(pcout[90]), .B(cyc2), .Z(pcout_in[90]) );
  GTECH_AND2 C361 ( .A(pcout[89]), .B(cyc2), .Z(pcout_in[89]) );
  GTECH_AND2 C362 ( .A(pcout[88]), .B(cyc2), .Z(pcout_in[88]) );
  GTECH_AND2 C363 ( .A(pcout[87]), .B(cyc2), .Z(pcout_in[87]) );
  GTECH_AND2 C364 ( .A(pcout[86]), .B(cyc2), .Z(pcout_in[86]) );
  GTECH_AND2 C365 ( .A(pcout[85]), .B(cyc2), .Z(pcout_in[85]) );
  GTECH_AND2 C366 ( .A(pcout[84]), .B(cyc2), .Z(pcout_in[84]) );
  GTECH_AND2 C367 ( .A(pcout[83]), .B(cyc2), .Z(pcout_in[83]) );
  GTECH_AND2 C368 ( .A(pcout[82]), .B(cyc2), .Z(pcout_in[82]) );
  GTECH_AND2 C369 ( .A(pcout[81]), .B(cyc2), .Z(pcout_in[81]) );
  GTECH_AND2 C370 ( .A(pcout[80]), .B(cyc2), .Z(pcout_in[80]) );
  GTECH_AND2 C371 ( .A(pcout[79]), .B(cyc2), .Z(pcout_in[79]) );
  GTECH_AND2 C372 ( .A(pcout[78]), .B(cyc2), .Z(pcout_in[78]) );
  GTECH_AND2 C373 ( .A(pcout[77]), .B(cyc2), .Z(pcout_in[77]) );
  GTECH_AND2 C374 ( .A(pcout[76]), .B(cyc2), .Z(pcout_in[76]) );
  GTECH_AND2 C375 ( .A(pcout[75]), .B(cyc2), .Z(pcout_in[75]) );
  GTECH_AND2 C376 ( .A(pcout[74]), .B(cyc2), .Z(pcout_in[74]) );
  GTECH_AND2 C377 ( .A(pcout[73]), .B(cyc2), .Z(pcout_in[73]) );
  GTECH_AND2 C378 ( .A(pcout[72]), .B(cyc2), .Z(pcout_in[72]) );
  GTECH_AND2 C379 ( .A(pcout[71]), .B(cyc2), .Z(pcout_in[71]) );
  GTECH_AND2 C380 ( .A(pcout[70]), .B(cyc2), .Z(pcout_in[70]) );
  GTECH_AND2 C381 ( .A(pcout[69]), .B(cyc2), .Z(pcout_in[69]) );
  GTECH_AND2 C382 ( .A(pcout[68]), .B(cyc2), .Z(pcout_in[68]) );
  GTECH_AND2 C383 ( .A(pcout[67]), .B(cyc2), .Z(pcout_in[67]) );
  GTECH_AND2 C384 ( .A(pcout[66]), .B(cyc2), .Z(pcout_in[66]) );
  GTECH_AND2 C385 ( .A(pcout[65]), .B(cyc2), .Z(pcout_in[65]) );
  GTECH_AND2 C386 ( .A(pcout[64]), .B(cyc2), .Z(pcout_in[64]) );
  GTECH_AND2 C387 ( .A(pcout[63]), .B(cyc2), .Z(pcout_in[63]) );
  GTECH_AND2 C388 ( .A(pcout[62]), .B(cyc2), .Z(pcout_in[62]) );
  GTECH_AND2 C389 ( .A(pcout[61]), .B(cyc2), .Z(pcout_in[61]) );
  GTECH_AND2 C390 ( .A(pcout[60]), .B(cyc2), .Z(pcout_in[60]) );
  GTECH_AND2 C391 ( .A(pcout[59]), .B(cyc2), .Z(pcout_in[59]) );
  GTECH_AND2 C392 ( .A(pcout[58]), .B(cyc2), .Z(pcout_in[58]) );
  GTECH_AND2 C393 ( .A(pcout[57]), .B(cyc2), .Z(pcout_in[57]) );
  GTECH_AND2 C394 ( .A(pcout[56]), .B(cyc2), .Z(pcout_in[56]) );
  GTECH_AND2 C395 ( .A(pcout[55]), .B(cyc2), .Z(pcout_in[55]) );
  GTECH_AND2 C396 ( .A(pcout[54]), .B(cyc2), .Z(pcout_in[54]) );
  GTECH_AND2 C397 ( .A(pcout[53]), .B(cyc2), .Z(pcout_in[53]) );
  GTECH_AND2 C398 ( .A(pcout[52]), .B(cyc2), .Z(pcout_in[52]) );
  GTECH_AND2 C399 ( .A(pcout[51]), .B(cyc2), .Z(pcout_in[51]) );
  GTECH_AND2 C400 ( .A(pcout[50]), .B(cyc2), .Z(pcout_in[50]) );
  GTECH_AND2 C401 ( .A(pcout[49]), .B(cyc2), .Z(pcout_in[49]) );
  GTECH_AND2 C402 ( .A(pcout[48]), .B(cyc2), .Z(pcout_in[48]) );
  GTECH_AND2 C403 ( .A(pcout[47]), .B(cyc2), .Z(pcout_in[47]) );
  GTECH_AND2 C404 ( .A(pcout[46]), .B(cyc2), .Z(pcout_in[46]) );
  GTECH_AND2 C405 ( .A(pcout[45]), .B(cyc2), .Z(pcout_in[45]) );
  GTECH_AND2 C406 ( .A(pcout[44]), .B(cyc2), .Z(pcout_in[44]) );
  GTECH_AND2 C407 ( .A(pcout[43]), .B(cyc2), .Z(pcout_in[43]) );
  GTECH_AND2 C408 ( .A(pcout[42]), .B(cyc2), .Z(pcout_in[42]) );
  GTECH_AND2 C409 ( .A(pcout[41]), .B(cyc2), .Z(pcout_in[41]) );
  GTECH_AND2 C410 ( .A(pcout[40]), .B(cyc2), .Z(pcout_in[40]) );
  GTECH_AND2 C411 ( .A(pcout[39]), .B(cyc2), .Z(pcout_in[39]) );
  GTECH_AND2 C412 ( .A(pcout[38]), .B(cyc2), .Z(pcout_in[38]) );
  GTECH_AND2 C413 ( .A(pcout[37]), .B(cyc2), .Z(pcout_in[37]) );
  GTECH_AND2 C414 ( .A(pcout[36]), .B(cyc2), .Z(pcout_in[36]) );
  GTECH_AND2 C415 ( .A(pcout[35]), .B(cyc2), .Z(pcout_in[35]) );
  GTECH_AND2 C416 ( .A(pcout[34]), .B(cyc2), .Z(pcout_in[34]) );
  GTECH_AND2 C417 ( .A(pcout[33]), .B(cyc2), .Z(pcout_in[33]) );
  GTECH_AND2 C418 ( .A(pcout[32]), .B(cyc2), .Z(pcout_in[32]) );
  GTECH_AND2 C419 ( .A(pcout[31]), .B(cyc2), .Z(pcout_in[31]) );
  GTECH_AND2 C420 ( .A(pcout[30]), .B(x2_c2), .Z(pcout_in[30]) );
  GTECH_AND2 C421 ( .A(add_co31), .B(cyc3), .Z(add_cin) );
endmodule


module fpu_mul ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_mul, 
        mul_dest_rdy, mul_dest_rdya, fmul_clken_l, fmul_clken_l_buf1, arst_l, 
        grst_l, rclk, mul_pipe_active, m1stg_step, m6stg_fmul_in, m6stg_id_in, 
        mul_exc_out, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, 
        mul_exp_out, mul_frac_out, se_mul, se_mul64, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] m6stg_id_in;
  output [4:0] mul_exc_out;
  output [10:0] mul_exp_out;
  output [51:0] mul_frac_out;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_mul, mul_dest_rdy, mul_dest_rdya,
         fmul_clken_l, fmul_clken_l_buf1, arst_l, grst_l, rclk, se_mul,
         se_mul64, si;
  output mul_pipe_active, m1stg_step, m6stg_fmul_in, m6stg_fmul_dbl_dst,
         m6stg_fmuls, mul_sign_out, so;
  wire   m5stg_fracadd_cout, m5stg_frac_neq_0, m5stg_frac_dbl_nx,
         m5stg_frac_sng_nx, m3stg_expadd_eq_0, m3stg_expadd_lte_0_inv,
         m4stg_frac_105, mul_rst_l, m1stg_snan_sng_in1, m1stg_snan_dbl_in1,
         m1stg_snan_sng_in2, m1stg_snan_dbl_in2, m1stg_sngop, m1stg_dblop,
         m1stg_dblop_inv, m1stg_fmul, m1stg_fsmuld, m2stg_fmuls, m2stg_fmuld,
         m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda, m6stg_step,
         m5stg_in_of, m2stg_frac1_dbl_norm, m2stg_frac1_dbl_dnrm,
         m2stg_frac1_sng_norm, m2stg_frac1_sng_dnrm, m2stg_frac1_inf,
         m2stg_frac2_dbl_norm, m2stg_frac2_dbl_dnrm, m2stg_frac2_sng_norm,
         m2stg_frac2_sng_dnrm, m2stg_frac2_inf, m1stg_inf_zero_in,
         m1stg_inf_zero_in_dbl, m2stg_exp_expadd, m2stg_exp_0bff,
         m2stg_exp_017f, m2stg_exp_04ff, m2stg_exp_zero, m4stg_inc_exp_54,
         m4stg_inc_exp_55, m4stg_inc_exp_105, m4stg_left_shift_step,
         m4stg_right_shift_step, m5stg_to_0, m5stg_to_0_inv,
         mul_frac_out_fracadd, mul_frac_out_frac, mul_exp_out_exp_plus1,
         mul_exp_out_exp, scan_out_fpu_mul_ctl, m4stg_shl_54, m4stg_shl_55,
         scan_out_fpu_mul_exp_dp, scan_out_fpu_mul_frac_dp;
  wire   [12:0] m5stg_exp;
  wire   [5:0] m1stg_ld0_1;
  wire   [5:0] m1stg_ld0_2;
  wire   [12:0] m3stg_exp;
  wire   [6:0] m3stg_ld0_inv;
  wire   [12:0] m4stg_exp;
  wire   [32:0] m5stg_frac_32_0;
  wire   [6:0] m3bstg_ld0_inv;
  wire   [5:0] m4stg_sh_cnt_in;
  wire   [105:0] m4stg_frac;
  wire   [52:0] m2stg_frac1_array_in;
  wire   [52:0] m2stg_frac2_array_in;
  wire   [29:0] m4stg_frac_unused;

  fpu_mul_ctl fpu_mul_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_51(inq_in2[51]), .inq_in2_54(
        inq_in2[54]), .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(inq_op), .inq_mul(
        inq_mul), .inq_rnd_mode(inq_rnd_mode), .inq_id(inq_id), .inq_in1_63(
        inq_in1[63]), .inq_in2_63(inq_in2[63]), .mul_dest_rdy(mul_dest_rdy), 
        .mul_dest_rdya(mul_dest_rdya), .m5stg_exp(m5stg_exp), 
        .m5stg_fracadd_cout(m5stg_fracadd_cout), .m5stg_frac_neq_0(
        m5stg_frac_neq_0), .m5stg_frac_dbl_nx(m5stg_frac_dbl_nx), 
        .m5stg_frac_sng_nx(m5stg_frac_sng_nx), .m1stg_ld0_1(m1stg_ld0_1), 
        .m1stg_ld0_2(m1stg_ld0_2), .m3stg_exp(m3stg_exp), .m3stg_expadd_eq_0(
        m3stg_expadd_eq_0), .m3stg_expadd_lte_0_inv(m3stg_expadd_lte_0_inv), 
        .m3stg_ld0_inv(m3stg_ld0_inv[5:0]), .m4stg_exp(m4stg_exp), 
        .m4stg_frac_105(m4stg_frac_105), .m5stg_frac(m5stg_frac_32_0), 
        .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), .mul_pipe_active(
        mul_pipe_active), .m1stg_snan_sng_in1(m1stg_snan_sng_in1), 
        .m1stg_snan_dbl_in1(m1stg_snan_dbl_in1), .m1stg_snan_sng_in2(
        m1stg_snan_sng_in2), .m1stg_snan_dbl_in2(m1stg_snan_dbl_in2), 
        .m1stg_step(m1stg_step), .m1stg_sngop(m1stg_sngop), .m1stg_dblop(
        m1stg_dblop), .m1stg_dblop_inv(m1stg_dblop_inv), .m1stg_fmul(
        m1stg_fmul), .m1stg_fsmuld(m1stg_fsmuld), .m2stg_fmuls(m2stg_fmuls), 
        .m2stg_fmuld(m2stg_fmuld), .m2stg_fsmuld(m2stg_fsmuld), .m5stg_fmuls(
        m5stg_fmuls), .m5stg_fmuld(m5stg_fmuld), .m5stg_fmulda(m5stg_fmulda), 
        .m6stg_fmul_in(m6stg_fmul_in), .m6stg_id_in(m6stg_id_in), 
        .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), .m6stg_fmuls(m6stg_fmuls), 
        .m6stg_step(m6stg_step), .mul_sign_out(mul_sign_out), .m5stg_in_of(
        m5stg_in_of), .mul_exc_out(mul_exc_out), .m2stg_frac1_dbl_norm(
        m2stg_frac1_dbl_norm), .m2stg_frac1_dbl_dnrm(m2stg_frac1_dbl_dnrm), 
        .m2stg_frac1_sng_norm(m2stg_frac1_sng_norm), .m2stg_frac1_sng_dnrm(
        m2stg_frac1_sng_dnrm), .m2stg_frac1_inf(m2stg_frac1_inf), 
        .m2stg_frac2_dbl_norm(m2stg_frac2_dbl_norm), .m2stg_frac2_dbl_dnrm(
        m2stg_frac2_dbl_dnrm), .m2stg_frac2_sng_norm(m2stg_frac2_sng_norm), 
        .m2stg_frac2_sng_dnrm(m2stg_frac2_sng_dnrm), .m2stg_frac2_inf(
        m2stg_frac2_inf), .m1stg_inf_zero_in(m1stg_inf_zero_in), 
        .m1stg_inf_zero_in_dbl(m1stg_inf_zero_in_dbl), .m2stg_exp_expadd(
        m2stg_exp_expadd), .m2stg_exp_0bff(m2stg_exp_0bff), .m2stg_exp_017f(
        m2stg_exp_017f), .m2stg_exp_04ff(m2stg_exp_04ff), .m2stg_exp_zero(
        m2stg_exp_zero), .m3bstg_ld0_inv(m3bstg_ld0_inv), .m4stg_sh_cnt_in(
        m4stg_sh_cnt_in), .m4stg_inc_exp_54(m4stg_inc_exp_54), 
        .m4stg_inc_exp_55(m4stg_inc_exp_55), .m4stg_inc_exp_105(
        m4stg_inc_exp_105), .m4stg_left_shift_step(m4stg_left_shift_step), 
        .m4stg_right_shift_step(m4stg_right_shift_step), .m5stg_to_0(
        m5stg_to_0), .m5stg_to_0_inv(m5stg_to_0_inv), .mul_frac_out_fracadd(
        mul_frac_out_fracadd), .mul_frac_out_frac(mul_frac_out_frac), 
        .mul_exp_out_exp_plus1(mul_exp_out_exp_plus1), .mul_exp_out_exp(
        mul_exp_out_exp), .mula_rst_l(mul_rst_l), .se(se_mul), .si(si), .so(
        scan_out_fpu_mul_ctl) );
  fpu_mul_exp_dp fpu_mul_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .m6stg_step(m6stg_step), .m1stg_dblop(m1stg_dblop), 
        .m1stg_sngop(m1stg_sngop), .m2stg_exp_expadd(m2stg_exp_expadd), 
        .m2stg_exp_0bff(m2stg_exp_0bff), .m2stg_exp_017f(m2stg_exp_017f), 
        .m2stg_exp_04ff(m2stg_exp_04ff), .m2stg_exp_zero(m2stg_exp_zero), 
        .m1stg_fsmuld(m1stg_fsmuld), .m2stg_fmuld(m2stg_fmuld), .m2stg_fmuls(
        m2stg_fmuls), .m2stg_fsmuld(m2stg_fsmuld), .m3stg_ld0_inv(
        m3stg_ld0_inv), .m5stg_fracadd_cout(m5stg_fracadd_cout), 
        .mul_exp_out_exp_plus1(mul_exp_out_exp_plus1), .mul_exp_out_exp(
        mul_exp_out_exp), .m5stg_in_of(m5stg_in_of), .m5stg_fmuld(m5stg_fmuld), 
        .m5stg_to_0_inv(m5stg_to_0_inv), .m4stg_shl_54(m4stg_shl_54), 
        .m4stg_shl_55(m4stg_shl_55), .m4stg_inc_exp_54(m4stg_inc_exp_54), 
        .m4stg_inc_exp_55(m4stg_inc_exp_55), .m4stg_inc_exp_105(
        m4stg_inc_exp_105), .fmul_clken_l(fmul_clken_l_buf1), .rclk(rclk), 
        .m3stg_exp(m3stg_exp), .m3stg_expadd_eq_0(m3stg_expadd_eq_0), 
        .m3stg_expadd_lte_0_inv(m3stg_expadd_lte_0_inv), .m4stg_exp(m4stg_exp), 
        .m5stg_exp(m5stg_exp), .mul_exp_out(mul_exp_out), .se(se_mul), .si(
        scan_out_fpu_mul_ctl), .so(scan_out_fpu_mul_exp_dp) );
  fpu_mul_frac_dp fpu_mul_frac_dp ( .inq_in1(inq_in1[54:0]), .inq_in2(
        inq_in2[54:0]), .m6stg_step(m6stg_step), .m2stg_frac1_dbl_norm(
        m2stg_frac1_dbl_norm), .m2stg_frac1_dbl_dnrm(m2stg_frac1_dbl_dnrm), 
        .m2stg_frac1_sng_norm(m2stg_frac1_sng_norm), .m2stg_frac1_sng_dnrm(
        m2stg_frac1_sng_dnrm), .m2stg_frac1_inf(m2stg_frac1_inf), 
        .m1stg_snan_dbl_in1(m1stg_snan_dbl_in1), .m1stg_snan_sng_in1(
        m1stg_snan_sng_in1), .m2stg_frac2_dbl_norm(m2stg_frac2_dbl_norm), 
        .m2stg_frac2_dbl_dnrm(m2stg_frac2_dbl_dnrm), .m2stg_frac2_sng_norm(
        m2stg_frac2_sng_norm), .m2stg_frac2_sng_dnrm(m2stg_frac2_sng_dnrm), 
        .m2stg_frac2_inf(m2stg_frac2_inf), .m1stg_snan_dbl_in2(
        m1stg_snan_dbl_in2), .m1stg_snan_sng_in2(m1stg_snan_sng_in2), 
        .m1stg_inf_zero_in(m1stg_inf_zero_in), .m1stg_inf_zero_in_dbl(
        m1stg_inf_zero_in_dbl), .m1stg_dblop(m1stg_dblop), .m1stg_dblop_inv(
        m1stg_dblop_inv), .m4stg_frac(m4stg_frac), .m4stg_sh_cnt_in(
        m4stg_sh_cnt_in), .m3bstg_ld0_inv(m3bstg_ld0_inv), 
        .m4stg_left_shift_step(m4stg_left_shift_step), 
        .m4stg_right_shift_step(m4stg_right_shift_step), .m5stg_fmuls(
        m5stg_fmuls), .m5stg_fmulda(m5stg_fmulda), .mul_frac_out_fracadd(
        mul_frac_out_fracadd), .mul_frac_out_frac(mul_frac_out_frac), 
        .m5stg_in_of(m5stg_in_of), .m5stg_to_0(m5stg_to_0), .fmul_clken_l(
        fmul_clken_l), .rclk(rclk), .m2stg_frac1_array_in(m2stg_frac1_array_in), .m2stg_frac2_array_in(m2stg_frac2_array_in), .m1stg_ld0_1(m1stg_ld0_1), 
        .m1stg_ld0_2(m1stg_ld0_2), .m4stg_frac_105(m4stg_frac_105), 
        .m3stg_ld0_inv(m3stg_ld0_inv), .m4stg_shl_54(m4stg_shl_54), 
        .m4stg_shl_55(m4stg_shl_55), .m5stg_frac_32_0(m5stg_frac_32_0), 
        .m5stg_frac_dbl_nx(m5stg_frac_dbl_nx), .m5stg_frac_sng_nx(
        m5stg_frac_sng_nx), .m5stg_frac_neq_0(m5stg_frac_neq_0), 
        .m5stg_fracadd_cout(m5stg_fracadd_cout), .mul_frac_out(mul_frac_out), 
        .se(se_mul), .si(scan_out_fpu_mul_exp_dp), .so(
        scan_out_fpu_mul_frac_dp) );
  mul64 i_m4stg_frac ( .rs1_l({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, m2stg_frac1_array_in}), .rs2({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m2stg_frac2_array_in}), 
        .valid(m1stg_fmul), .areg({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .accreg({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .x2(1'b0), .out({m4stg_frac_unused, m4stg_frac}), 
        .rclk(rclk), .si(scan_out_fpu_mul_frac_dp), .so(so), .se(se_mul64), 
        .mul_rst_l(mul_rst_l), .mul_step(m6stg_step) );
endmodule


module dffr_SIZE8 ( din, clk, rst, q, se, si, so );
  input [7:0] din;
  output [7:0] q;
  input [7:0] si;
  output [7:0] so;
  input clk, rst, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21;
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C31 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({N13, N12, N11, N10, N9, 
        N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  GTECH_BUF B_1 ( .A(N5), .Z(N1) );
  SELECT_OP C32 ( .DATA1(si), .DATA2({N13, N12, N11, N10, N9, N8, N7, N6}), 
        .CONTROL1(N2), .CONTROL2(N3), .Z({N21, N20, N19, N18, N17, N16, N15, 
        N14}) );
  GTECH_BUF B_2 ( .A(se), .Z(N2) );
  GTECH_BUF B_3 ( .A(N4), .Z(N3) );
  GTECH_NOT I_0 ( .A(se), .Z(N4) );
  GTECH_NOT I_1 ( .A(rst), .Z(N5) );
endmodule


module dffr_SIZE3 ( din, clk, rst, q, se, si, so );
  input [2:0] din;
  output [2:0] q;
  input [2:0] si;
  output [2:0] so;
  input clk, rst, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11;
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C21 ( .DATA1({1'b0, 1'b0, 1'b0}), .DATA2(din), .CONTROL1(N0), 
        .CONTROL2(N1), .Z({N8, N7, N6}) );
  GTECH_BUF B_0 ( .A(rst), .Z(N0) );
  GTECH_BUF B_1 ( .A(N5), .Z(N1) );
  SELECT_OP C22 ( .DATA1(si), .DATA2({N8, N7, N6}), .CONTROL1(N2), .CONTROL2(
        N3), .Z({N11, N10, N9}) );
  GTECH_BUF B_2 ( .A(se), .Z(N2) );
  GTECH_BUF B_3 ( .A(N4), .Z(N3) );
  GTECH_NOT I_0 ( .A(se), .Z(N4) );
  GTECH_NOT I_1 ( .A(rst), .Z(N5) );
endmodule


module fpu_div_ctl ( inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, inq_op, div_exp1, div_dest_rdy, inq_rnd_mode, 
        inq_id, inq_in1_63, inq_in2_63, inq_div, div_exp_out, 
        div_frac_add_52_inva, div_frac_add_in1_neq_0, div_frac_out_54, 
        d6stg_frac_0, d6stg_frac_1, d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, 
        d6stg_frac_31, div_frac_out_53, div_expadd2_12, arst_l, grst_l, rclk, 
        div_pipe_active, d1stg_snan_sng_in1, d1stg_snan_dbl_in1, 
        d1stg_snan_sng_in2, d1stg_snan_dbl_in2, d1stg_step, d1stg_dblop, 
        d234stg_fdiv, d3stg_fdiv, d4stg_fdiv, d5stg_fdiva, d5stg_fdivb, 
        d5stg_fdivs, d5stg_fdivd, d6stg_fdiv, d6stg_fdivs, d6stg_fdivd, 
        d7stg_fdiv, d7stg_fdivd, d8stg_fdiv_in, d8stg_fdivs, d8stg_fdivd, 
        div_id_out_in, div_sign_out, div_exc_out, div_norm_frac_in1_dbl_norm, 
        div_norm_frac_in1_dbl_dnrm, div_norm_frac_in1_sng_norm, 
        div_norm_frac_in1_sng_dnrm, div_norm_frac_in2_dbl_norm, 
        div_norm_frac_in2_dbl_dnrm, div_norm_frac_in2_sng_norm, 
        div_norm_frac_in2_sng_dnrm, div_norm_inf, div_norm_qnan, div_norm_zero, 
        div_frac_add_in2_load, d6stg_frac_out_shl1, d6stg_frac_out_nosh, 
        div_frac_add_in1_add, div_frac_add_in1_load, d7stg_rndup_inv, 
        d7stg_to_0, d7stg_to_0_inv, div_frac_out_add_in1, div_frac_out_add, 
        div_frac_out_shl1_dbl, div_frac_out_shl1_sng, div_frac_out_of, 
        div_frac_out_load, div_expadd1_in1_dbl, div_expadd1_in1_sng, 
        div_expadd1_in2_exp_in2_dbl, div_expadd1_in2_exp_in2_sng, 
        div_exp1_expadd1, div_exp1_0835, div_exp1_0118, div_exp1_zero, 
        div_exp1_load, div_expadd2_in1_exp_out, div_expadd2_no_decr_inv, 
        div_expadd2_cin, div_exp_out_expadd22_inv, div_exp_out_expadd2, 
        div_exp_out_of, div_exp_out_exp_out, div_exp_out_load, se, si, so );
  input [7:0] inq_op;
  input [12:0] div_exp1;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [12:0] div_exp_out;
  output [9:0] div_id_out_in;
  output [4:0] div_exc_out;
  input inq_in1_51, inq_in1_54, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs,
         inq_in2_51, inq_in2_54, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs,
         div_dest_rdy, inq_in1_63, inq_in2_63, inq_div, div_frac_add_52_inva,
         div_frac_add_in1_neq_0, div_frac_out_54, d6stg_frac_0, d6stg_frac_1,
         d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, d6stg_frac_31,
         div_frac_out_53, div_expadd2_12, arst_l, grst_l, rclk, se, si;
  output div_pipe_active, d1stg_snan_sng_in1, d1stg_snan_dbl_in1,
         d1stg_snan_sng_in2, d1stg_snan_dbl_in2, d1stg_step, d1stg_dblop,
         d234stg_fdiv, d3stg_fdiv, d4stg_fdiv, d5stg_fdiva, d5stg_fdivb,
         d5stg_fdivs, d5stg_fdivd, d6stg_fdiv, d6stg_fdivs, d6stg_fdivd,
         d7stg_fdiv, d7stg_fdivd, d8stg_fdiv_in, d8stg_fdivs, d8stg_fdivd,
         div_sign_out, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm,
         div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm,
         div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm,
         div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf,
         div_norm_qnan, div_norm_zero, div_frac_add_in2_load,
         d6stg_frac_out_shl1, d6stg_frac_out_nosh, div_frac_add_in1_add,
         div_frac_add_in1_load, d7stg_rndup_inv, d7stg_to_0, d7stg_to_0_inv,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, div_frac_out_load,
         div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl,
         div_expadd1_in2_exp_in2_sng, div_exp1_expadd1, div_exp1_0835,
         div_exp1_0118, div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd22_inv,
         div_exp_out_expadd2, div_exp_out_of, div_exp_out_exp_out,
         div_exp_out_load, so;
  wire   div_ctl_rst_l, reset, div_frac_in1_51, div_frac_in1_54,
         div_frac_in1_53_0_neq_0, div_frac_in1_50_0_neq_0,
         div_frac_in1_53_32_neq_0, div_exp_in1_exp_eq_0,
         div_exp_in1_exp_neq_ffs, div_frac_in2_51, div_frac_in2_54,
         div_frac_in2_53_0_neq_0, div_frac_in2_50_0_neq_0,
         div_frac_in2_53_32_neq_0, div_exp_in2_exp_eq_0,
         div_exp_in2_exp_neq_ffs, d1stg_denorm_sng_in1, d1stg_denorm_dbl_in1,
         d1stg_denorm_sng_in2, d1stg_denorm_dbl_in2, d2stg_denorm_sng_in2,
         d2stg_denorm_dbl_in2, d1stg_norm_sng_in1, d1stg_norm_dbl_in1,
         d1stg_norm_sng_in2, d1stg_norm_dbl_in2, d2stg_norm_sng_in2,
         d2stg_norm_dbl_in2, d1stg_qnan_sng_in1, d1stg_qnan_dbl_in1,
         d1stg_qnan_sng_in2, d1stg_qnan_dbl_in2, d1stg_snan_in1,
         d1stg_snan_in2, d1stg_qnan_in1, d1stg_qnan_in2, d1stg_nan_sng_in1,
         d1stg_nan_dbl_in1, d1stg_nan_sng_in2, d1stg_nan_dbl_in2,
         d1stg_nan_in1, d1stg_nan_in2, d1stg_nan_in, d2stg_snan_in1,
         d2stg_snan_in2, d2stg_qnan_in1, d2stg_qnan_in2, d2stg_nan_in2,
         d2stg_nan_in, d1stg_inf_sng_in1, d1stg_inf_dbl_in1, d1stg_inf_sng_in2,
         d1stg_inf_dbl_in2, d1stg_inf_in1, d1stg_inf_in2, d1stg_inf_in,
         d1stg_2inf_in, d2stg_inf_in1, d2stg_inf_in2, d2stg_2inf_in,
         d1stg_infnan_sng_in1, d1stg_infnan_dbl_in1, d1stg_infnan_sng_in2,
         d1stg_infnan_dbl_in2, d1stg_infnan_in1, d1stg_infnan_in2,
         d1stg_infnan_in, d2stg_infnan_in1, d2stg_infnan_in2, d2stg_infnan_in,
         d1stg_zero_in1, d1stg_zero_in2, d1stg_zero_in, d1stg_2zero_in,
         d2stg_zero_in1, d2stg_zero_in2, d2stg_zero_in, d2stg_2zero_in,
         d1stg_div, divs_cnt_lt_23, divd_cnt_lt_52, d1stg_hold,
         divs_cnt_lt_23a, divd_cnt_lt_52a, d1stg_holda, d1stg_stepa,
         d1stg_div_in, d234stg_fdiv_in, d6stg_step, d5stg_step, d5stg_fdivb_in,
         N0, N1, d8stg_step, N2, d8stg_hold, div_pipe_active_in, d1stg_sign1,
         d1stg_sign2, N3, d1stg_sign, div_bkend_step, div_cnt_step,
         div_cnt_lt_step, N4, divs_cnt_lt_23_in, N5, divd_cnt_lt_52_in,
         div_exc_step, div_of_mask_in, div_of_mask, div_nv_out_in,
         div_dz_out_in, N6, d7stg_in_of, d7stg_rndup, div_of_out_tmp1_in,
         div_of_out_tmp1, div_of_out_tmp2, div_out_52_inv, d7stg_grd,
         d7stg_stk, div_uf_out_in, div_nx_out_in, div_nx_out, d1stg_spc_rslt,
         d7stg_lsb_in, d7stg_grd_in, d7stg_stk_in, d7stg_lsb, N7,
         div_expadd1_in1_dbl_in, div_expadd1_in1_sng_in, d2stg_max_exp,
         d2stg_zero_exp, div_expadd2_in1_exp_out_in, N8, N9, N10,
         div_expadd2_no_decr_inv_in, div_expadd2_no_decr_load,
         div_exp_out_zero, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279,
         N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290,
         N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301,
         N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312,
         N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323,
         N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367,
         N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378,
         N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422,
         N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433,
         N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444,
         N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455,
         N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477,
         N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510,
         N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521,
         N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532,
         N533, N534, N535, N536, N537, N538, N539, N540, net12866, net12867,
         net12868, net12869, net12870, net12871, net12872, net12873, net12874,
         net12875, net12876, net12877, net12878, net12879, net12880, net12881,
         net12882, net12883, net12884, net12885, net12886, net12887, net12888,
         net12889, net12890, net12891, net12892, net12893, net12894, net12895,
         net12896, net12897, net12898, net12899, net12900, net12901, net12902,
         net12903, net12904, net12905, net12906, net12907, net12908, net12909,
         net12910, net12911, net12912, net12913, net12914, net12915, net12916,
         net12917, net12918, net12919, net12920, net12921, net12922, net12923,
         net12924, net12925, net12926, net12927, net12928, net12929, net12930,
         net12931, net12932, net12933, net12934, net12935, net12936, net12937,
         net12938, net12939, net12940, net12941, net12942, net12943, net12944,
         net12945, net12946, net12947, net12948, net12949, net12950, net12951,
         net12952, net12953, net12954, net12955, net12956, net12957, net12958,
         net12959, net12960, net12961, net12962, net12963, net12964, net12965,
         net12966, net12967, net12968, net12969, net12970, net12971, net12972,
         net12973, net12974, net12975, net12976, net12977, net12978, net12979,
         net12980, net12981, net12982, net12983, net12984, net12985, net12986,
         net12987, net12988, net12989, net12990, net12991, net12992, net12993;
  wire   [4:0] d1stg_sngopa;
  wire   [4:0] d1stg_dblopa;
  wire   [7:0] d1stg_op_in;
  wire   [7:0] d1stg_op;
  wire   [2:2] d1stg_opdec;
  wire   [2:2] d2stg_opdec;
  wire   [1:0] d3stg_opdec;
  wire   [1:0] d4stg_opdec;
  wire   [2:2] d5stg_opdec;
  wire   [5:0] div_cnt;
  wire   [2:0] d6stg_opdec_in;
  wire   [1:1] d7stg_opdec;
  wire   [2:2] d8stg_opdec;
  wire   [1:0] d1stg_rnd_mode;
  wire   [4:0] d1stg_id;
  wire   [1:0] div_rnd_mode;
  wire   [9:0] div_id_out;
  wire   [5:0] div_cnt_plus1;
  wire   [5:0] div_cnt_in;

  dffrl_async_SIZE1 dffrl_div_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(div_ctl_rst_l), .se(se), .si(net12993) );
  dffe_SIZE1 i_div_frac_in1_51 ( .din(inq_in1_51), .en(d1stg_step), .clk(rclk), 
        .q(div_frac_in1_51), .se(se), .si(net12992) );
  dffe_SIZE1 i_div_frac_in1_54 ( .din(inq_in1_54), .en(d1stg_step), .clk(rclk), 
        .q(div_frac_in1_54), .se(se), .si(net12991) );
  dffe_SIZE1 i_div_frac_in1_53_0_neq_0 ( .din(inq_in1_53_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_53_0_neq_0), .se(se), .si(
        net12990) );
  dffe_SIZE1 i_div_frac_in1_50_0_neq_0 ( .din(inq_in1_50_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_50_0_neq_0), .se(se), .si(
        net12989) );
  dffe_SIZE1 i_div_frac_in1_53_32_neq_0 ( .din(inq_in1_53_32_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in1_53_32_neq_0), .se(se), .si(
        net12988) );
  dffe_SIZE1 i_div_exp_in1_exp_eq_0 ( .din(inq_in1_exp_eq_0), .en(d1stg_step), 
        .clk(rclk), .q(div_exp_in1_exp_eq_0), .se(se), .si(net12987) );
  dffe_SIZE1 i_div_exp_in1_exp_neq_ffs ( .din(inq_in1_exp_neq_ffs), .en(
        d1stg_step), .clk(rclk), .q(div_exp_in1_exp_neq_ffs), .se(se), .si(
        net12986) );
  dffe_SIZE1 i_div_frac_in2_51 ( .din(inq_in2_51), .en(d1stg_step), .clk(rclk), 
        .q(div_frac_in2_51), .se(se), .si(net12985) );
  dffe_SIZE1 i_div_frac_in2_54 ( .din(inq_in2_54), .en(d1stg_step), .clk(rclk), 
        .q(div_frac_in2_54), .se(se), .si(net12984) );
  dffe_SIZE1 i_div_frac_in2_53_0_neq_0 ( .din(inq_in2_53_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_53_0_neq_0), .se(se), .si(
        net12983) );
  dffe_SIZE1 i_div_frac_in2_50_0_neq_0 ( .din(inq_in2_50_0_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_50_0_neq_0), .se(se), .si(
        net12982) );
  dffe_SIZE1 i_div_frac_in2_53_32_neq_0 ( .din(inq_in2_53_32_neq_0), .en(
        d1stg_step), .clk(rclk), .q(div_frac_in2_53_32_neq_0), .se(se), .si(
        net12981) );
  dffe_SIZE1 i_div_exp_in2_exp_eq_0 ( .din(inq_in2_exp_eq_0), .en(d1stg_step), 
        .clk(rclk), .q(div_exp_in2_exp_eq_0), .se(se), .si(net12980) );
  dffe_SIZE1 i_div_exp_in2_exp_neq_ffs ( .din(inq_in2_exp_neq_ffs), .en(
        d1stg_step), .clk(rclk), .q(div_exp_in2_exp_neq_ffs), .se(se), .si(
        net12979) );
  dff_SIZE1 i_d2stg_denorm_sng_in2 ( .din(d1stg_denorm_sng_in2), .clk(rclk), 
        .q(d2stg_denorm_sng_in2), .se(se), .si(net12978) );
  dff_SIZE1 i_d2stg_denorm_dbl_in2 ( .din(d1stg_denorm_dbl_in2), .clk(rclk), 
        .q(d2stg_denorm_dbl_in2), .se(se), .si(net12977) );
  dff_SIZE1 i_d2stg_norm_sng_in2 ( .din(d1stg_norm_sng_in2), .clk(rclk), .q(
        d2stg_norm_sng_in2), .se(se), .si(net12976) );
  dff_SIZE1 i_d2stg_norm_dbl_in2 ( .din(d1stg_norm_dbl_in2), .clk(rclk), .q(
        d2stg_norm_dbl_in2), .se(se), .si(net12975) );
  dff_SIZE1 i_d2stg_snan_in1 ( .din(d1stg_snan_in1), .clk(rclk), .q(
        d2stg_snan_in1), .se(se), .si(net12974) );
  dff_SIZE1 i_d2stg_snan_in2 ( .din(d1stg_snan_in2), .clk(rclk), .q(
        d2stg_snan_in2), .se(se), .si(net12973) );
  dff_SIZE1 i_d2stg_qnan_in1 ( .din(d1stg_qnan_in1), .clk(rclk), .q(
        d2stg_qnan_in1), .se(se), .si(net12972) );
  dff_SIZE1 i_d2stg_qnan_in2 ( .din(d1stg_qnan_in2), .clk(rclk), .q(
        d2stg_qnan_in2), .se(se), .si(net12971) );
  dff_SIZE1 i_d2stg_nan_in2 ( .din(d1stg_nan_in2), .clk(rclk), .q(
        d2stg_nan_in2), .se(se), .si(net12970) );
  dff_SIZE1 i_d2stg_nan_in ( .din(d1stg_nan_in), .clk(rclk), .q(d2stg_nan_in), 
        .se(se), .si(net12969) );
  dff_SIZE1 i_d2stg_inf_in1 ( .din(d1stg_inf_in1), .clk(rclk), .q(
        d2stg_inf_in1), .se(se), .si(net12968) );
  dff_SIZE1 i_d2stg_inf_in2 ( .din(d1stg_inf_in2), .clk(rclk), .q(
        d2stg_inf_in2), .se(se), .si(net12967) );
  dff_SIZE1 i_d2stg_2inf_in ( .din(d1stg_2inf_in), .clk(rclk), .q(
        d2stg_2inf_in), .se(se), .si(net12966) );
  dff_SIZE1 i_d2stg_infnan_in1 ( .din(d1stg_infnan_in1), .clk(rclk), .q(
        d2stg_infnan_in1), .se(se), .si(net12965) );
  dff_SIZE1 i_d2stg_infnan_in2 ( .din(d1stg_infnan_in2), .clk(rclk), .q(
        d2stg_infnan_in2), .se(se), .si(net12964) );
  dff_SIZE1 i_d2stg_infnan_in ( .din(d1stg_infnan_in), .clk(rclk), .q(
        d2stg_infnan_in), .se(se), .si(net12963) );
  dff_SIZE1 i_d2stg_zero_in1 ( .din(d1stg_zero_in1), .clk(rclk), .q(
        d2stg_zero_in1), .se(se), .si(net12962) );
  dff_SIZE1 i_d2stg_zero_in2 ( .din(d1stg_zero_in2), .clk(rclk), .q(
        d2stg_zero_in2), .se(se), .si(net12961) );
  dff_SIZE1 i_d2stg_zero_in ( .din(d1stg_zero_in), .clk(rclk), .q(
        d2stg_zero_in), .se(se), .si(net12960) );
  dff_SIZE1 i_d2stg_2zero_in ( .din(d1stg_2zero_in), .clk(rclk), .q(
        d2stg_2zero_in), .se(se), .si(net12959) );
  dffr_SIZE8 i_d1stg_op ( .din(d1stg_op_in), .clk(rclk), .rst(reset), .q(
        d1stg_op), .se(se), .si({net12951, net12952, net12953, net12954, 
        net12955, net12956, net12957, net12958}) );
  dffr_SIZE1 i_d1stg_div ( .din(d1stg_div_in), .clk(rclk), .rst(reset), .q(
        d1stg_div), .se(se), .si(net12950) );
  dffe_SIZE5 i_d1stg_sngopa ( .din({inq_op[0], inq_op[0], inq_op[0], inq_op[0], 
        inq_op[0]}), .en(d1stg_stepa), .clk(rclk), .q(d1stg_sngopa), .se(se), 
        .si({net12945, net12946, net12947, net12948, net12949}) );
  dffe_SIZE1 i_d1stg_dblop ( .din(inq_op[1]), .en(d1stg_stepa), .clk(rclk), 
        .q(d1stg_dblop), .se(se), .si(net12944) );
  dffe_SIZE5 i_d1stg_dblopa ( .din({inq_op[1], inq_op[1], inq_op[1], inq_op[1], 
        inq_op[1]}), .en(d1stg_stepa), .clk(rclk), .q(d1stg_dblopa), .se(se), 
        .si({net12939, net12940, net12941, net12942, net12943}) );
  dffr_SIZE3 i_d2stg_opdec ( .din({d1stg_opdec[2], N22, N31}), .clk(rclk), 
        .rst(reset), .q({d2stg_opdec[2], div_expadd1_in2_exp_in2_sng, 
        div_expadd1_in2_exp_in2_dbl}), .se(se), .si({net12936, net12937, 
        net12938}) );
  dffr_SIZE1 i_d234stg_fdiv ( .din(d234stg_fdiv_in), .clk(rclk), .rst(reset), 
        .q(d234stg_fdiv), .se(se), .si(net12935) );
  dffr_SIZE3 i_d3stg_opdec ( .din({d2stg_opdec[2], div_expadd1_in2_exp_in2_sng, 
        div_expadd1_in2_exp_in2_dbl}), .clk(rclk), .rst(reset), .q({d3stg_fdiv, 
        d3stg_opdec}), .se(se), .si({net12932, net12933, net12934}) );
  dffr_SIZE3 i_d4stg_opdec ( .din({d3stg_fdiv, d3stg_opdec}), .clk(rclk), 
        .rst(reset), .q({d4stg_fdiv, d4stg_opdec}), .se(se), .si({net12929, 
        net12930, net12931}) );
  dffre_SIZE3 i_d5stg_opdec ( .din({d4stg_fdiv, d4stg_opdec}), .rst(reset), 
        .en(d5stg_step), .clk(rclk), .q({d5stg_opdec[2], d5stg_fdivs, 
        d5stg_fdivd}), .se(se), .si({net12926, net12927, net12928}) );
  dffre_SIZE1 i_d5stg_fdiva ( .din(d4stg_fdiv), .rst(reset), .en(d5stg_step), 
        .clk(rclk), .q(d5stg_fdiva), .se(se), .si(net12925) );
  dff_SIZE1 i_d5stg_fdivb ( .din(d5stg_fdivb_in), .clk(rclk), .q(d5stg_fdivb), 
        .se(se), .si(net12924) );
  EQ_UNS_OP eq_1308_3 ( .A(div_cnt), .B(div_exp1), .Z(N0) );
  EQ_UNS_OP eq_1308_4 ( .A(div_cnt), .B(div_exp1), .Z(N1) );
  dffr_SIZE3 i_d6stg_opdec ( .din(d6stg_opdec_in), .clk(rclk), .rst(reset), 
        .q({d6stg_fdiv, d6stg_fdivs, d6stg_fdivd}), .se(se), .si({net12921, 
        net12922, net12923}) );
  dffr_SIZE3 i_d7stg_opdec ( .din({d6stg_fdiv, d6stg_fdivs, d6stg_fdivd}), 
        .clk(rclk), .rst(reset), .q({d7stg_fdiv, d7stg_opdec[1], d7stg_fdivd}), 
        .se(se), .si({net12918, net12919, net12920}) );
  dffre_SIZE3 i_d8stg_opdec ( .din({d7stg_fdiv, d7stg_opdec[1], d7stg_fdivd}), 
        .rst(reset), .en(d8stg_step), .clk(rclk), .q({d8stg_opdec[2], 
        d8stg_fdivs, d8stg_fdivd}), .se(se), .si({net12915, net12916, net12917}) );
  dffre_SIZE1 i_div_pipe_active ( .din(div_pipe_active_in), .rst(reset), .en(
        1'b1), .clk(rclk), .q(div_pipe_active), .se(se), .si(net12914) );
  dffe_SIZE2 i_d1stg_rnd_mode ( .din(inq_rnd_mode), .en(d1stg_stepa), .clk(
        rclk), .q(d1stg_rnd_mode), .se(se), .si({net12912, net12913}) );
  dffe_SIZE5 i_d1stg_id ( .din(inq_id), .en(d1stg_stepa), .clk(rclk), .q(
        d1stg_id), .se(se), .si({net12907, net12908, net12909, net12910, 
        net12911}) );
  dffe_SIZE1 i_d1stg_sign1 ( .din(inq_in1_63), .en(d1stg_stepa), .clk(rclk), 
        .q(d1stg_sign1), .se(se), .si(net12906) );
  dffe_SIZE1 i_d1stg_sign2 ( .din(inq_in2_63), .en(d1stg_stepa), .clk(rclk), 
        .q(d1stg_sign2), .se(se), .si(net12905) );
  dffe_SIZE2 i_div_rnd_mode ( .din(d1stg_rnd_mode), .en(div_bkend_step), .clk(
        rclk), .q(div_rnd_mode), .se(se), .si({net12903, net12904}) );
  dff_SIZE10 i_div_id_out ( .din(div_id_out_in), .clk(rclk), .q(div_id_out), 
        .se(se), .si({net12893, net12894, net12895, net12896, net12897, 
        net12898, net12899, net12900, net12901, net12902}) );
  dffe_SIZE1 i_div_sign_out ( .din(d1stg_sign), .en(div_bkend_step), .clk(rclk), .q(div_sign_out), .se(se), .si(net12892) );
  dffre_SIZE6 i_div_cnt ( .din(div_cnt_in), .rst(reset), .en(div_cnt_step), 
        .clk(rclk), .q(div_cnt), .se(se), .si({net12886, net12887, net12888, 
        net12889, net12890, net12891}) );
  LT_UNS_OP lt_1579 ( .A(div_cnt_plus1), .B({1'b1, 1'b0, 1'b1, 1'b1, 1'b1}), 
        .Z(N4) );
  dffre_SIZE1 i_divs_cnt_lt_23 ( .din(divs_cnt_lt_23_in), .rst(reset), .en(
        div_cnt_lt_step), .clk(rclk), .q(divs_cnt_lt_23), .se(se), .si(
        net12885) );
  dffre_SIZE1 i_divs_cnt_lt_23a ( .din(divs_cnt_lt_23_in), .rst(reset), .en(
        div_cnt_lt_step), .clk(rclk), .q(divs_cnt_lt_23a), .se(se), .si(
        net12884) );
  LT_UNS_OP lt_1608 ( .A(div_cnt_plus1), .B({1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 
        1'b0}), .Z(N5) );
  dffre_SIZE1 i_divd_cnt_lt_52 ( .din(divd_cnt_lt_52_in), .rst(reset), .en(
        div_cnt_lt_step), .clk(rclk), .q(divd_cnt_lt_52), .se(se), .si(
        net12883) );
  dffre_SIZE1 i_divd_cnt_lt_52a ( .din(divd_cnt_lt_52_in), .rst(reset), .en(
        div_cnt_lt_step), .clk(rclk), .q(divd_cnt_lt_52a), .se(se), .si(
        net12882) );
  dffe_SIZE1 i_div_of_mask ( .din(div_of_mask_in), .en(div_exc_step), .clk(
        rclk), .q(div_of_mask), .se(se), .si(net12881) );
  dffe_SIZE1 i_div_nv_out ( .din(div_nv_out_in), .en(div_exc_step), .clk(rclk), 
        .q(div_exc_out[4]), .se(se), .si(net12880) );
  dffe_SIZE1 i_div_dz_out ( .din(div_dz_out_in), .en(div_exc_step), .clk(rclk), 
        .q(div_exc_out[1]), .se(se), .si(net12879) );
  dffe_SIZE1 i_div_of_out_tmp1 ( .din(div_of_out_tmp1_in), .en(d7stg_fdiv), 
        .clk(rclk), .q(div_of_out_tmp1), .se(se), .si(net12878) );
  dffe_SIZE1 i_div_of_out_tmp2 ( .din(d7stg_in_of), .en(d7stg_fdiv), .clk(rclk), .q(div_of_out_tmp2), .se(se), .si(net12877) );
  dffe_SIZE1 i_div_out_52_inv ( .din(div_frac_add_52_inva), .en(d7stg_fdiv), 
        .clk(rclk), .q(div_out_52_inv), .se(se), .si(net12876) );
  dffe_SIZE1 i_div_uf_out ( .din(div_uf_out_in), .en(d7stg_fdiv), .clk(rclk), 
        .q(div_exc_out[2]), .se(se), .si(net12875) );
  dffe_SIZE1 i_div_nx_out ( .din(div_nx_out_in), .en(d7stg_fdiv), .clk(rclk), 
        .q(div_nx_out), .se(se), .si(net12874) );
  dffe_SIZE1 i_d7stg_lsb ( .din(d7stg_lsb_in), .en(d6stg_fdiv), .clk(rclk), 
        .q(d7stg_lsb), .se(se), .si(net12873) );
  dffe_SIZE1 i_d7stg_grd ( .din(d7stg_grd_in), .en(d6stg_fdiv), .clk(rclk), 
        .q(d7stg_grd), .se(se), .si(net12872) );
  dffe_SIZE1 i_d7stg_stk ( .din(d7stg_stk_in), .en(d6stg_fdiv), .clk(rclk), 
        .q(d7stg_stk), .se(se), .si(net12871) );
  dff_SIZE1 i_div_expadd1_in1_dbl ( .din(div_expadd1_in1_dbl_in), .clk(rclk), 
        .q(div_expadd1_in1_dbl), .se(se), .si(net12870) );
  dff_SIZE1 i_div_expadd1_in1_sng ( .din(div_expadd1_in1_sng_in), .clk(rclk), 
        .q(div_expadd1_in1_sng), .se(se), .si(net12869) );
  dffr_SIZE1 i_div_expadd2_in1_exp_out ( .din(div_expadd2_in1_exp_out_in), 
        .clk(rclk), .rst(reset), .q(div_expadd2_in1_exp_out), .se(se), .si(
        net12868) );
  EQ_UNS_OP eq_2107 ( .A(div_exp1[11:0]), .B({N8, N9, d5stg_fdivs, N8, 1'b0, 
        N8}), .Z(N10) );
  dffe_SIZE1 i_div_expadd2_no_decr_inv ( .din(div_expadd2_no_decr_inv_in), 
        .en(div_expadd2_no_decr_load), .clk(rclk), .q(div_expadd2_no_decr_inv), 
        .se(se), .si(net12867) );
  GTECH_NOT I_0 ( .A(d1stg_op[6]), .Z(N11) );
  GTECH_NOT I_1 ( .A(d1stg_op[3]), .Z(N12) );
  GTECH_NOT I_2 ( .A(d1stg_op[2]), .Z(N13) );
  GTECH_NOT I_3 ( .A(d1stg_op[0]), .Z(N14) );
  GTECH_OR2 C171 ( .A(N11), .B(d1stg_op[7]), .Z(N15) );
  GTECH_OR2 C172 ( .A(d1stg_op[5]), .B(N15), .Z(N16) );
  GTECH_OR2 C173 ( .A(d1stg_op[4]), .B(N16), .Z(N17) );
  GTECH_OR2 C174 ( .A(N12), .B(N17), .Z(N18) );
  GTECH_OR2 C175 ( .A(N13), .B(N18), .Z(N19) );
  GTECH_OR2 C176 ( .A(d1stg_op[1]), .B(N19), .Z(N20) );
  GTECH_OR2 C177 ( .A(N14), .B(N20), .Z(N21) );
  GTECH_NOT I_4 ( .A(N21), .Z(N22) );
  GTECH_NOT I_5 ( .A(d1stg_op[1]), .Z(N23) );
  GTECH_OR2 C183 ( .A(N11), .B(d1stg_op[7]), .Z(N24) );
  GTECH_OR2 C184 ( .A(d1stg_op[5]), .B(N24), .Z(N25) );
  GTECH_OR2 C185 ( .A(d1stg_op[4]), .B(N25), .Z(N26) );
  GTECH_OR2 C186 ( .A(N12), .B(N26), .Z(N27) );
  GTECH_OR2 C187 ( .A(N13), .B(N27), .Z(N28) );
  GTECH_OR2 C188 ( .A(N23), .B(N28), .Z(N29) );
  GTECH_OR2 C189 ( .A(d1stg_op[0]), .B(N29), .Z(N30) );
  GTECH_NOT I_6 ( .A(N30), .Z(N31) );
  GTECH_AND2 C191 ( .A(d1stg_id[3]), .B(d1stg_id[4]), .Z(N32) );
  GTECH_AND2 C192 ( .A(d1stg_id[2]), .B(N32), .Z(N33) );
  GTECH_NOT I_7 ( .A(d1stg_id[4]), .Z(N34) );
  GTECH_NOT I_8 ( .A(d1stg_id[3]), .Z(N35) );
  GTECH_OR2 C195 ( .A(N35), .B(N34), .Z(N36) );
  GTECH_OR2 C196 ( .A(d1stg_id[2]), .B(N36), .Z(N37) );
  GTECH_NOT I_9 ( .A(N37), .Z(N38) );
  GTECH_NOT I_10 ( .A(d1stg_id[2]), .Z(N39) );
  GTECH_OR2 C200 ( .A(d1stg_id[3]), .B(N34), .Z(N40) );
  GTECH_OR2 C201 ( .A(N39), .B(N40), .Z(N41) );
  GTECH_NOT I_11 ( .A(N41), .Z(N42) );
  GTECH_OR2 C204 ( .A(d1stg_id[3]), .B(N34), .Z(N43) );
  GTECH_OR2 C205 ( .A(d1stg_id[2]), .B(N43), .Z(N44) );
  GTECH_NOT I_12 ( .A(N44), .Z(N45) );
  GTECH_OR2 C209 ( .A(N35), .B(d1stg_id[4]), .Z(N46) );
  GTECH_OR2 C210 ( .A(N39), .B(N46), .Z(N47) );
  GTECH_NOT I_13 ( .A(N47), .Z(N48) );
  GTECH_OR2 C213 ( .A(N35), .B(d1stg_id[4]), .Z(N49) );
  GTECH_OR2 C214 ( .A(d1stg_id[2]), .B(N49), .Z(N50) );
  GTECH_NOT I_14 ( .A(N50), .Z(N51) );
  GTECH_OR2 C217 ( .A(d1stg_id[3]), .B(d1stg_id[4]), .Z(N52) );
  GTECH_OR2 C218 ( .A(N39), .B(N52), .Z(N53) );
  GTECH_NOT I_15 ( .A(N53), .Z(N54) );
  GTECH_OR2 C220 ( .A(d1stg_id[3]), .B(d1stg_id[4]), .Z(N55) );
  GTECH_OR2 C221 ( .A(d1stg_id[2]), .B(N55), .Z(N56) );
  GTECH_NOT I_16 ( .A(N56), .Z(N57) );
  GTECH_OR2 C223 ( .A(div_cnt[4]), .B(div_cnt[5]), .Z(N58) );
  GTECH_OR2 C224 ( .A(div_cnt[3]), .B(N58), .Z(N59) );
  GTECH_OR2 C225 ( .A(div_cnt[2]), .B(N59), .Z(N60) );
  GTECH_OR2 C226 ( .A(div_cnt[1]), .B(N60), .Z(N61) );
  GTECH_OR2 C227 ( .A(div_cnt[0]), .B(N61), .Z(N62) );
  GTECH_NOT I_17 ( .A(N62), .Z(N63) );
  GTECH_OR2 C229 ( .A(div_cnt[4]), .B(div_cnt[5]), .Z(N64) );
  GTECH_OR2 C230 ( .A(div_cnt[3]), .B(N64), .Z(N65) );
  GTECH_OR2 C231 ( .A(div_cnt[2]), .B(N65), .Z(N66) );
  GTECH_OR2 C232 ( .A(div_cnt[1]), .B(N66), .Z(N67) );
  GTECH_OR2 C233 ( .A(div_cnt[0]), .B(N67), .Z(N68) );
  GTECH_NOT I_18 ( .A(N68), .Z(N69) );
  GTECH_OR2 C235 ( .A(div_cnt[4]), .B(div_cnt[5]), .Z(N70) );
  GTECH_OR2 C236 ( .A(div_cnt[3]), .B(N70), .Z(N71) );
  GTECH_OR2 C237 ( .A(div_cnt[2]), .B(N71), .Z(N72) );
  GTECH_OR2 C238 ( .A(div_cnt[1]), .B(N72), .Z(N73) );
  GTECH_OR2 C239 ( .A(div_cnt[0]), .B(N73), .Z(N74) );
  GTECH_NOT I_19 ( .A(N74), .Z(N75) );
  GTECH_OR2 C241 ( .A(div_cnt[4]), .B(div_cnt[5]), .Z(N76) );
  GTECH_OR2 C242 ( .A(div_cnt[3]), .B(N76), .Z(N77) );
  GTECH_OR2 C243 ( .A(div_cnt[2]), .B(N77), .Z(N78) );
  GTECH_OR2 C244 ( .A(div_cnt[1]), .B(N78), .Z(N79) );
  GTECH_OR2 C245 ( .A(div_cnt[0]), .B(N79), .Z(N80) );
  GTECH_NOT I_20 ( .A(N80), .Z(N81) );
  GTECH_OR2 C247 ( .A(div_cnt[4]), .B(div_cnt[5]), .Z(N82) );
  GTECH_OR2 C248 ( .A(div_cnt[3]), .B(N82), .Z(N83) );
  GTECH_OR2 C249 ( .A(div_cnt[2]), .B(N83), .Z(N84) );
  GTECH_OR2 C250 ( .A(div_cnt[1]), .B(N84), .Z(N85) );
  GTECH_OR2 C251 ( .A(div_cnt[0]), .B(N85), .Z(N86) );
  GTECH_NOT I_21 ( .A(N86), .Z(N87) );
  GTECH_OR2 C253 ( .A(div_exp_out[10]), .B(div_exp_out[11]), .Z(N88) );
  GTECH_OR2 C254 ( .A(div_exp_out[9]), .B(N88), .Z(N89) );
  GTECH_OR2 C255 ( .A(div_exp_out[8]), .B(N89), .Z(N90) );
  GTECH_OR2 C256 ( .A(div_exp_out[7]), .B(N90), .Z(N91) );
  GTECH_OR2 C257 ( .A(div_exp_out[6]), .B(N91), .Z(N92) );
  GTECH_OR2 C258 ( .A(div_exp_out[5]), .B(N92), .Z(N93) );
  GTECH_OR2 C259 ( .A(div_exp_out[4]), .B(N93), .Z(N94) );
  GTECH_OR2 C260 ( .A(div_exp_out[3]), .B(N94), .Z(N95) );
  GTECH_OR2 C261 ( .A(div_exp_out[2]), .B(N95), .Z(N96) );
  GTECH_OR2 C262 ( .A(div_exp_out[1]), .B(N96), .Z(N97) );
  GTECH_NOT I_22 ( .A(div_rnd_mode[0]), .Z(N98) );
  GTECH_OR2 C266 ( .A(N98), .B(div_rnd_mode[1]), .Z(N99) );
  GTECH_NOT I_23 ( .A(N99), .Z(N100) );
  GTECH_NOT I_24 ( .A(div_rnd_mode[1]), .Z(N101) );
  GTECH_OR2 C269 ( .A(div_rnd_mode[0]), .B(N101), .Z(N102) );
  GTECH_NOT I_25 ( .A(N102), .Z(N103) );
  GTECH_AND2 C271 ( .A(div_rnd_mode[0]), .B(div_rnd_mode[1]), .Z(N104) );
  GTECH_OR2 C273 ( .A(div_rnd_mode[0]), .B(N101), .Z(N105) );
  GTECH_NOT I_26 ( .A(N105), .Z(N106) );
  GTECH_AND2 C275 ( .A(div_rnd_mode[0]), .B(div_rnd_mode[1]), .Z(N107) );
  GTECH_OR2 C276 ( .A(div_rnd_mode[0]), .B(div_rnd_mode[1]), .Z(N108) );
  GTECH_NOT I_27 ( .A(N108), .Z(N109) );
  GTECH_OR2 C282 ( .A(N11), .B(d1stg_op[7]), .Z(N110) );
  GTECH_OR2 C283 ( .A(d1stg_op[5]), .B(N110), .Z(N111) );
  GTECH_OR2 C284 ( .A(d1stg_op[4]), .B(N111), .Z(N112) );
  GTECH_OR2 C285 ( .A(N12), .B(N112), .Z(N113) );
  GTECH_OR2 C286 ( .A(N13), .B(N113), .Z(N114) );
  GTECH_OR2 C287 ( .A(d1stg_op[1]), .B(N114), .Z(N115) );
  GTECH_OR2 C288 ( .A(N14), .B(N115), .Z(N116) );
  GTECH_NOT I_28 ( .A(N116), .Z(N117) );
  GTECH_OR2 C294 ( .A(N11), .B(d1stg_op[7]), .Z(N118) );
  GTECH_OR2 C295 ( .A(d1stg_op[5]), .B(N118), .Z(N119) );
  GTECH_OR2 C296 ( .A(d1stg_op[4]), .B(N119), .Z(N120) );
  GTECH_OR2 C297 ( .A(N12), .B(N120), .Z(N121) );
  GTECH_OR2 C298 ( .A(N13), .B(N121), .Z(N122) );
  GTECH_OR2 C299 ( .A(N23), .B(N122), .Z(N123) );
  GTECH_OR2 C300 ( .A(d1stg_op[0]), .B(N123), .Z(N124) );
  GTECH_NOT I_29 ( .A(N124), .Z(N125) );
  GTECH_NOT I_30 ( .A(div_cnt[5]), .Z(N126) );
  GTECH_NOT I_31 ( .A(div_cnt[4]), .Z(N127) );
  GTECH_NOT I_32 ( .A(div_cnt[2]), .Z(N128) );
  GTECH_NOT I_33 ( .A(div_cnt[1]), .Z(N129) );
  GTECH_OR2 C306 ( .A(N127), .B(N126), .Z(N130) );
  GTECH_OR2 C307 ( .A(div_cnt[3]), .B(N130), .Z(N131) );
  GTECH_OR2 C308 ( .A(N128), .B(N131), .Z(N132) );
  GTECH_OR2 C309 ( .A(N129), .B(N132), .Z(N133) );
  GTECH_OR2 C310 ( .A(div_cnt[0]), .B(N133), .Z(N134) );
  GTECH_NOT I_34 ( .A(N134), .Z(N135) );
  GTECH_NOT I_35 ( .A(div_cnt[3]), .Z(N136) );
  GTECH_NOT I_36 ( .A(div_cnt[0]), .Z(N137) );
  GTECH_OR2 C315 ( .A(N127), .B(div_cnt[5]), .Z(N138) );
  GTECH_OR2 C316 ( .A(N136), .B(N138), .Z(N139) );
  GTECH_OR2 C317 ( .A(div_cnt[2]), .B(N139), .Z(N140) );
  GTECH_OR2 C318 ( .A(div_cnt[1]), .B(N140), .Z(N141) );
  GTECH_OR2 C319 ( .A(N137), .B(N141), .Z(N142) );
  GTECH_NOT I_37 ( .A(N142), .Z(N143) );
  GTECH_OR2 C321 ( .A(div_exp1[11]), .B(div_exp1[12]), .Z(N144) );
  GTECH_OR2 C322 ( .A(div_exp1[10]), .B(N144), .Z(N145) );
  GTECH_OR2 C323 ( .A(div_exp1[9]), .B(N145), .Z(N146) );
  GTECH_OR2 C324 ( .A(div_exp1[8]), .B(N146), .Z(N147) );
  GTECH_OR2 C325 ( .A(div_exp1[7]), .B(N147), .Z(N148) );
  GTECH_OR2 C326 ( .A(div_exp1[6]), .B(N148), .Z(N149) );
  GTECH_OR2 C327 ( .A(div_exp1[5]), .B(N149), .Z(N150) );
  GTECH_OR2 C328 ( .A(div_exp1[4]), .B(N150), .Z(N151) );
  GTECH_OR2 C329 ( .A(div_exp1[3]), .B(N151), .Z(N152) );
  GTECH_OR2 C330 ( .A(div_exp1[2]), .B(N152), .Z(N153) );
  GTECH_OR2 C331 ( .A(div_exp1[1]), .B(N153), .Z(N154) );
  GTECH_OR2 C332 ( .A(div_exp1[0]), .B(N154), .Z(N155) );
  GTECH_OR2 C335 ( .A(div_exp1[11]), .B(div_exp1[12]), .Z(N156) );
  GTECH_OR2 C336 ( .A(div_exp1[10]), .B(N156), .Z(N157) );
  GTECH_OR2 C337 ( .A(div_exp1[9]), .B(N157), .Z(N158) );
  GTECH_OR2 C338 ( .A(div_exp1[8]), .B(N158), .Z(N159) );
  GTECH_OR2 C339 ( .A(div_exp1[7]), .B(N159), .Z(N160) );
  GTECH_OR2 C340 ( .A(div_exp1[6]), .B(N160), .Z(N161) );
  GTECH_OR2 C341 ( .A(div_exp1[5]), .B(N161), .Z(N162) );
  GTECH_OR2 C342 ( .A(div_exp1[4]), .B(N162), .Z(N163) );
  GTECH_OR2 C343 ( .A(div_exp1[3]), .B(N163), .Z(N164) );
  GTECH_OR2 C344 ( .A(div_exp1[2]), .B(N164), .Z(N165) );
  GTECH_OR2 C345 ( .A(div_exp1[1]), .B(N165), .Z(N166) );
  GTECH_OR2 C346 ( .A(div_exp1[0]), .B(N166), .Z(N167) );
  GTECH_NOT I_38 ( .A(N167), .Z(N168) );
  ADD_UNS_OP add_1554 ( .A(div_cnt), .B(1'b1), .Z(div_cnt_plus1) );
  GTECH_NOT I_39 ( .A(div_ctl_rst_l), .Z(reset) );
  GTECH_AND2 C351 ( .A(div_exp_in1_exp_eq_0), .B(d1stg_sngopa[0]), .Z(
        d1stg_denorm_sng_in1) );
  GTECH_AND2 C352 ( .A(div_exp_in1_exp_eq_0), .B(d1stg_dblopa[0]), .Z(
        d1stg_denorm_dbl_in1) );
  GTECH_AND2 C353 ( .A(div_exp_in2_exp_eq_0), .B(d1stg_sngopa[0]), .Z(
        d1stg_denorm_sng_in2) );
  GTECH_AND2 C354 ( .A(div_exp_in2_exp_eq_0), .B(d1stg_dblopa[0]), .Z(
        d1stg_denorm_dbl_in2) );
  GTECH_AND2 C355 ( .A(N169), .B(d1stg_sngopa[0]), .Z(d1stg_norm_sng_in1) );
  GTECH_NOT I_40 ( .A(div_exp_in1_exp_eq_0), .Z(N169) );
  GTECH_AND2 C357 ( .A(N169), .B(d1stg_dblopa[0]), .Z(d1stg_norm_dbl_in1) );
  GTECH_AND2 C359 ( .A(N170), .B(d1stg_sngopa[0]), .Z(d1stg_norm_sng_in2) );
  GTECH_NOT I_41 ( .A(div_exp_in2_exp_eq_0), .Z(N170) );
  GTECH_AND2 C361 ( .A(N170), .B(d1stg_dblopa[0]), .Z(d1stg_norm_dbl_in2) );
  GTECH_AND2 C363 ( .A(N174), .B(d1stg_sngopa[1]), .Z(d1stg_snan_sng_in1) );
  GTECH_AND2 C364 ( .A(N173), .B(div_frac_in1_53_32_neq_0), .Z(N174) );
  GTECH_AND2 C365 ( .A(N171), .B(N172), .Z(N173) );
  GTECH_NOT I_42 ( .A(div_exp_in1_exp_neq_ffs), .Z(N171) );
  GTECH_NOT I_43 ( .A(div_frac_in1_54), .Z(N172) );
  GTECH_AND2 C368 ( .A(N177), .B(d1stg_dblopa[1]), .Z(d1stg_snan_dbl_in1) );
  GTECH_AND2 C369 ( .A(N176), .B(div_frac_in1_50_0_neq_0), .Z(N177) );
  GTECH_AND2 C370 ( .A(N171), .B(N175), .Z(N176) );
  GTECH_NOT I_44 ( .A(div_frac_in1_51), .Z(N175) );
  GTECH_AND2 C373 ( .A(N181), .B(d1stg_sngopa[1]), .Z(d1stg_snan_sng_in2) );
  GTECH_AND2 C374 ( .A(N180), .B(div_frac_in2_53_32_neq_0), .Z(N181) );
  GTECH_AND2 C375 ( .A(N178), .B(N179), .Z(N180) );
  GTECH_NOT I_45 ( .A(div_exp_in2_exp_neq_ffs), .Z(N178) );
  GTECH_NOT I_46 ( .A(div_frac_in2_54), .Z(N179) );
  GTECH_AND2 C378 ( .A(N184), .B(d1stg_dblopa[1]), .Z(d1stg_snan_dbl_in2) );
  GTECH_AND2 C379 ( .A(N183), .B(div_frac_in2_50_0_neq_0), .Z(N184) );
  GTECH_AND2 C380 ( .A(N178), .B(N182), .Z(N183) );
  GTECH_NOT I_47 ( .A(div_frac_in2_51), .Z(N182) );
  GTECH_AND2 C383 ( .A(N185), .B(d1stg_sngopa[1]), .Z(d1stg_qnan_sng_in1) );
  GTECH_AND2 C384 ( .A(N171), .B(div_frac_in1_54), .Z(N185) );
  GTECH_AND2 C386 ( .A(N186), .B(d1stg_dblopa[1]), .Z(d1stg_qnan_dbl_in1) );
  GTECH_AND2 C387 ( .A(N171), .B(div_frac_in1_51), .Z(N186) );
  GTECH_AND2 C389 ( .A(N187), .B(d1stg_sngopa[1]), .Z(d1stg_qnan_sng_in2) );
  GTECH_AND2 C390 ( .A(N178), .B(div_frac_in2_54), .Z(N187) );
  GTECH_AND2 C392 ( .A(N188), .B(d1stg_dblopa[1]), .Z(d1stg_qnan_dbl_in2) );
  GTECH_AND2 C393 ( .A(N178), .B(div_frac_in2_51), .Z(N188) );
  GTECH_OR2 C395 ( .A(d1stg_snan_sng_in1), .B(d1stg_snan_dbl_in1), .Z(
        d1stg_snan_in1) );
  GTECH_OR2 C396 ( .A(d1stg_snan_sng_in2), .B(d1stg_snan_dbl_in2), .Z(
        d1stg_snan_in2) );
  GTECH_OR2 C397 ( .A(d1stg_qnan_sng_in1), .B(d1stg_qnan_dbl_in1), .Z(
        d1stg_qnan_in1) );
  GTECH_OR2 C398 ( .A(d1stg_qnan_sng_in2), .B(d1stg_qnan_dbl_in2), .Z(
        d1stg_qnan_in2) );
  GTECH_AND2 C399 ( .A(N190), .B(d1stg_sngopa[2]), .Z(d1stg_nan_sng_in1) );
  GTECH_AND2 C400 ( .A(N171), .B(N189), .Z(N190) );
  GTECH_OR2 C402 ( .A(div_frac_in1_54), .B(div_frac_in1_53_32_neq_0), .Z(N189)
         );
  GTECH_AND2 C403 ( .A(N192), .B(d1stg_dblopa[2]), .Z(d1stg_nan_dbl_in1) );
  GTECH_AND2 C404 ( .A(N171), .B(N191), .Z(N192) );
  GTECH_OR2 C406 ( .A(div_frac_in1_51), .B(div_frac_in1_50_0_neq_0), .Z(N191)
         );
  GTECH_AND2 C407 ( .A(N194), .B(d1stg_sngopa[2]), .Z(d1stg_nan_sng_in2) );
  GTECH_AND2 C408 ( .A(N178), .B(N193), .Z(N194) );
  GTECH_OR2 C410 ( .A(div_frac_in2_54), .B(div_frac_in2_53_32_neq_0), .Z(N193)
         );
  GTECH_AND2 C411 ( .A(N196), .B(d1stg_dblopa[2]), .Z(d1stg_nan_dbl_in2) );
  GTECH_AND2 C412 ( .A(N178), .B(N195), .Z(N196) );
  GTECH_OR2 C414 ( .A(div_frac_in2_51), .B(div_frac_in2_50_0_neq_0), .Z(N195)
         );
  GTECH_OR2 C415 ( .A(d1stg_nan_sng_in1), .B(d1stg_nan_dbl_in1), .Z(
        d1stg_nan_in1) );
  GTECH_OR2 C416 ( .A(d1stg_nan_sng_in2), .B(d1stg_nan_dbl_in2), .Z(
        d1stg_nan_in2) );
  GTECH_OR2 C417 ( .A(d1stg_nan_in1), .B(d1stg_nan_in2), .Z(d1stg_nan_in) );
  GTECH_AND2 C418 ( .A(N199), .B(d1stg_sngopa[2]), .Z(d1stg_inf_sng_in1) );
  GTECH_AND2 C419 ( .A(N197), .B(N198), .Z(N199) );
  GTECH_AND2 C420 ( .A(N171), .B(N172), .Z(N197) );
  GTECH_NOT I_48 ( .A(div_frac_in1_53_32_neq_0), .Z(N198) );
  GTECH_AND2 C424 ( .A(N202), .B(d1stg_dblopa[2]), .Z(d1stg_inf_dbl_in1) );
  GTECH_AND2 C425 ( .A(N200), .B(N201), .Z(N202) );
  GTECH_AND2 C426 ( .A(N171), .B(N175), .Z(N200) );
  GTECH_NOT I_49 ( .A(div_frac_in1_50_0_neq_0), .Z(N201) );
  GTECH_AND2 C430 ( .A(N205), .B(d1stg_sngopa[2]), .Z(d1stg_inf_sng_in2) );
  GTECH_AND2 C431 ( .A(N203), .B(N204), .Z(N205) );
  GTECH_AND2 C432 ( .A(N178), .B(N179), .Z(N203) );
  GTECH_NOT I_50 ( .A(div_frac_in2_53_32_neq_0), .Z(N204) );
  GTECH_AND2 C436 ( .A(N208), .B(d1stg_dblopa[2]), .Z(d1stg_inf_dbl_in2) );
  GTECH_AND2 C437 ( .A(N206), .B(N207), .Z(N208) );
  GTECH_AND2 C438 ( .A(N178), .B(N182), .Z(N206) );
  GTECH_NOT I_51 ( .A(div_frac_in2_50_0_neq_0), .Z(N207) );
  GTECH_OR2 C442 ( .A(d1stg_inf_sng_in1), .B(d1stg_inf_dbl_in1), .Z(
        d1stg_inf_in1) );
  GTECH_OR2 C443 ( .A(d1stg_inf_sng_in2), .B(d1stg_inf_dbl_in2), .Z(
        d1stg_inf_in2) );
  GTECH_OR2 C444 ( .A(d1stg_inf_in1), .B(d1stg_inf_in2), .Z(d1stg_inf_in) );
  GTECH_AND2 C445 ( .A(d1stg_inf_in1), .B(d1stg_inf_in2), .Z(d1stg_2inf_in) );
  GTECH_AND2 C446 ( .A(N171), .B(d1stg_sngopa[3]), .Z(d1stg_infnan_sng_in1) );
  GTECH_AND2 C448 ( .A(N171), .B(d1stg_dblopa[3]), .Z(d1stg_infnan_dbl_in1) );
  GTECH_AND2 C450 ( .A(N178), .B(d1stg_sngopa[3]), .Z(d1stg_infnan_sng_in2) );
  GTECH_AND2 C452 ( .A(N178), .B(d1stg_dblopa[3]), .Z(d1stg_infnan_dbl_in2) );
  GTECH_OR2 C454 ( .A(d1stg_infnan_sng_in1), .B(d1stg_infnan_dbl_in1), .Z(
        d1stg_infnan_in1) );
  GTECH_OR2 C455 ( .A(d1stg_infnan_sng_in2), .B(d1stg_infnan_dbl_in2), .Z(
        d1stg_infnan_in2) );
  GTECH_OR2 C456 ( .A(d1stg_infnan_in1), .B(d1stg_infnan_in2), .Z(
        d1stg_infnan_in) );
  GTECH_AND2 C457 ( .A(N210), .B(N172), .Z(d1stg_zero_in1) );
  GTECH_AND2 C458 ( .A(div_exp_in1_exp_eq_0), .B(N209), .Z(N210) );
  GTECH_NOT I_52 ( .A(div_frac_in1_53_0_neq_0), .Z(N209) );
  GTECH_AND2 C461 ( .A(N212), .B(N179), .Z(d1stg_zero_in2) );
  GTECH_AND2 C462 ( .A(div_exp_in2_exp_eq_0), .B(N211), .Z(N212) );
  GTECH_NOT I_53 ( .A(div_frac_in2_53_0_neq_0), .Z(N211) );
  GTECH_OR2 C465 ( .A(d1stg_zero_in1), .B(d1stg_zero_in2), .Z(d1stg_zero_in)
         );
  GTECH_AND2 C466 ( .A(d1stg_zero_in1), .B(d1stg_zero_in2), .Z(d1stg_2zero_in)
         );
  GTECH_OR2 C467 ( .A(N214), .B(divd_cnt_lt_52), .Z(d1stg_hold) );
  GTECH_OR2 C468 ( .A(N213), .B(divs_cnt_lt_23), .Z(N214) );
  GTECH_OR2 C469 ( .A(d1stg_div), .B(d234stg_fdiv), .Z(N213) );
  GTECH_OR2 C470 ( .A(N216), .B(divd_cnt_lt_52a), .Z(d1stg_holda) );
  GTECH_OR2 C471 ( .A(N215), .B(divs_cnt_lt_23a), .Z(N216) );
  GTECH_OR2 C472 ( .A(d1stg_div), .B(d234stg_fdiv), .Z(N215) );
  GTECH_NOT I_54 ( .A(d1stg_hold), .Z(d1stg_step) );
  GTECH_NOT I_55 ( .A(d1stg_holda), .Z(d1stg_stepa) );
  GTECH_AND2 C475 ( .A(d1stg_stepa), .B(N217), .Z(d1stg_op_in[7]) );
  GTECH_AND2 C476 ( .A(inq_op[7]), .B(inq_div), .Z(N217) );
  GTECH_AND2 C477 ( .A(d1stg_stepa), .B(N218), .Z(d1stg_op_in[6]) );
  GTECH_AND2 C478 ( .A(inq_op[6]), .B(inq_div), .Z(N218) );
  GTECH_AND2 C479 ( .A(d1stg_stepa), .B(N219), .Z(d1stg_op_in[5]) );
  GTECH_AND2 C480 ( .A(inq_op[5]), .B(inq_div), .Z(N219) );
  GTECH_AND2 C481 ( .A(d1stg_stepa), .B(N220), .Z(d1stg_op_in[4]) );
  GTECH_AND2 C482 ( .A(inq_op[4]), .B(inq_div), .Z(N220) );
  GTECH_AND2 C483 ( .A(d1stg_stepa), .B(N221), .Z(d1stg_op_in[3]) );
  GTECH_AND2 C484 ( .A(inq_op[3]), .B(inq_div), .Z(N221) );
  GTECH_AND2 C485 ( .A(d1stg_stepa), .B(N222), .Z(d1stg_op_in[2]) );
  GTECH_AND2 C486 ( .A(inq_op[2]), .B(inq_div), .Z(N222) );
  GTECH_AND2 C487 ( .A(d1stg_stepa), .B(N223), .Z(d1stg_op_in[1]) );
  GTECH_AND2 C488 ( .A(inq_op[1]), .B(inq_div), .Z(N223) );
  GTECH_AND2 C489 ( .A(d1stg_stepa), .B(N224), .Z(d1stg_op_in[0]) );
  GTECH_AND2 C490 ( .A(inq_op[0]), .B(inq_div), .Z(N224) );
  GTECH_AND2 C491 ( .A(inq_div), .B(d1stg_stepa), .Z(d1stg_div_in) );
  GTECH_OR2 C492 ( .A(N117), .B(N125), .Z(d1stg_opdec[2]) );
  GTECH_OR2 C493 ( .A(N225), .B(d3stg_fdiv), .Z(d234stg_fdiv_in) );
  GTECH_OR2 C494 ( .A(d1stg_opdec[2]), .B(d2stg_opdec[2]), .Z(N225) );
  GTECH_OR2 C495 ( .A(N226), .B(d6stg_step), .Z(d5stg_step) );
  GTECH_NOT I_56 ( .A(d5stg_opdec[2]), .Z(N226) );
  GTECH_AND2 C497 ( .A(N230), .B(N231), .Z(d5stg_fdivb_in) );
  GTECH_OR2 C498 ( .A(N227), .B(N229), .Z(N230) );
  GTECH_AND2 C499 ( .A(d5stg_step), .B(d4stg_fdiv), .Z(N227) );
  GTECH_AND2 C500 ( .A(N228), .B(d5stg_opdec[2]), .Z(N229) );
  GTECH_NOT I_57 ( .A(d5stg_step), .Z(N228) );
  GTECH_NOT I_58 ( .A(reset), .Z(N231) );
  GTECH_OR2 C503 ( .A(N234), .B(N241), .Z(d6stg_step) );
  GTECH_OR2 C504 ( .A(N232), .B(N233), .Z(N234) );
  GTECH_AND2 C505 ( .A(d5stg_fdivd), .B(N135), .Z(N232) );
  GTECH_AND2 C506 ( .A(d5stg_fdivs), .B(N143), .Z(N233) );
  GTECH_AND2 C507 ( .A(d5stg_opdec[2]), .B(N240), .Z(N241) );
  GTECH_OR2 C508 ( .A(N238), .B(N239), .Z(N240) );
  GTECH_OR2 C509 ( .A(N235), .B(N237), .Z(N238) );
  GTECH_AND2 C510 ( .A(N0), .B(N155), .Z(N235) );
  GTECH_AND2 C511 ( .A(N236), .B(d8stg_step), .Z(N237) );
  GTECH_AND2 C512 ( .A(N1), .B(N168), .Z(N236) );
  GTECH_AND2 C513 ( .A(div_exp1[12]), .B(d8stg_step), .Z(N239) );
  GTECH_AND2 C514 ( .A(d6stg_step), .B(d5stg_opdec[2]), .Z(d6stg_opdec_in[2])
         );
  GTECH_AND2 C515 ( .A(d6stg_step), .B(d5stg_fdivs), .Z(d6stg_opdec_in[1]) );
  GTECH_AND2 C516 ( .A(d6stg_step), .B(d5stg_fdivd), .Z(d6stg_opdec_in[0]) );
  GTECH_NOT I_59 ( .A(reset), .Z(N2) );
  GTECH_OR2 C518 ( .A(N243), .B(N246), .Z(d8stg_fdiv_in) );
  GTECH_AND2 C519 ( .A(N242), .B(d7stg_fdiv), .Z(N243) );
  GTECH_AND2 C520 ( .A(d8stg_step), .B(N2), .Z(N242) );
  GTECH_AND2 C521 ( .A(N245), .B(d8stg_opdec[2]), .Z(N246) );
  GTECH_AND2 C522 ( .A(N244), .B(N2), .Z(N245) );
  GTECH_NOT I_60 ( .A(d8stg_step), .Z(N244) );
  GTECH_AND2 C524 ( .A(d8stg_opdec[2]), .B(N247), .Z(d8stg_hold) );
  GTECH_NOT I_61 ( .A(div_dest_rdy), .Z(N247) );
  GTECH_NOT I_62 ( .A(d8stg_hold), .Z(d8stg_step) );
  GTECH_OR2 C527 ( .A(N253), .B(d8stg_opdec[2]), .Z(div_pipe_active_in) );
  GTECH_OR2 C528 ( .A(N252), .B(d7stg_fdiv), .Z(N253) );
  GTECH_OR2 C529 ( .A(N251), .B(d6stg_fdiv), .Z(N252) );
  GTECH_OR2 C530 ( .A(N249), .B(N250), .Z(N251) );
  GTECH_OR2 C531 ( .A(N248), .B(d3stg_fdiv), .Z(N249) );
  GTECH_OR2 C532 ( .A(d1stg_opdec[2]), .B(d2stg_opdec[2]), .Z(N248) );
  GTECH_OR2 C533 ( .A(d4stg_fdiv), .B(d5stg_opdec[2]), .Z(N250) );
  GTECH_NOT I_63 ( .A(d2stg_snan_in2), .Z(N3) );
  GTECH_AND2 C535 ( .A(N266), .B(N268), .Z(d1stg_sign) );
  GTECH_XOR2 C536 ( .A(N258), .B(N265), .Z(N266) );
  GTECH_AND2 C537 ( .A(N254), .B(N257), .Z(N258) );
  GTECH_AND2 C538 ( .A(d1stg_sign1), .B(N3), .Z(N254) );
  GTECH_NOT I_64 ( .A(N256), .Z(N257) );
  GTECH_AND2 C540 ( .A(d2stg_qnan_in2), .B(N255), .Z(N256) );
  GTECH_NOT I_65 ( .A(d2stg_snan_in1), .Z(N255) );
  GTECH_AND2 C542 ( .A(N261), .B(N264), .Z(N265) );
  GTECH_AND2 C543 ( .A(d1stg_sign2), .B(N260), .Z(N261) );
  GTECH_NOT I_66 ( .A(N259), .Z(N260) );
  GTECH_AND2 C545 ( .A(d2stg_snan_in1), .B(N3), .Z(N259) );
  GTECH_NOT I_67 ( .A(N263), .Z(N264) );
  GTECH_AND2 C547 ( .A(d2stg_qnan_in1), .B(N262), .Z(N263) );
  GTECH_NOT I_68 ( .A(d2stg_nan_in2), .Z(N262) );
  GTECH_NOT I_69 ( .A(N267), .Z(N268) );
  GTECH_OR2 C550 ( .A(d2stg_2inf_in), .B(d2stg_2zero_in), .Z(N267) );
  GTECH_AND2 C551 ( .A(N269), .B(d8stg_step), .Z(div_bkend_step) );
  GTECH_AND2 C552 ( .A(d5stg_opdec[2]), .B(N87), .Z(N269) );
  GTECH_OR2 C553 ( .A(N270), .B(N272), .Z(div_id_out_in[9]) );
  GTECH_AND2 C554 ( .A(div_bkend_step), .B(N33), .Z(N270) );
  GTECH_AND2 C555 ( .A(N271), .B(div_id_out[9]), .Z(N272) );
  GTECH_NOT I_70 ( .A(div_bkend_step), .Z(N271) );
  GTECH_OR2 C557 ( .A(N273), .B(N275), .Z(div_id_out_in[8]) );
  GTECH_AND2 C558 ( .A(div_bkend_step), .B(N38), .Z(N273) );
  GTECH_AND2 C559 ( .A(N274), .B(div_id_out[8]), .Z(N275) );
  GTECH_NOT I_71 ( .A(div_bkend_step), .Z(N274) );
  GTECH_OR2 C561 ( .A(N276), .B(N278), .Z(div_id_out_in[7]) );
  GTECH_AND2 C562 ( .A(div_bkend_step), .B(N42), .Z(N276) );
  GTECH_AND2 C563 ( .A(N277), .B(div_id_out[7]), .Z(N278) );
  GTECH_NOT I_72 ( .A(div_bkend_step), .Z(N277) );
  GTECH_OR2 C565 ( .A(N279), .B(N281), .Z(div_id_out_in[6]) );
  GTECH_AND2 C566 ( .A(div_bkend_step), .B(N45), .Z(N279) );
  GTECH_AND2 C567 ( .A(N280), .B(div_id_out[6]), .Z(N281) );
  GTECH_NOT I_73 ( .A(div_bkend_step), .Z(N280) );
  GTECH_OR2 C569 ( .A(N282), .B(N284), .Z(div_id_out_in[5]) );
  GTECH_AND2 C570 ( .A(div_bkend_step), .B(N48), .Z(N282) );
  GTECH_AND2 C571 ( .A(N283), .B(div_id_out[5]), .Z(N284) );
  GTECH_NOT I_74 ( .A(div_bkend_step), .Z(N283) );
  GTECH_OR2 C573 ( .A(N285), .B(N287), .Z(div_id_out_in[4]) );
  GTECH_AND2 C574 ( .A(div_bkend_step), .B(N51), .Z(N285) );
  GTECH_AND2 C575 ( .A(N286), .B(div_id_out[4]), .Z(N287) );
  GTECH_NOT I_75 ( .A(div_bkend_step), .Z(N286) );
  GTECH_OR2 C577 ( .A(N288), .B(N290), .Z(div_id_out_in[3]) );
  GTECH_AND2 C578 ( .A(div_bkend_step), .B(N54), .Z(N288) );
  GTECH_AND2 C579 ( .A(N289), .B(div_id_out[3]), .Z(N290) );
  GTECH_NOT I_76 ( .A(div_bkend_step), .Z(N289) );
  GTECH_OR2 C581 ( .A(N291), .B(N293), .Z(div_id_out_in[2]) );
  GTECH_AND2 C582 ( .A(div_bkend_step), .B(N57), .Z(N291) );
  GTECH_AND2 C583 ( .A(N292), .B(div_id_out[2]), .Z(N293) );
  GTECH_NOT I_77 ( .A(div_bkend_step), .Z(N292) );
  GTECH_OR2 C585 ( .A(N294), .B(N296), .Z(div_id_out_in[1]) );
  GTECH_AND2 C586 ( .A(div_bkend_step), .B(d1stg_id[1]), .Z(N294) );
  GTECH_AND2 C587 ( .A(N295), .B(div_id_out[1]), .Z(N296) );
  GTECH_NOT I_78 ( .A(div_bkend_step), .Z(N295) );
  GTECH_OR2 C589 ( .A(N297), .B(N299), .Z(div_id_out_in[0]) );
  GTECH_AND2 C590 ( .A(div_bkend_step), .B(d1stg_id[0]), .Z(N297) );
  GTECH_AND2 C591 ( .A(N298), .B(div_id_out[0]), .Z(N299) );
  GTECH_NOT I_79 ( .A(div_bkend_step), .Z(N298) );
  GTECH_AND2 C593 ( .A(N300), .B(div_cnt_plus1[5]), .Z(div_cnt_in[5]) );
  GTECH_AND2 C594 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N300) );
  GTECH_AND2 C595 ( .A(N301), .B(div_cnt_plus1[4]), .Z(div_cnt_in[4]) );
  GTECH_AND2 C596 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N301) );
  GTECH_AND2 C597 ( .A(N302), .B(div_cnt_plus1[3]), .Z(div_cnt_in[3]) );
  GTECH_AND2 C598 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N302) );
  GTECH_AND2 C599 ( .A(N303), .B(div_cnt_plus1[2]), .Z(div_cnt_in[2]) );
  GTECH_AND2 C600 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N303) );
  GTECH_AND2 C601 ( .A(N304), .B(div_cnt_plus1[1]), .Z(div_cnt_in[1]) );
  GTECH_AND2 C602 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N304) );
  GTECH_AND2 C603 ( .A(N305), .B(div_cnt_plus1[0]), .Z(div_cnt_in[0]) );
  GTECH_AND2 C604 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N305) );
  GTECH_OR2 C605 ( .A(N306), .B(d4stg_fdiv), .Z(div_cnt_step) );
  GTECH_AND2 C606 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(N306) );
  GTECH_OR2 C607 ( .A(N307), .B(d8stg_step), .Z(div_cnt_lt_step) );
  GTECH_OR2 C608 ( .A(N226), .B(d6stg_step), .Z(N307) );
  GTECH_OR2 C610 ( .A(d4stg_opdec[1]), .B(N310), .Z(divs_cnt_lt_23_in) );
  GTECH_AND2 C611 ( .A(N309), .B(N4), .Z(N310) );
  GTECH_AND2 C612 ( .A(d5stg_fdivs), .B(N308), .Z(N309) );
  GTECH_NOT I_80 ( .A(d6stg_step), .Z(N308) );
  GTECH_OR2 C614 ( .A(d4stg_opdec[0]), .B(N312), .Z(divd_cnt_lt_52_in) );
  GTECH_AND2 C615 ( .A(N311), .B(N5), .Z(N312) );
  GTECH_AND2 C616 ( .A(d5stg_fdivd), .B(N308), .Z(N311) );
  GTECH_AND2 C618 ( .A(N313), .B(d8stg_step), .Z(div_exc_step) );
  GTECH_AND2 C619 ( .A(d5stg_opdec[2]), .B(N81), .Z(N313) );
  GTECH_NOT I_81 ( .A(N314), .Z(div_of_mask_in) );
  GTECH_OR2 C621 ( .A(d1stg_infnan_in), .B(d1stg_zero_in), .Z(N314) );
  GTECH_OR2 C622 ( .A(N316), .B(d1stg_2zero_in), .Z(div_nv_out_in) );
  GTECH_OR2 C623 ( .A(N315), .B(d1stg_2inf_in), .Z(N316) );
  GTECH_OR2 C624 ( .A(d1stg_snan_in1), .B(d1stg_snan_in2), .Z(N315) );
  GTECH_AND2 C625 ( .A(N318), .B(N319), .Z(div_dz_out_in) );
  GTECH_AND2 C626 ( .A(d1stg_zero_in2), .B(N317), .Z(N318) );
  GTECH_NOT I_82 ( .A(d1stg_zero_in1), .Z(N317) );
  GTECH_NOT I_83 ( .A(d1stg_infnan_in1), .Z(N319) );
  GTECH_NOT I_84 ( .A(div_exp_out[12]), .Z(N6) );
  GTECH_OR2 C630 ( .A(N333), .B(N347), .Z(d7stg_in_of) );
  GTECH_AND2 C631 ( .A(N332), .B(div_of_mask), .Z(N333) );
  GTECH_AND2 C632 ( .A(N320), .B(N331), .Z(N332) );
  GTECH_AND2 C633 ( .A(N6), .B(d7stg_fdivd), .Z(N320) );
  GTECH_OR2 C634 ( .A(div_exp_out[11]), .B(N330), .Z(N331) );
  GTECH_AND2 C635 ( .A(N329), .B(div_exp_out[0]), .Z(N330) );
  GTECH_AND2 C636 ( .A(N328), .B(div_exp_out[1]), .Z(N329) );
  GTECH_AND2 C637 ( .A(N327), .B(div_exp_out[2]), .Z(N328) );
  GTECH_AND2 C638 ( .A(N326), .B(div_exp_out[3]), .Z(N327) );
  GTECH_AND2 C639 ( .A(N325), .B(div_exp_out[4]), .Z(N326) );
  GTECH_AND2 C640 ( .A(N324), .B(div_exp_out[5]), .Z(N325) );
  GTECH_AND2 C641 ( .A(N323), .B(div_exp_out[6]), .Z(N324) );
  GTECH_AND2 C642 ( .A(N322), .B(div_exp_out[7]), .Z(N323) );
  GTECH_AND2 C643 ( .A(N321), .B(div_exp_out[8]), .Z(N322) );
  GTECH_AND2 C644 ( .A(div_exp_out[10]), .B(div_exp_out[9]), .Z(N321) );
  GTECH_AND2 C645 ( .A(N346), .B(div_of_mask), .Z(N347) );
  GTECH_AND2 C646 ( .A(N334), .B(N345), .Z(N346) );
  GTECH_AND2 C647 ( .A(N6), .B(d7stg_opdec[1]), .Z(N334) );
  GTECH_OR2 C648 ( .A(N337), .B(N344), .Z(N345) );
  GTECH_OR2 C649 ( .A(N336), .B(div_exp_out[8]), .Z(N337) );
  GTECH_OR2 C650 ( .A(N335), .B(div_exp_out[9]), .Z(N336) );
  GTECH_OR2 C651 ( .A(div_exp_out[11]), .B(div_exp_out[10]), .Z(N335) );
  GTECH_AND2 C652 ( .A(N343), .B(div_exp_out[0]), .Z(N344) );
  GTECH_AND2 C653 ( .A(N342), .B(div_exp_out[1]), .Z(N343) );
  GTECH_AND2 C654 ( .A(N341), .B(div_exp_out[2]), .Z(N342) );
  GTECH_AND2 C655 ( .A(N340), .B(div_exp_out[3]), .Z(N341) );
  GTECH_AND2 C656 ( .A(N339), .B(div_exp_out[4]), .Z(N340) );
  GTECH_AND2 C657 ( .A(N338), .B(div_exp_out[5]), .Z(N339) );
  GTECH_AND2 C658 ( .A(div_exp_out[7]), .B(div_exp_out[6]), .Z(N338) );
  GTECH_OR2 C659 ( .A(N360), .B(N370), .Z(div_of_out_tmp1_in) );
  GTECH_AND2 C660 ( .A(N359), .B(div_of_mask), .Z(N360) );
  GTECH_AND2 C661 ( .A(N358), .B(d7stg_rndup), .Z(N359) );
  GTECH_AND2 C662 ( .A(N348), .B(N357), .Z(N358) );
  GTECH_AND2 C663 ( .A(N6), .B(d7stg_fdivd), .Z(N348) );
  GTECH_AND2 C664 ( .A(N356), .B(div_exp_out[1]), .Z(N357) );
  GTECH_AND2 C665 ( .A(N355), .B(div_exp_out[2]), .Z(N356) );
  GTECH_AND2 C666 ( .A(N354), .B(div_exp_out[3]), .Z(N355) );
  GTECH_AND2 C667 ( .A(N353), .B(div_exp_out[4]), .Z(N354) );
  GTECH_AND2 C668 ( .A(N352), .B(div_exp_out[5]), .Z(N353) );
  GTECH_AND2 C669 ( .A(N351), .B(div_exp_out[6]), .Z(N352) );
  GTECH_AND2 C670 ( .A(N350), .B(div_exp_out[7]), .Z(N351) );
  GTECH_AND2 C671 ( .A(N349), .B(div_exp_out[8]), .Z(N350) );
  GTECH_AND2 C672 ( .A(div_exp_out[10]), .B(div_exp_out[9]), .Z(N349) );
  GTECH_AND2 C673 ( .A(N369), .B(div_of_mask), .Z(N370) );
  GTECH_AND2 C674 ( .A(N368), .B(d7stg_rndup), .Z(N369) );
  GTECH_AND2 C675 ( .A(N361), .B(N367), .Z(N368) );
  GTECH_AND2 C676 ( .A(N6), .B(d7stg_opdec[1]), .Z(N361) );
  GTECH_AND2 C677 ( .A(N366), .B(div_exp_out[1]), .Z(N367) );
  GTECH_AND2 C678 ( .A(N365), .B(div_exp_out[2]), .Z(N366) );
  GTECH_AND2 C679 ( .A(N364), .B(div_exp_out[3]), .Z(N365) );
  GTECH_AND2 C680 ( .A(N363), .B(div_exp_out[4]), .Z(N364) );
  GTECH_AND2 C681 ( .A(N362), .B(div_exp_out[5]), .Z(N363) );
  GTECH_AND2 C682 ( .A(div_exp_out[7]), .B(div_exp_out[6]), .Z(N362) );
  GTECH_OR2 C683 ( .A(div_of_out_tmp2), .B(N372), .Z(div_exc_out[3]) );
  GTECH_AND2 C684 ( .A(div_of_out_tmp1), .B(N371), .Z(N372) );
  GTECH_NOT I_85 ( .A(div_out_52_inv), .Z(N371) );
  GTECH_OR2 C686 ( .A(N388), .B(N389), .Z(div_uf_out_in) );
  GTECH_AND2 C687 ( .A(N387), .B(div_of_mask), .Z(N388) );
  GTECH_AND2 C688 ( .A(N384), .B(N386), .Z(N387) );
  GTECH_NOT I_86 ( .A(N383), .Z(N384) );
  GTECH_OR2 C690 ( .A(N382), .B(div_exp_out[0]), .Z(N383) );
  GTECH_OR2 C691 ( .A(N381), .B(div_exp_out[1]), .Z(N382) );
  GTECH_OR2 C692 ( .A(N380), .B(div_exp_out[2]), .Z(N381) );
  GTECH_OR2 C693 ( .A(N379), .B(div_exp_out[3]), .Z(N380) );
  GTECH_OR2 C694 ( .A(N378), .B(div_exp_out[4]), .Z(N379) );
  GTECH_OR2 C695 ( .A(N377), .B(div_exp_out[5]), .Z(N378) );
  GTECH_OR2 C696 ( .A(N376), .B(div_exp_out[6]), .Z(N377) );
  GTECH_OR2 C697 ( .A(N375), .B(div_exp_out[7]), .Z(N376) );
  GTECH_OR2 C698 ( .A(N374), .B(div_exp_out[8]), .Z(N375) );
  GTECH_OR2 C699 ( .A(N373), .B(div_exp_out[9]), .Z(N374) );
  GTECH_OR2 C700 ( .A(div_exp_out[11]), .B(div_exp_out[10]), .Z(N373) );
  GTECH_OR2 C701 ( .A(N385), .B(d7stg_stk), .Z(N386) );
  GTECH_OR2 C702 ( .A(div_frac_add_in1_neq_0), .B(d7stg_grd), .Z(N385) );
  GTECH_AND2 C703 ( .A(div_exp_out[12]), .B(div_of_mask), .Z(N389) );
  GTECH_OR2 C704 ( .A(d7stg_grd), .B(d7stg_stk), .Z(div_nx_out_in) );
  GTECH_OR2 C705 ( .A(div_nx_out), .B(div_exc_out[3]), .Z(div_exc_out[0]) );
  GTECH_AND2 C706 ( .A(N390), .B(N391), .Z(d1stg_spc_rslt) );
  GTECH_OR2 C707 ( .A(d1stg_inf_in), .B(d1stg_zero_in), .Z(N390) );
  GTECH_NOT I_87 ( .A(d1stg_nan_in), .Z(N391) );
  GTECH_AND2 C709 ( .A(N397), .B(N398), .Z(div_norm_frac_in1_dbl_norm) );
  GTECH_AND2 C710 ( .A(N394), .B(N396), .Z(N397) );
  GTECH_AND2 C711 ( .A(N392), .B(N393), .Z(N394) );
  GTECH_AND2 C712 ( .A(d1stg_opdec[2]), .B(d1stg_norm_dbl_in1), .Z(N392) );
  GTECH_NOT I_88 ( .A(d1stg_snan_dbl_in2), .Z(N393) );
  GTECH_OR2 C714 ( .A(N395), .B(d1stg_snan_dbl_in1), .Z(N396) );
  GTECH_NOT I_89 ( .A(d1stg_qnan_dbl_in2), .Z(N395) );
  GTECH_NOT I_90 ( .A(d1stg_spc_rslt), .Z(N398) );
  GTECH_AND2 C717 ( .A(N401), .B(N398), .Z(div_norm_frac_in1_dbl_dnrm) );
  GTECH_AND2 C718 ( .A(N400), .B(N395), .Z(N401) );
  GTECH_AND2 C719 ( .A(N399), .B(N393), .Z(N400) );
  GTECH_AND2 C720 ( .A(d1stg_opdec[2]), .B(d1stg_denorm_dbl_in1), .Z(N399) );
  GTECH_AND2 C724 ( .A(N407), .B(N398), .Z(div_norm_frac_in1_sng_norm) );
  GTECH_AND2 C725 ( .A(N404), .B(N406), .Z(N407) );
  GTECH_AND2 C726 ( .A(N402), .B(N403), .Z(N404) );
  GTECH_AND2 C727 ( .A(d1stg_opdec[2]), .B(d1stg_norm_sng_in1), .Z(N402) );
  GTECH_NOT I_91 ( .A(d1stg_snan_sng_in2), .Z(N403) );
  GTECH_OR2 C729 ( .A(N405), .B(d1stg_snan_sng_in1), .Z(N406) );
  GTECH_NOT I_92 ( .A(d1stg_qnan_sng_in2), .Z(N405) );
  GTECH_AND2 C732 ( .A(N410), .B(N398), .Z(div_norm_frac_in1_sng_dnrm) );
  GTECH_AND2 C733 ( .A(N409), .B(N405), .Z(N410) );
  GTECH_AND2 C734 ( .A(N408), .B(N403), .Z(N409) );
  GTECH_AND2 C735 ( .A(d1stg_opdec[2]), .B(d1stg_denorm_sng_in1), .Z(N408) );
  GTECH_OR2 C739 ( .A(N417), .B(N420), .Z(div_norm_frac_in2_dbl_norm) );
  GTECH_OR2 C740 ( .A(N415), .B(N416), .Z(N417) );
  GTECH_AND2 C741 ( .A(N413), .B(N414), .Z(N415) );
  GTECH_AND2 C742 ( .A(N411), .B(N412), .Z(N413) );
  GTECH_AND2 C743 ( .A(d2stg_opdec[2]), .B(d2stg_norm_dbl_in2), .Z(N411) );
  GTECH_NOT I_93 ( .A(d2stg_infnan_in), .Z(N412) );
  GTECH_NOT I_94 ( .A(d2stg_zero_in), .Z(N414) );
  GTECH_AND2 C746 ( .A(d1stg_opdec[2]), .B(d1stg_snan_dbl_in2), .Z(N416) );
  GTECH_AND2 C747 ( .A(N418), .B(N419), .Z(N420) );
  GTECH_AND2 C748 ( .A(d1stg_opdec[2]), .B(d1stg_qnan_dbl_in2), .Z(N418) );
  GTECH_NOT I_95 ( .A(d1stg_snan_dbl_in1), .Z(N419) );
  GTECH_AND2 C750 ( .A(N422), .B(N414), .Z(div_norm_frac_in2_dbl_dnrm) );
  GTECH_AND2 C751 ( .A(N421), .B(N412), .Z(N422) );
  GTECH_AND2 C752 ( .A(d2stg_opdec[2]), .B(d2stg_denorm_dbl_in2), .Z(N421) );
  GTECH_OR2 C755 ( .A(N427), .B(N430), .Z(div_norm_frac_in2_sng_norm) );
  GTECH_OR2 C756 ( .A(N425), .B(N426), .Z(N427) );
  GTECH_AND2 C757 ( .A(N424), .B(N414), .Z(N425) );
  GTECH_AND2 C758 ( .A(N423), .B(N412), .Z(N424) );
  GTECH_AND2 C759 ( .A(d2stg_opdec[2]), .B(d2stg_norm_sng_in2), .Z(N423) );
  GTECH_AND2 C762 ( .A(d1stg_opdec[2]), .B(d1stg_snan_sng_in2), .Z(N426) );
  GTECH_AND2 C763 ( .A(N428), .B(N429), .Z(N430) );
  GTECH_AND2 C764 ( .A(d1stg_opdec[2]), .B(d1stg_qnan_sng_in2), .Z(N428) );
  GTECH_NOT I_96 ( .A(d1stg_snan_sng_in1), .Z(N429) );
  GTECH_AND2 C766 ( .A(N432), .B(N414), .Z(div_norm_frac_in2_sng_dnrm) );
  GTECH_AND2 C767 ( .A(N431), .B(N412), .Z(N432) );
  GTECH_AND2 C768 ( .A(d2stg_opdec[2]), .B(d2stg_denorm_sng_in2), .Z(N431) );
  GTECH_OR2 C771 ( .A(N434), .B(N442), .Z(div_norm_inf) );
  GTECH_AND2 C772 ( .A(d2stg_opdec[2]), .B(N433), .Z(N434) );
  GTECH_OR2 C773 ( .A(d2stg_infnan_in), .B(d2stg_zero_in), .Z(N433) );
  GTECH_AND2 C774 ( .A(d1stg_opdec[2]), .B(N441), .Z(N442) );
  GTECH_OR2 C775 ( .A(N436), .B(N440), .Z(N441) );
  GTECH_AND2 C776 ( .A(d1stg_inf_in1), .B(N435), .Z(N436) );
  GTECH_NOT I_97 ( .A(d1stg_infnan_in2), .Z(N435) );
  GTECH_AND2 C778 ( .A(N438), .B(N439), .Z(N440) );
  GTECH_AND2 C779 ( .A(d1stg_zero_in2), .B(N437), .Z(N438) );
  GTECH_NOT I_98 ( .A(d1stg_infnan_in1), .Z(N437) );
  GTECH_NOT I_99 ( .A(d1stg_zero_in1), .Z(N439) );
  GTECH_AND2 C782 ( .A(d1stg_opdec[2]), .B(N443), .Z(div_norm_qnan) );
  GTECH_OR2 C783 ( .A(d1stg_2inf_in), .B(d1stg_2zero_in), .Z(N443) );
  GTECH_AND2 C784 ( .A(d1stg_opdec[2]), .B(N450), .Z(div_norm_zero) );
  GTECH_OR2 C785 ( .A(N445), .B(N449), .Z(N450) );
  GTECH_AND2 C786 ( .A(d1stg_inf_in2), .B(N444), .Z(N445) );
  GTECH_NOT I_100 ( .A(d1stg_infnan_in1), .Z(N444) );
  GTECH_AND2 C788 ( .A(N447), .B(N448), .Z(N449) );
  GTECH_AND2 C789 ( .A(d1stg_zero_in1), .B(N446), .Z(N447) );
  GTECH_NOT I_101 ( .A(d1stg_infnan_in2), .Z(N446) );
  GTECH_NOT I_102 ( .A(d1stg_zero_in2), .Z(N448) );
  GTECH_OR2 C792 ( .A(d4stg_fdiv), .B(d6stg_fdiv), .Z(div_frac_add_in2_load)
         );
  GTECH_AND2 C793 ( .A(N452), .B(N97), .Z(d6stg_frac_out_shl1) );
  GTECH_AND2 C794 ( .A(N451), .B(N6), .Z(N452) );
  GTECH_NOT I_103 ( .A(div_frac_out_54), .Z(N451) );
  GTECH_NOT I_104 ( .A(d6stg_frac_out_shl1), .Z(d6stg_frac_out_nosh) );
  GTECH_AND2 C798 ( .A(N454), .B(d8stg_step), .Z(div_frac_add_in1_add) );
  GTECH_AND2 C799 ( .A(d5stg_opdec[2]), .B(N453), .Z(N454) );
  GTECH_NOT I_105 ( .A(div_exp1[12]), .Z(N453) );
  GTECH_OR2 C801 ( .A(N457), .B(d6stg_fdiv), .Z(div_frac_add_in1_load) );
  GTECH_OR2 C802 ( .A(d4stg_fdiv), .B(N456), .Z(N457) );
  GTECH_AND2 C803 ( .A(N455), .B(d8stg_step), .Z(N456) );
  GTECH_AND2 C804 ( .A(d5stg_opdec[2]), .B(N453), .Z(N455) );
  GTECH_OR2 C806 ( .A(N458), .B(N460), .Z(d7stg_lsb_in) );
  GTECH_AND2 C807 ( .A(d6stg_fdivd), .B(d6stg_frac_2), .Z(N458) );
  GTECH_AND2 C808 ( .A(N459), .B(d6stg_frac_31), .Z(N460) );
  GTECH_NOT I_106 ( .A(d6stg_fdivd), .Z(N459) );
  GTECH_OR2 C810 ( .A(N461), .B(N463), .Z(d7stg_grd_in) );
  GTECH_AND2 C811 ( .A(d6stg_fdivd), .B(d6stg_frac_1), .Z(N461) );
  GTECH_AND2 C812 ( .A(N462), .B(d6stg_frac_30), .Z(N463) );
  GTECH_NOT I_107 ( .A(d6stg_fdivd), .Z(N462) );
  GTECH_OR2 C814 ( .A(N467), .B(div_frac_add_in1_neq_0), .Z(d7stg_stk_in) );
  GTECH_OR2 C815 ( .A(N464), .B(N466), .Z(N467) );
  GTECH_AND2 C816 ( .A(d6stg_fdivd), .B(d6stg_frac_0), .Z(N464) );
  GTECH_AND2 C817 ( .A(N465), .B(d6stg_frac_29), .Z(N466) );
  GTECH_NOT I_108 ( .A(d6stg_fdivd), .Z(N465) );
  GTECH_OR2 C819 ( .A(d7stg_grd), .B(d7stg_stk), .Z(N7) );
  GTECH_OR2 C820 ( .A(N473), .B(N479), .Z(d7stg_rndup) );
  GTECH_OR2 C821 ( .A(N470), .B(N472), .Z(N473) );
  GTECH_AND2 C822 ( .A(N469), .B(N7), .Z(N470) );
  GTECH_AND2 C823 ( .A(N106), .B(N468), .Z(N469) );
  GTECH_NOT I_109 ( .A(div_sign_out), .Z(N468) );
  GTECH_AND2 C825 ( .A(N471), .B(N7), .Z(N472) );
  GTECH_AND2 C826 ( .A(N107), .B(div_sign_out), .Z(N471) );
  GTECH_AND2 C827 ( .A(N109), .B(N478), .Z(N479) );
  GTECH_OR2 C828 ( .A(N474), .B(N477), .Z(N478) );
  GTECH_AND2 C829 ( .A(d7stg_grd), .B(d7stg_stk), .Z(N474) );
  GTECH_AND2 C830 ( .A(N476), .B(d7stg_lsb), .Z(N477) );
  GTECH_AND2 C831 ( .A(d7stg_grd), .B(N475), .Z(N476) );
  GTECH_NOT I_110 ( .A(d7stg_stk), .Z(N475) );
  GTECH_NOT I_111 ( .A(d7stg_rndup), .Z(d7stg_rndup_inv) );
  GTECH_OR2 C834 ( .A(N481), .B(N482), .Z(d7stg_to_0) );
  GTECH_OR2 C835 ( .A(N100), .B(N480), .Z(N481) );
  GTECH_AND2 C836 ( .A(N103), .B(div_sign_out), .Z(N480) );
  GTECH_AND2 C837 ( .A(N104), .B(N468), .Z(N482) );
  GTECH_NOT I_112 ( .A(d7stg_to_0), .Z(d7stg_to_0_inv) );
  GTECH_AND2 C840 ( .A(N484), .B(N485), .Z(div_frac_out_add_in1) );
  GTECH_AND2 C841 ( .A(d7stg_fdiv), .B(N483), .Z(N484) );
  GTECH_NOT I_113 ( .A(d7stg_rndup), .Z(N483) );
  GTECH_NOT I_114 ( .A(d7stg_in_of), .Z(N485) );
  GTECH_AND2 C844 ( .A(N486), .B(N487), .Z(div_frac_out_add) );
  GTECH_AND2 C845 ( .A(d7stg_fdiv), .B(d7stg_rndup), .Z(N486) );
  GTECH_NOT I_115 ( .A(d7stg_in_of), .Z(N487) );
  GTECH_AND2 C847 ( .A(N488), .B(d8stg_step), .Z(div_frac_out_shl1_dbl) );
  GTECH_AND2 C848 ( .A(d5stg_fdivd), .B(N453), .Z(N488) );
  GTECH_AND2 C850 ( .A(N489), .B(d8stg_step), .Z(div_frac_out_shl1_sng) );
  GTECH_AND2 C851 ( .A(d5stg_fdivs), .B(N453), .Z(N489) );
  GTECH_AND2 C853 ( .A(d7stg_fdiv), .B(d7stg_in_of), .Z(div_frac_out_of) );
  GTECH_OR2 C854 ( .A(N491), .B(div_frac_out_shl1_sng), .Z(div_frac_out_load)
         );
  GTECH_OR2 C855 ( .A(N490), .B(div_frac_out_shl1_dbl), .Z(N491) );
  GTECH_OR2 C856 ( .A(d4stg_fdiv), .B(d7stg_fdiv), .Z(N490) );
  GTECH_AND2 C857 ( .A(N495), .B(N500), .Z(div_expadd1_in1_dbl_in) );
  GTECH_OR2 C858 ( .A(N492), .B(N494), .Z(N495) );
  GTECH_AND2 C859 ( .A(d1stg_stepa), .B(inq_op[1]), .Z(N492) );
  GTECH_AND2 C860 ( .A(N493), .B(d1stg_dblopa[4]), .Z(N494) );
  GTECH_NOT I_116 ( .A(d1stg_stepa), .Z(N493) );
  GTECH_NOT I_117 ( .A(N499), .Z(N500) );
  GTECH_AND2 C863 ( .A(N497), .B(N498), .Z(N499) );
  GTECH_OR2 C864 ( .A(N496), .B(d3stg_fdiv), .Z(N497) );
  GTECH_OR2 C865 ( .A(d1stg_opdec[2]), .B(d2stg_opdec[2]), .Z(N496) );
  GTECH_NOT I_118 ( .A(reset), .Z(N498) );
  GTECH_AND2 C867 ( .A(N504), .B(N509), .Z(div_expadd1_in1_sng_in) );
  GTECH_OR2 C868 ( .A(N501), .B(N503), .Z(N504) );
  GTECH_AND2 C869 ( .A(d1stg_stepa), .B(inq_op[0]), .Z(N501) );
  GTECH_AND2 C870 ( .A(N502), .B(d1stg_sngopa[4]), .Z(N503) );
  GTECH_NOT I_119 ( .A(d1stg_stepa), .Z(N502) );
  GTECH_NOT I_120 ( .A(N508), .Z(N509) );
  GTECH_AND2 C873 ( .A(N506), .B(N507), .Z(N508) );
  GTECH_OR2 C874 ( .A(N505), .B(d3stg_fdiv), .Z(N506) );
  GTECH_OR2 C875 ( .A(d1stg_opdec[2]), .B(d2stg_opdec[2]), .Z(N505) );
  GTECH_NOT I_121 ( .A(reset), .Z(N507) );
  GTECH_OR2 C877 ( .A(N513), .B(d4stg_fdiv), .Z(div_exp1_expadd1) );
  GTECH_OR2 C878 ( .A(N512), .B(d3stg_fdiv), .Z(N513) );
  GTECH_OR2 C879 ( .A(d1stg_opdec[2]), .B(N511), .Z(N512) );
  GTECH_AND2 C880 ( .A(N510), .B(N414), .Z(N511) );
  GTECH_AND2 C881 ( .A(d2stg_opdec[2]), .B(N412), .Z(N510) );
  GTECH_AND2 C884 ( .A(div_expadd1_in2_exp_in2_dbl), .B(d2stg_max_exp), .Z(
        div_exp1_0835) );
  GTECH_AND2 C885 ( .A(div_expadd1_in2_exp_in2_sng), .B(d2stg_max_exp), .Z(
        div_exp1_0118) );
  GTECH_AND2 C886 ( .A(d2stg_opdec[2]), .B(d2stg_zero_exp), .Z(div_exp1_zero)
         );
  GTECH_OR2 C887 ( .A(N514), .B(d2stg_zero_in2), .Z(d2stg_max_exp) );
  GTECH_OR2 C888 ( .A(d2stg_nan_in), .B(d2stg_inf_in1), .Z(N514) );
  GTECH_OR2 C889 ( .A(N516), .B(N520), .Z(d2stg_zero_exp) );
  GTECH_AND2 C890 ( .A(d2stg_inf_in2), .B(N515), .Z(N516) );
  GTECH_NOT I_122 ( .A(d2stg_infnan_in1), .Z(N515) );
  GTECH_AND2 C892 ( .A(N518), .B(N519), .Z(N520) );
  GTECH_AND2 C893 ( .A(d2stg_zero_in1), .B(N517), .Z(N518) );
  GTECH_NOT I_123 ( .A(d2stg_infnan_in2), .Z(N517) );
  GTECH_NOT I_124 ( .A(d2stg_zero_in2), .Z(N519) );
  GTECH_OR2 C896 ( .A(N522), .B(d4stg_fdiv), .Z(div_exp1_load) );
  GTECH_OR2 C897 ( .A(N521), .B(d3stg_fdiv), .Z(N522) );
  GTECH_OR2 C898 ( .A(d1stg_opdec[2]), .B(d2stg_opdec[2]), .Z(N521) );
  GTECH_OR2 C899 ( .A(d6stg_opdec_in[2]), .B(d6stg_fdiv), .Z(
        div_expadd2_in1_exp_out_in) );
  GTECH_NOT I_125 ( .A(d5stg_fdivs), .Z(N8) );
  GTECH_OR2 C901 ( .A(N8), .B(d5stg_fdivs), .Z(N9) );
  GTECH_NOT I_126 ( .A(N524), .Z(div_expadd2_no_decr_inv_in) );
  GTECH_OR2 C906 ( .A(N523), .B(div_expadd2_12), .Z(N524) );
  GTECH_OR2 C907 ( .A(div_frac_out_53), .B(N10), .Z(N523) );
  GTECH_AND2 C908 ( .A(d5stg_opdec[2]), .B(d8stg_step), .Z(
        div_expadd2_no_decr_load) );
  GTECH_OR2 C909 ( .A(d5stg_opdec[2]), .B(d7stg_fdiv), .Z(div_expadd2_cin) );
  GTECH_AND2 C910 ( .A(d7stg_fdiv), .B(div_exp_out[12]), .Z(div_exp_out_zero)
         );
  GTECH_NOT I_127 ( .A(N527), .Z(div_exp_out_expadd22_inv) );
  GTECH_OR2 C912 ( .A(d6stg_fdiv), .B(N526), .Z(N527) );
  GTECH_AND2 C913 ( .A(N525), .B(d8stg_step), .Z(N526) );
  GTECH_AND2 C914 ( .A(d5stg_opdec[2]), .B(N63), .Z(N525) );
  GTECH_AND2 C915 ( .A(N534), .B(N535), .Z(div_exp_out_expadd2) );
  GTECH_OR2 C916 ( .A(N533), .B(d6stg_fdiv), .Z(N534) );
  GTECH_OR2 C917 ( .A(N530), .B(N532), .Z(N533) );
  GTECH_AND2 C918 ( .A(N528), .B(N529), .Z(N530) );
  GTECH_AND2 C919 ( .A(d7stg_fdiv), .B(d7stg_rndup), .Z(N528) );
  GTECH_NOT I_128 ( .A(d7stg_in_of), .Z(N529) );
  GTECH_AND2 C921 ( .A(N531), .B(d8stg_step), .Z(N532) );
  GTECH_AND2 C922 ( .A(d5stg_opdec[2]), .B(N69), .Z(N531) );
  GTECH_NOT I_129 ( .A(div_exp_out_zero), .Z(N535) );
  GTECH_AND2 C924 ( .A(d7stg_fdiv), .B(d7stg_in_of), .Z(div_exp_out_of) );
  GTECH_AND2 C925 ( .A(N537), .B(N535), .Z(div_exp_out_exp_out) );
  GTECH_AND2 C926 ( .A(d7stg_fdiv), .B(N536), .Z(N537) );
  GTECH_NOT I_130 ( .A(d7stg_in_of), .Z(N536) );
  GTECH_OR2 C929 ( .A(N540), .B(d7stg_fdiv), .Z(div_exp_out_load) );
  GTECH_OR2 C930 ( .A(N539), .B(d6stg_fdiv), .Z(N540) );
  GTECH_AND2 C931 ( .A(N538), .B(d8stg_step), .Z(N539) );
  GTECH_AND2 C932 ( .A(d5stg_opdec[2]), .B(N75), .Z(N538) );
endmodule


module fpu_div_exp_dp ( inq_in1, inq_in2, d1stg_step, d234stg_fdiv, 
        div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl, 
        div_expadd1_in2_exp_in2_sng, d3stg_fdiv, d4stg_fdiv, div_shl_cnt, 
        div_exp1_expadd1, div_exp1_0835, div_exp1_0118, div_exp1_zero, 
        div_exp1_load, div_expadd2_in1_exp_out, d5stg_fdiva, d5stg_fdivd, 
        d5stg_fdivs, d6stg_fdiv, d7stg_fdiv, div_expadd2_no_decr_inv, 
        div_expadd2_cin, div_exp_out_expadd2, div_exp_out_expadd22_inv, 
        div_exp_out_of, d7stg_to_0_inv, d7stg_fdivd, div_exp_out_exp_out, 
        d7stg_rndup_inv, div_frac_add_52_inv, div_exp_out_load, fdiv_clken_l, 
        rclk, div_exp1, div_expadd2_12, div_exp_out, div_exp_outa, se, si, so
 );
  input [62:52] inq_in1;
  input [62:52] inq_in2;
  input [5:0] div_shl_cnt;
  output [12:0] div_exp1;
  output [12:0] div_exp_out;
  output [10:0] div_exp_outa;
  input d1stg_step, d234stg_fdiv, div_expadd1_in1_dbl, div_expadd1_in1_sng,
         div_expadd1_in2_exp_in2_dbl, div_expadd1_in2_exp_in2_sng, d3stg_fdiv,
         d4stg_fdiv, div_exp1_expadd1, div_exp1_0835, div_exp1_0118,
         div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out, d5stg_fdiva,
         d5stg_fdivd, d5stg_fdivs, d6stg_fdiv, d7stg_fdiv,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd2,
         div_exp_out_expadd22_inv, div_exp_out_of, d7stg_to_0_inv, d7stg_fdivd,
         div_exp_out_exp_out, d7stg_rndup_inv, div_frac_add_52_inv,
         div_exp_out_load, fdiv_clken_l, rclk, se, si;
  output div_expadd2_12, so;
  wire   se_l, clk, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13,
         N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, net12817, net12818,
         net12819, net12820, net12821, net12822, net12823, net12824, net12825,
         net12826, net12827, net12828, net12829, net12830, net12831, net12832,
         net12833, net12834, net12835, net12836, net12837, net12838, net12839,
         net12840, net12841, net12842, net12843, net12844, net12845, net12846,
         net12847, net12848, net12849, net12850, net12851, net12852, net12853,
         net12854, net12855, net12856, net12857, net12858, net12859, net12860,
         net12861, net12862, net12863, net12864, net12865;
  wire   [10:0] div_exp_in1;
  wire   [10:0] div_exp_in2;
  wire   [12:0] div_expadd1_in1;
  wire   [12:0] div_expadd1_in2;
  wire   [12:0] div_expadd1;
  wire   [12:0] div_exp1_in;
  wire   [12:0] div_expadd2_in1;
  wire   [12:0] div_expadd2_in2;
  wire   [11:0] div_expadd2;
  wire   [12:0] div_exp_out_in;
  assign div_exp_outa[10] = div_exp_out[10];
  assign div_exp_outa[9] = div_exp_out[9];
  assign div_exp_outa[8] = div_exp_out[8];
  assign div_exp_outa[7] = div_exp_out[7];
  assign div_exp_outa[6] = div_exp_out[6];
  assign div_exp_outa[5] = div_exp_out[5];
  assign div_exp_outa[4] = div_exp_out[4];
  assign div_exp_outa[3] = div_exp_out[3];
  assign div_exp_outa[2] = div_exp_out[2];
  assign div_exp_outa[1] = div_exp_out[1];
  assign div_exp_outa[0] = div_exp_out[0];

  clken_buf ckbuf_div_exp_dp ( .clk(clk), .rclk(rclk), .enb_l(fdiv_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE11 i_div_exp_in1 ( .din(inq_in1), .en(d1stg_step), .clk(clk), .q(
        div_exp_in1), .se(se), .si({net12855, net12856, net12857, net12858, 
        net12859, net12860, net12861, net12862, net12863, net12864, net12865})
         );
  dffe_SIZE11 i_div_exp_in2 ( .din(inq_in2), .en(d1stg_step), .clk(clk), .q(
        div_exp_in2), .se(se), .si({net12844, net12845, net12846, net12847, 
        net12848, net12849, net12850, net12851, net12852, net12853, net12854})
         );
  dffe_SIZE13 i_div_exp1 ( .din(div_exp1_in), .en(div_exp1_load), .clk(clk), 
        .q(div_exp1), .se(se), .si({net12831, net12832, net12833, net12834, 
        net12835, net12836, net12837, net12838, net12839, net12840, net12841, 
        net12842, net12843}) );
  dffe_SIZE13 i_div_exp_out ( .din(div_exp_out_in), .en(div_exp_out_load), 
        .clk(clk), .q(div_exp_out), .se(se), .si({net12818, net12819, net12820, 
        net12821, net12822, net12823, net12824, net12825, net12826, net12827, 
        net12828, net12829, net12830}) );
  ADD_UNS_OP add_205 ( .A(div_expadd1_in1), .B(div_expadd1_in2), .Z(
        div_expadd1) );
  ADD_UNS_OP add_249 ( .A(div_expadd2_in1), .B(div_expadd2_in2), .Z({N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  ADD_UNS_OP add_249_2 ( .A({N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, 
        N0}), .B(div_expadd2_cin), .Z({div_expadd2_12, div_expadd2}) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_AND2 C86 ( .A(d234stg_fdiv), .B(div_exp1[12]), .Z(div_expadd1_in1[12])
         );
  GTECH_AND2 C87 ( .A(d234stg_fdiv), .B(div_exp1[11]), .Z(div_expadd1_in1[11])
         );
  GTECH_OR2 C88 ( .A(N13), .B(N14), .Z(div_expadd1_in1[10]) );
  GTECH_AND2 C89 ( .A(d234stg_fdiv), .B(div_exp1[10]), .Z(N13) );
  GTECH_AND2 C90 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[10]), .Z(N14) );
  GTECH_OR2 C91 ( .A(N15), .B(N16), .Z(div_expadd1_in1[9]) );
  GTECH_AND2 C92 ( .A(d234stg_fdiv), .B(div_exp1[9]), .Z(N15) );
  GTECH_AND2 C93 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[9]), .Z(N16) );
  GTECH_OR2 C94 ( .A(N17), .B(N18), .Z(div_expadd1_in1[8]) );
  GTECH_AND2 C95 ( .A(d234stg_fdiv), .B(div_exp1[8]), .Z(N17) );
  GTECH_AND2 C96 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[8]), .Z(N18) );
  GTECH_OR2 C97 ( .A(N21), .B(N22), .Z(div_expadd1_in1[7]) );
  GTECH_OR2 C98 ( .A(N19), .B(N20), .Z(N21) );
  GTECH_AND2 C99 ( .A(d234stg_fdiv), .B(div_exp1[7]), .Z(N19) );
  GTECH_AND2 C100 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[7]), .Z(N20) );
  GTECH_AND2 C101 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[10]), .Z(N22) );
  GTECH_OR2 C102 ( .A(N25), .B(N26), .Z(div_expadd1_in1[6]) );
  GTECH_OR2 C103 ( .A(N23), .B(N24), .Z(N25) );
  GTECH_AND2 C104 ( .A(d234stg_fdiv), .B(div_exp1[6]), .Z(N23) );
  GTECH_AND2 C105 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[6]), .Z(N24) );
  GTECH_AND2 C106 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[9]), .Z(N26) );
  GTECH_OR2 C107 ( .A(N29), .B(N30), .Z(div_expadd1_in1[5]) );
  GTECH_OR2 C108 ( .A(N27), .B(N28), .Z(N29) );
  GTECH_AND2 C109 ( .A(d234stg_fdiv), .B(div_exp1[5]), .Z(N27) );
  GTECH_AND2 C110 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[5]), .Z(N28) );
  GTECH_AND2 C111 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[8]), .Z(N30) );
  GTECH_OR2 C112 ( .A(N33), .B(N34), .Z(div_expadd1_in1[4]) );
  GTECH_OR2 C113 ( .A(N31), .B(N32), .Z(N33) );
  GTECH_AND2 C114 ( .A(d234stg_fdiv), .B(div_exp1[4]), .Z(N31) );
  GTECH_AND2 C115 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[4]), .Z(N32) );
  GTECH_AND2 C116 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[7]), .Z(N34) );
  GTECH_OR2 C117 ( .A(N37), .B(N38), .Z(div_expadd1_in1[3]) );
  GTECH_OR2 C118 ( .A(N35), .B(N36), .Z(N37) );
  GTECH_AND2 C119 ( .A(d234stg_fdiv), .B(div_exp1[3]), .Z(N35) );
  GTECH_AND2 C120 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[3]), .Z(N36) );
  GTECH_AND2 C121 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[6]), .Z(N38) );
  GTECH_OR2 C122 ( .A(N41), .B(N42), .Z(div_expadd1_in1[2]) );
  GTECH_OR2 C123 ( .A(N39), .B(N40), .Z(N41) );
  GTECH_AND2 C124 ( .A(d234stg_fdiv), .B(div_exp1[2]), .Z(N39) );
  GTECH_AND2 C125 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[2]), .Z(N40) );
  GTECH_AND2 C126 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[5]), .Z(N42) );
  GTECH_OR2 C127 ( .A(N45), .B(N46), .Z(div_expadd1_in1[1]) );
  GTECH_OR2 C128 ( .A(N43), .B(N44), .Z(N45) );
  GTECH_AND2 C129 ( .A(d234stg_fdiv), .B(div_exp1[1]), .Z(N43) );
  GTECH_AND2 C130 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[1]), .Z(N44) );
  GTECH_AND2 C131 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[4]), .Z(N46) );
  GTECH_OR2 C132 ( .A(N49), .B(N50), .Z(div_expadd1_in1[0]) );
  GTECH_OR2 C133 ( .A(N47), .B(N48), .Z(N49) );
  GTECH_AND2 C134 ( .A(d234stg_fdiv), .B(div_exp1[0]), .Z(N47) );
  GTECH_AND2 C135 ( .A(div_expadd1_in1_dbl), .B(div_exp_in1[0]), .Z(N48) );
  GTECH_AND2 C136 ( .A(div_expadd1_in1_sng), .B(div_exp_in1[3]), .Z(N50) );
  GTECH_OR2 C137 ( .A(N51), .B(d3stg_fdiv), .Z(div_expadd1_in2[12]) );
  GTECH_OR2 C138 ( .A(div_expadd1_in2_exp_in2_dbl), .B(
        div_expadd1_in2_exp_in2_sng), .Z(N51) );
  GTECH_OR2 C139 ( .A(N52), .B(d3stg_fdiv), .Z(div_expadd1_in2[11]) );
  GTECH_OR2 C140 ( .A(div_expadd1_in2_exp_in2_dbl), .B(
        div_expadd1_in2_exp_in2_sng), .Z(N52) );
  GTECH_OR2 C141 ( .A(N56), .B(d3stg_fdiv), .Z(div_expadd1_in2[10]) );
  GTECH_OR2 C142 ( .A(N55), .B(div_expadd1_in2_exp_in2_sng), .Z(N56) );
  GTECH_OR2 C143 ( .A(div_expadd1_in1_dbl), .B(N54), .Z(N55) );
  GTECH_AND2 C144 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N53), .Z(N54) );
  GTECH_NOT I_1 ( .A(div_exp_in2[10]), .Z(N53) );
  GTECH_OR2 C146 ( .A(N59), .B(d3stg_fdiv), .Z(div_expadd1_in2[9]) );
  GTECH_OR2 C147 ( .A(N58), .B(div_expadd1_in2_exp_in2_sng), .Z(N59) );
  GTECH_AND2 C148 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N57), .Z(N58) );
  GTECH_NOT I_2 ( .A(div_exp_in2[9]), .Z(N57) );
  GTECH_OR2 C150 ( .A(N62), .B(d3stg_fdiv), .Z(div_expadd1_in2[8]) );
  GTECH_OR2 C151 ( .A(N61), .B(div_expadd1_in2_exp_in2_sng), .Z(N62) );
  GTECH_AND2 C152 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N60), .Z(N61) );
  GTECH_NOT I_3 ( .A(div_exp_in2[8]), .Z(N60) );
  GTECH_OR2 C154 ( .A(N67), .B(d3stg_fdiv), .Z(div_expadd1_in2[7]) );
  GTECH_OR2 C155 ( .A(N65), .B(N66), .Z(N67) );
  GTECH_OR2 C156 ( .A(div_expadd1_in1_sng), .B(N64), .Z(N65) );
  GTECH_AND2 C157 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N63), .Z(N64) );
  GTECH_NOT I_4 ( .A(div_exp_in2[7]), .Z(N63) );
  GTECH_AND2 C159 ( .A(div_expadd1_in2_exp_in2_sng), .B(N53), .Z(N66) );
  GTECH_OR2 C161 ( .A(N71), .B(d3stg_fdiv), .Z(div_expadd1_in2[6]) );
  GTECH_OR2 C162 ( .A(N69), .B(N70), .Z(N71) );
  GTECH_AND2 C163 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N68), .Z(N69) );
  GTECH_NOT I_5 ( .A(div_exp_in2[6]), .Z(N68) );
  GTECH_AND2 C165 ( .A(div_expadd1_in2_exp_in2_sng), .B(N57), .Z(N70) );
  GTECH_OR2 C167 ( .A(N79), .B(N80), .Z(div_expadd1_in2[5]) );
  GTECH_OR2 C168 ( .A(N76), .B(N78), .Z(N79) );
  GTECH_OR2 C169 ( .A(N74), .B(N75), .Z(N76) );
  GTECH_OR2 C170 ( .A(div_expadd1_in1_dbl), .B(N73), .Z(N74) );
  GTECH_AND2 C171 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N72), .Z(N73) );
  GTECH_NOT I_6 ( .A(div_exp_in2[5]), .Z(N72) );
  GTECH_AND2 C173 ( .A(div_expadd1_in2_exp_in2_sng), .B(N60), .Z(N75) );
  GTECH_AND2 C175 ( .A(d3stg_fdiv), .B(N77), .Z(N78) );
  GTECH_NOT I_7 ( .A(div_shl_cnt[5]), .Z(N77) );
  GTECH_AND2 C177 ( .A(d4stg_fdiv), .B(div_shl_cnt[5]), .Z(N80) );
  GTECH_OR2 C178 ( .A(N89), .B(N90), .Z(div_expadd1_in2[4]) );
  GTECH_OR2 C179 ( .A(N86), .B(N88), .Z(N89) );
  GTECH_OR2 C180 ( .A(N84), .B(N85), .Z(N86) );
  GTECH_OR2 C181 ( .A(N81), .B(N83), .Z(N84) );
  GTECH_OR2 C182 ( .A(div_expadd1_in1_dbl), .B(div_expadd1_in1_sng), .Z(N81)
         );
  GTECH_AND2 C183 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N82), .Z(N83) );
  GTECH_NOT I_8 ( .A(div_exp_in2[4]), .Z(N82) );
  GTECH_AND2 C185 ( .A(div_expadd1_in2_exp_in2_sng), .B(N63), .Z(N85) );
  GTECH_AND2 C187 ( .A(d3stg_fdiv), .B(N87), .Z(N88) );
  GTECH_NOT I_9 ( .A(div_shl_cnt[4]), .Z(N87) );
  GTECH_AND2 C189 ( .A(d4stg_fdiv), .B(div_shl_cnt[4]), .Z(N90) );
  GTECH_OR2 C190 ( .A(N98), .B(N99), .Z(div_expadd1_in2[3]) );
  GTECH_OR2 C191 ( .A(N95), .B(N97), .Z(N98) );
  GTECH_OR2 C192 ( .A(N93), .B(N94), .Z(N95) );
  GTECH_OR2 C193 ( .A(div_expadd1_in1_sng), .B(N92), .Z(N93) );
  GTECH_AND2 C194 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N91), .Z(N92) );
  GTECH_NOT I_10 ( .A(div_exp_in2[3]), .Z(N91) );
  GTECH_AND2 C196 ( .A(div_expadd1_in2_exp_in2_sng), .B(N68), .Z(N94) );
  GTECH_AND2 C198 ( .A(d3stg_fdiv), .B(N96), .Z(N97) );
  GTECH_NOT I_11 ( .A(div_shl_cnt[3]), .Z(N96) );
  GTECH_AND2 C200 ( .A(d4stg_fdiv), .B(div_shl_cnt[3]), .Z(N99) );
  GTECH_OR2 C201 ( .A(N107), .B(N108), .Z(div_expadd1_in2[2]) );
  GTECH_OR2 C202 ( .A(N104), .B(N106), .Z(N107) );
  GTECH_OR2 C203 ( .A(N102), .B(N103), .Z(N104) );
  GTECH_OR2 C204 ( .A(div_expadd1_in1_dbl), .B(N101), .Z(N102) );
  GTECH_AND2 C205 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N100), .Z(N101) );
  GTECH_NOT I_12 ( .A(div_exp_in2[2]), .Z(N100) );
  GTECH_AND2 C207 ( .A(div_expadd1_in2_exp_in2_sng), .B(N72), .Z(N103) );
  GTECH_AND2 C209 ( .A(d3stg_fdiv), .B(N105), .Z(N106) );
  GTECH_NOT I_13 ( .A(div_shl_cnt[2]), .Z(N105) );
  GTECH_AND2 C211 ( .A(d4stg_fdiv), .B(div_shl_cnt[2]), .Z(N108) );
  GTECH_OR2 C212 ( .A(N116), .B(N117), .Z(div_expadd1_in2[1]) );
  GTECH_OR2 C213 ( .A(N113), .B(N115), .Z(N116) );
  GTECH_OR2 C214 ( .A(N111), .B(N112), .Z(N113) );
  GTECH_OR2 C215 ( .A(div_expadd1_in1_dbl), .B(N110), .Z(N111) );
  GTECH_AND2 C216 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N109), .Z(N110) );
  GTECH_NOT I_14 ( .A(div_exp_in2[1]), .Z(N109) );
  GTECH_AND2 C218 ( .A(div_expadd1_in2_exp_in2_sng), .B(N82), .Z(N112) );
  GTECH_AND2 C220 ( .A(d3stg_fdiv), .B(N114), .Z(N115) );
  GTECH_NOT I_15 ( .A(div_shl_cnt[1]), .Z(N114) );
  GTECH_AND2 C222 ( .A(d4stg_fdiv), .B(div_shl_cnt[1]), .Z(N117) );
  GTECH_OR2 C223 ( .A(N125), .B(N126), .Z(div_expadd1_in2[0]) );
  GTECH_OR2 C224 ( .A(N122), .B(N124), .Z(N125) );
  GTECH_OR2 C225 ( .A(N120), .B(N121), .Z(N122) );
  GTECH_OR2 C226 ( .A(div_expadd1_in1_sng), .B(N119), .Z(N120) );
  GTECH_AND2 C227 ( .A(div_expadd1_in2_exp_in2_dbl), .B(N118), .Z(N119) );
  GTECH_NOT I_16 ( .A(div_exp_in2[0]), .Z(N118) );
  GTECH_AND2 C229 ( .A(div_expadd1_in2_exp_in2_sng), .B(N91), .Z(N121) );
  GTECH_AND2 C231 ( .A(d3stg_fdiv), .B(N123), .Z(N124) );
  GTECH_NOT I_17 ( .A(div_shl_cnt[0]), .Z(N123) );
  GTECH_AND2 C233 ( .A(d4stg_fdiv), .B(div_shl_cnt[0]), .Z(N126) );
  GTECH_AND2 C234 ( .A(div_exp1_expadd1), .B(div_expadd1[12]), .Z(
        div_exp1_in[12]) );
  GTECH_OR2 C235 ( .A(N127), .B(div_exp1_0835), .Z(div_exp1_in[11]) );
  GTECH_AND2 C236 ( .A(div_exp1_expadd1), .B(div_expadd1[11]), .Z(N127) );
  GTECH_AND2 C237 ( .A(div_exp1_expadd1), .B(div_expadd1[10]), .Z(
        div_exp1_in[10]) );
  GTECH_AND2 C238 ( .A(div_exp1_expadd1), .B(div_expadd1[9]), .Z(
        div_exp1_in[9]) );
  GTECH_OR2 C239 ( .A(N128), .B(div_exp1_0118), .Z(div_exp1_in[8]) );
  GTECH_AND2 C240 ( .A(div_exp1_expadd1), .B(div_expadd1[8]), .Z(N128) );
  GTECH_AND2 C241 ( .A(div_exp1_expadd1), .B(div_expadd1[7]), .Z(
        div_exp1_in[7]) );
  GTECH_AND2 C242 ( .A(div_exp1_expadd1), .B(div_expadd1[6]), .Z(
        div_exp1_in[6]) );
  GTECH_OR2 C243 ( .A(N129), .B(div_exp1_0835), .Z(div_exp1_in[5]) );
  GTECH_AND2 C244 ( .A(div_exp1_expadd1), .B(div_expadd1[5]), .Z(N129) );
  GTECH_OR2 C245 ( .A(N131), .B(div_exp1_0118), .Z(div_exp1_in[4]) );
  GTECH_OR2 C246 ( .A(N130), .B(div_exp1_0835), .Z(N131) );
  GTECH_AND2 C247 ( .A(div_exp1_expadd1), .B(div_expadd1[4]), .Z(N130) );
  GTECH_OR2 C248 ( .A(N132), .B(div_exp1_0118), .Z(div_exp1_in[3]) );
  GTECH_AND2 C249 ( .A(div_exp1_expadd1), .B(div_expadd1[3]), .Z(N132) );
  GTECH_OR2 C250 ( .A(N133), .B(div_exp1_0835), .Z(div_exp1_in[2]) );
  GTECH_AND2 C251 ( .A(div_exp1_expadd1), .B(div_expadd1[2]), .Z(N133) );
  GTECH_AND2 C252 ( .A(div_exp1_expadd1), .B(div_expadd1[1]), .Z(
        div_exp1_in[1]) );
  GTECH_OR2 C253 ( .A(N134), .B(div_exp1_0835), .Z(div_exp1_in[0]) );
  GTECH_AND2 C254 ( .A(div_exp1_expadd1), .B(div_expadd1[0]), .Z(N134) );
  GTECH_OR2 C255 ( .A(N135), .B(N136), .Z(div_expadd2_in1[12]) );
  GTECH_AND2 C256 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[12]), .Z(N135)
         );
  GTECH_AND2 C257 ( .A(d5stg_fdiva), .B(div_exp1[12]), .Z(N136) );
  GTECH_OR2 C258 ( .A(N137), .B(N138), .Z(div_expadd2_in1[11]) );
  GTECH_AND2 C259 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[11]), .Z(N137)
         );
  GTECH_AND2 C260 ( .A(d5stg_fdiva), .B(div_exp1[11]), .Z(N138) );
  GTECH_OR2 C261 ( .A(N139), .B(N140), .Z(div_expadd2_in1[10]) );
  GTECH_AND2 C262 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[10]), .Z(N139)
         );
  GTECH_AND2 C263 ( .A(d5stg_fdiva), .B(div_exp1[10]), .Z(N140) );
  GTECH_OR2 C264 ( .A(N141), .B(N142), .Z(div_expadd2_in1[9]) );
  GTECH_AND2 C265 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[9]), .Z(N141)
         );
  GTECH_AND2 C266 ( .A(d5stg_fdiva), .B(div_exp1[9]), .Z(N142) );
  GTECH_OR2 C267 ( .A(N143), .B(N144), .Z(div_expadd2_in1[8]) );
  GTECH_AND2 C268 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[8]), .Z(N143)
         );
  GTECH_AND2 C269 ( .A(d5stg_fdiva), .B(div_exp1[8]), .Z(N144) );
  GTECH_OR2 C270 ( .A(N145), .B(N146), .Z(div_expadd2_in1[7]) );
  GTECH_AND2 C271 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[7]), .Z(N145)
         );
  GTECH_AND2 C272 ( .A(d5stg_fdiva), .B(div_exp1[7]), .Z(N146) );
  GTECH_OR2 C273 ( .A(N147), .B(N148), .Z(div_expadd2_in1[6]) );
  GTECH_AND2 C274 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[6]), .Z(N147)
         );
  GTECH_AND2 C275 ( .A(d5stg_fdiva), .B(div_exp1[6]), .Z(N148) );
  GTECH_OR2 C276 ( .A(N149), .B(N150), .Z(div_expadd2_in1[5]) );
  GTECH_AND2 C277 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[5]), .Z(N149)
         );
  GTECH_AND2 C278 ( .A(d5stg_fdiva), .B(div_exp1[5]), .Z(N150) );
  GTECH_OR2 C279 ( .A(N151), .B(N152), .Z(div_expadd2_in1[4]) );
  GTECH_AND2 C280 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[4]), .Z(N151)
         );
  GTECH_AND2 C281 ( .A(d5stg_fdiva), .B(div_exp1[4]), .Z(N152) );
  GTECH_OR2 C282 ( .A(N153), .B(N154), .Z(div_expadd2_in1[3]) );
  GTECH_AND2 C283 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[3]), .Z(N153)
         );
  GTECH_AND2 C284 ( .A(d5stg_fdiva), .B(div_exp1[3]), .Z(N154) );
  GTECH_OR2 C285 ( .A(N155), .B(N156), .Z(div_expadd2_in1[2]) );
  GTECH_AND2 C286 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[2]), .Z(N155)
         );
  GTECH_AND2 C287 ( .A(d5stg_fdiva), .B(div_exp1[2]), .Z(N156) );
  GTECH_OR2 C288 ( .A(N157), .B(N158), .Z(div_expadd2_in1[1]) );
  GTECH_AND2 C289 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[1]), .Z(N157)
         );
  GTECH_AND2 C290 ( .A(d5stg_fdiva), .B(div_exp1[1]), .Z(N158) );
  GTECH_OR2 C291 ( .A(N159), .B(N160), .Z(div_expadd2_in1[0]) );
  GTECH_AND2 C292 ( .A(div_expadd2_in1_exp_out), .B(div_exp_out[0]), .Z(N159)
         );
  GTECH_AND2 C293 ( .A(d5stg_fdiva), .B(div_exp1[0]), .Z(N160) );
  GTECH_OR2 C294 ( .A(d5stg_fdiva), .B(N161), .Z(div_expadd2_in2[12]) );
  GTECH_AND2 C295 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N161) );
  GTECH_OR2 C296 ( .A(d5stg_fdiva), .B(N162), .Z(div_expadd2_in2[11]) );
  GTECH_AND2 C297 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N162) );
  GTECH_OR2 C298 ( .A(d5stg_fdiva), .B(N163), .Z(div_expadd2_in2[10]) );
  GTECH_AND2 C299 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N163) );
  GTECH_OR2 C300 ( .A(d5stg_fdiva), .B(N164), .Z(div_expadd2_in2[9]) );
  GTECH_AND2 C301 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N164) );
  GTECH_OR2 C302 ( .A(d5stg_fdiva), .B(N165), .Z(div_expadd2_in2[8]) );
  GTECH_AND2 C303 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N165) );
  GTECH_OR2 C304 ( .A(d5stg_fdiva), .B(N166), .Z(div_expadd2_in2[7]) );
  GTECH_AND2 C305 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N166) );
  GTECH_OR2 C306 ( .A(d5stg_fdiva), .B(N167), .Z(div_expadd2_in2[6]) );
  GTECH_AND2 C307 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N167) );
  GTECH_OR2 C308 ( .A(N168), .B(N169), .Z(div_expadd2_in2[5]) );
  GTECH_AND2 C309 ( .A(d5stg_fdiva), .B(d5stg_fdivs), .Z(N168) );
  GTECH_AND2 C310 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N169) );
  GTECH_AND2 C311 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(
        div_expadd2_in2[4]) );
  GTECH_OR2 C312 ( .A(N170), .B(N171), .Z(div_expadd2_in2[3]) );
  GTECH_AND2 C313 ( .A(d5stg_fdiva), .B(d5stg_fdivd), .Z(N170) );
  GTECH_AND2 C314 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N171) );
  GTECH_OR2 C315 ( .A(N172), .B(N173), .Z(div_expadd2_in2[2]) );
  GTECH_AND2 C316 ( .A(d5stg_fdiva), .B(d5stg_fdivs), .Z(N172) );
  GTECH_AND2 C317 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N173) );
  GTECH_OR2 C318 ( .A(d5stg_fdiva), .B(N174), .Z(div_expadd2_in2[1]) );
  GTECH_AND2 C319 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N174) );
  GTECH_OR2 C320 ( .A(N175), .B(N176), .Z(div_expadd2_in2[0]) );
  GTECH_AND2 C321 ( .A(d5stg_fdiva), .B(d5stg_fdivs), .Z(N175) );
  GTECH_AND2 C322 ( .A(d6stg_fdiv), .B(div_expadd2_no_decr_inv), .Z(N176) );
  GTECH_OR2 C323 ( .A(N180), .B(N183), .Z(div_exp_out_in[12]) );
  GTECH_AND2 C324 ( .A(N179), .B(div_expadd2_12), .Z(N180) );
  GTECH_AND2 C325 ( .A(div_exp_out_expadd2), .B(N178), .Z(N179) );
  GTECH_NOT I_18 ( .A(N177), .Z(N178) );
  GTECH_AND2 C327 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N177) );
  GTECH_AND2 C328 ( .A(N182), .B(div_exp_out[12]), .Z(N183) );
  GTECH_AND2 C329 ( .A(div_exp_out_exp_out), .B(N181), .Z(N182) );
  GTECH_OR2 C330 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N181) );
  GTECH_OR2 C331 ( .A(N187), .B(N190), .Z(div_exp_out_in[11]) );
  GTECH_AND2 C332 ( .A(N186), .B(div_expadd2[11]), .Z(N187) );
  GTECH_AND2 C333 ( .A(div_exp_out_expadd2), .B(N185), .Z(N186) );
  GTECH_NOT I_19 ( .A(N184), .Z(N185) );
  GTECH_AND2 C335 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N184) );
  GTECH_AND2 C336 ( .A(N189), .B(div_exp_out[11]), .Z(N190) );
  GTECH_AND2 C337 ( .A(div_exp_out_exp_out), .B(N188), .Z(N189) );
  GTECH_OR2 C338 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N188) );
  GTECH_OR2 C339 ( .A(N196), .B(N199), .Z(div_exp_out_in[10]) );
  GTECH_OR2 C340 ( .A(N194), .B(N195), .Z(N196) );
  GTECH_AND2 C341 ( .A(N193), .B(div_expadd2[10]), .Z(N194) );
  GTECH_AND2 C342 ( .A(div_exp_out_expadd2), .B(N192), .Z(N193) );
  GTECH_NOT I_20 ( .A(N191), .Z(N192) );
  GTECH_AND2 C344 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N191) );
  GTECH_AND2 C345 ( .A(div_exp_out_of), .B(d7stg_fdivd), .Z(N195) );
  GTECH_AND2 C346 ( .A(N198), .B(div_exp_out[10]), .Z(N199) );
  GTECH_AND2 C347 ( .A(div_exp_out_exp_out), .B(N197), .Z(N198) );
  GTECH_OR2 C348 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N197) );
  GTECH_OR2 C349 ( .A(N205), .B(N208), .Z(div_exp_out_in[9]) );
  GTECH_OR2 C350 ( .A(N203), .B(N204), .Z(N205) );
  GTECH_AND2 C351 ( .A(N202), .B(div_expadd2[9]), .Z(N203) );
  GTECH_AND2 C352 ( .A(div_exp_out_expadd2), .B(N201), .Z(N202) );
  GTECH_NOT I_21 ( .A(N200), .Z(N201) );
  GTECH_AND2 C354 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N200) );
  GTECH_AND2 C355 ( .A(div_exp_out_of), .B(d7stg_fdivd), .Z(N204) );
  GTECH_AND2 C356 ( .A(N207), .B(div_exp_out[9]), .Z(N208) );
  GTECH_AND2 C357 ( .A(div_exp_out_exp_out), .B(N206), .Z(N207) );
  GTECH_OR2 C358 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N206) );
  GTECH_OR2 C359 ( .A(N214), .B(N217), .Z(div_exp_out_in[8]) );
  GTECH_OR2 C360 ( .A(N212), .B(N213), .Z(N214) );
  GTECH_AND2 C361 ( .A(N211), .B(div_expadd2[8]), .Z(N212) );
  GTECH_AND2 C362 ( .A(div_exp_out_expadd2), .B(N210), .Z(N211) );
  GTECH_NOT I_22 ( .A(N209), .Z(N210) );
  GTECH_AND2 C364 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N209) );
  GTECH_AND2 C365 ( .A(div_exp_out_of), .B(d7stg_fdivd), .Z(N213) );
  GTECH_AND2 C366 ( .A(N216), .B(div_exp_out[8]), .Z(N217) );
  GTECH_AND2 C367 ( .A(div_exp_out_exp_out), .B(N215), .Z(N216) );
  GTECH_OR2 C368 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N215) );
  GTECH_OR2 C369 ( .A(N222), .B(N225), .Z(div_exp_out_in[7]) );
  GTECH_OR2 C370 ( .A(N221), .B(div_exp_out_of), .Z(N222) );
  GTECH_AND2 C371 ( .A(N220), .B(div_expadd2[7]), .Z(N221) );
  GTECH_AND2 C372 ( .A(div_exp_out_expadd2), .B(N219), .Z(N220) );
  GTECH_NOT I_23 ( .A(N218), .Z(N219) );
  GTECH_AND2 C374 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N218) );
  GTECH_AND2 C375 ( .A(N224), .B(div_exp_out[7]), .Z(N225) );
  GTECH_AND2 C376 ( .A(div_exp_out_exp_out), .B(N223), .Z(N224) );
  GTECH_OR2 C377 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N223) );
  GTECH_OR2 C378 ( .A(N230), .B(N233), .Z(div_exp_out_in[6]) );
  GTECH_OR2 C379 ( .A(N229), .B(div_exp_out_of), .Z(N230) );
  GTECH_AND2 C380 ( .A(N228), .B(div_expadd2[6]), .Z(N229) );
  GTECH_AND2 C381 ( .A(div_exp_out_expadd2), .B(N227), .Z(N228) );
  GTECH_NOT I_24 ( .A(N226), .Z(N227) );
  GTECH_AND2 C383 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N226) );
  GTECH_AND2 C384 ( .A(N232), .B(div_exp_out[6]), .Z(N233) );
  GTECH_AND2 C385 ( .A(div_exp_out_exp_out), .B(N231), .Z(N232) );
  GTECH_OR2 C386 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N231) );
  GTECH_OR2 C387 ( .A(N238), .B(N241), .Z(div_exp_out_in[5]) );
  GTECH_OR2 C388 ( .A(N237), .B(div_exp_out_of), .Z(N238) );
  GTECH_AND2 C389 ( .A(N236), .B(div_expadd2[5]), .Z(N237) );
  GTECH_AND2 C390 ( .A(div_exp_out_expadd2), .B(N235), .Z(N236) );
  GTECH_NOT I_25 ( .A(N234), .Z(N235) );
  GTECH_AND2 C392 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N234) );
  GTECH_AND2 C393 ( .A(N240), .B(div_exp_out[5]), .Z(N241) );
  GTECH_AND2 C394 ( .A(div_exp_out_exp_out), .B(N239), .Z(N240) );
  GTECH_OR2 C395 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N239) );
  GTECH_OR2 C396 ( .A(N246), .B(N249), .Z(div_exp_out_in[4]) );
  GTECH_OR2 C397 ( .A(N245), .B(div_exp_out_of), .Z(N246) );
  GTECH_AND2 C398 ( .A(N244), .B(div_expadd2[4]), .Z(N245) );
  GTECH_AND2 C399 ( .A(div_exp_out_expadd2), .B(N243), .Z(N244) );
  GTECH_NOT I_26 ( .A(N242), .Z(N243) );
  GTECH_AND2 C401 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N242) );
  GTECH_AND2 C402 ( .A(N248), .B(div_exp_out[4]), .Z(N249) );
  GTECH_AND2 C403 ( .A(div_exp_out_exp_out), .B(N247), .Z(N248) );
  GTECH_OR2 C404 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N247) );
  GTECH_OR2 C405 ( .A(N254), .B(N257), .Z(div_exp_out_in[3]) );
  GTECH_OR2 C406 ( .A(N253), .B(div_exp_out_of), .Z(N254) );
  GTECH_AND2 C407 ( .A(N252), .B(div_expadd2[3]), .Z(N253) );
  GTECH_AND2 C408 ( .A(div_exp_out_expadd2), .B(N251), .Z(N252) );
  GTECH_NOT I_27 ( .A(N250), .Z(N251) );
  GTECH_AND2 C410 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N250) );
  GTECH_AND2 C411 ( .A(N256), .B(div_exp_out[3]), .Z(N257) );
  GTECH_AND2 C412 ( .A(div_exp_out_exp_out), .B(N255), .Z(N256) );
  GTECH_OR2 C413 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N255) );
  GTECH_OR2 C414 ( .A(N262), .B(N265), .Z(div_exp_out_in[2]) );
  GTECH_OR2 C415 ( .A(N261), .B(div_exp_out_of), .Z(N262) );
  GTECH_AND2 C416 ( .A(N260), .B(div_expadd2[2]), .Z(N261) );
  GTECH_AND2 C417 ( .A(div_exp_out_expadd2), .B(N259), .Z(N260) );
  GTECH_NOT I_28 ( .A(N258), .Z(N259) );
  GTECH_AND2 C419 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N258) );
  GTECH_AND2 C420 ( .A(N264), .B(div_exp_out[2]), .Z(N265) );
  GTECH_AND2 C421 ( .A(div_exp_out_exp_out), .B(N263), .Z(N264) );
  GTECH_OR2 C422 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N263) );
  GTECH_OR2 C423 ( .A(N270), .B(N273), .Z(div_exp_out_in[1]) );
  GTECH_OR2 C424 ( .A(N269), .B(div_exp_out_of), .Z(N270) );
  GTECH_AND2 C425 ( .A(N268), .B(div_expadd2[1]), .Z(N269) );
  GTECH_AND2 C426 ( .A(div_exp_out_expadd2), .B(N267), .Z(N268) );
  GTECH_NOT I_29 ( .A(N266), .Z(N267) );
  GTECH_AND2 C428 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N266) );
  GTECH_AND2 C429 ( .A(N272), .B(div_exp_out[1]), .Z(N273) );
  GTECH_AND2 C430 ( .A(div_exp_out_exp_out), .B(N271), .Z(N272) );
  GTECH_OR2 C431 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N271) );
  GTECH_OR2 C432 ( .A(N279), .B(N282), .Z(div_exp_out_in[0]) );
  GTECH_OR2 C433 ( .A(N277), .B(N278), .Z(N279) );
  GTECH_AND2 C434 ( .A(N276), .B(div_expadd2[0]), .Z(N277) );
  GTECH_AND2 C435 ( .A(div_exp_out_expadd2), .B(N275), .Z(N276) );
  GTECH_NOT I_30 ( .A(N274), .Z(N275) );
  GTECH_AND2 C437 ( .A(div_frac_add_52_inv), .B(div_exp_out_expadd22_inv), .Z(
        N274) );
  GTECH_AND2 C438 ( .A(div_exp_out_of), .B(d7stg_to_0_inv), .Z(N278) );
  GTECH_AND2 C439 ( .A(N281), .B(div_exp_out[0]), .Z(N282) );
  GTECH_AND2 C440 ( .A(div_exp_out_exp_out), .B(N280), .Z(N281) );
  GTECH_OR2 C441 ( .A(div_frac_add_52_inv), .B(d7stg_rndup_inv), .Z(N280) );
endmodule


module dff_SIZE53 ( din, clk, q, se, si, so );
  input [52:0] din;
  output [52:0] q;
  input [52:0] si;
  output [52:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55;
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C63 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module dff_SIZE12 ( din, clk, q, se, si, so );
  input [11:0] din;
  output [11:0] q;
  input [11:0] si;
  output [11:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14;
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C22 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module fpu_div_frac_dp ( inq_in1, inq_in2, d1stg_step, 
        div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm, 
        div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm, 
        div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm, 
        div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf, 
        div_norm_qnan, d1stg_dblop, div_norm_zero, d1stg_snan_dbl_in1, 
        d1stg_snan_sng_in1, d1stg_snan_dbl_in2, d1stg_snan_sng_in2, d3stg_fdiv, 
        d6stg_fdiv, d6stg_fdivd, d6stg_fdivs, div_frac_add_in2_load, 
        d6stg_frac_out_shl1, d6stg_frac_out_nosh, d4stg_fdiv, 
        div_frac_add_in1_add, div_frac_add_in1_load, d5stg_fdivb, 
        div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl, 
        div_frac_out_shl1_sng, div_frac_out_of, d7stg_to_0, div_frac_out_load, 
        fdiv_clken_l, rclk, div_shl_cnt, d6stg_frac_0, d6stg_frac_1, 
        d6stg_frac_2, d6stg_frac_29, d6stg_frac_30, d6stg_frac_31, 
        div_frac_add_in1_neq_0, div_frac_add_52_inv, div_frac_add_52_inva, 
        div_frac_out_54_53, div_frac_outa, se, si, so );
  input [54:0] inq_in1;
  input [54:0] inq_in2;
  output [5:0] div_shl_cnt;
  output [1:0] div_frac_out_54_53;
  output [51:0] div_frac_outa;
  input d1stg_step, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm,
         div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm,
         div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm,
         div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf,
         div_norm_qnan, d1stg_dblop, div_norm_zero, d1stg_snan_dbl_in1,
         d1stg_snan_sng_in1, d1stg_snan_dbl_in2, d1stg_snan_sng_in2,
         d3stg_fdiv, d6stg_fdiv, d6stg_fdivd, d6stg_fdivs,
         div_frac_add_in2_load, d6stg_frac_out_shl1, d6stg_frac_out_nosh,
         d4stg_fdiv, div_frac_add_in1_add, div_frac_add_in1_load, d5stg_fdivb,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, d7stg_to_0, div_frac_out_load,
         fdiv_clken_l, rclk, se, si;
  output d6stg_frac_0, d6stg_frac_1, d6stg_frac_2, d6stg_frac_29,
         d6stg_frac_30, d6stg_frac_31, div_frac_add_in1_neq_0,
         div_frac_add_52_inv, div_frac_add_52_inva, so;
  wire   se_l, clk, d6stg_frac_53, d6stg_frac_52, d6stg_frac_51, d6stg_frac_50,
         d6stg_frac_49, d6stg_frac_48, d6stg_frac_47, d6stg_frac_46,
         d6stg_frac_45, d6stg_frac_44, d6stg_frac_43, d6stg_frac_42,
         d6stg_frac_41, d6stg_frac_40, d6stg_frac_39, d6stg_frac_38,
         d6stg_frac_37, d6stg_frac_36, d6stg_frac_35, d6stg_frac_34,
         d6stg_frac_33, d6stg_frac_32, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435,
         N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479,
         N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490,
         N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523,
         N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534,
         N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545,
         N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556,
         N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600,
         N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611,
         N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732,
         N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743,
         N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754,
         N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765,
         N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776,
         N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787,
         N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798,
         N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809,
         N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864,
         N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875,
         N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886,
         N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897,
         N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908,
         N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919,
         N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930,
         N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026,
         N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056,
         N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066,
         N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076,
         N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086,
         N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096,
         N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106,
         N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116,
         N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126,
         N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136,
         N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146,
         N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156,
         N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166,
         N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176,
         N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186,
         N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196,
         N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206,
         N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216,
         N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226,
         N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236,
         N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246,
         N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256,
         N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266,
         N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276,
         N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286,
         N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296,
         N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306,
         N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316,
         N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326,
         N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336,
         N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346,
         N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356,
         N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366,
         N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376,
         N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386,
         N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396,
         N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406,
         N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416,
         N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426,
         N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436,
         N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446,
         N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456,
         N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466,
         N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476,
         N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486,
         N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496,
         N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506,
         N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516,
         N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526,
         N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536,
         N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546,
         N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556,
         N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566,
         N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576,
         N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586,
         N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596,
         N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606,
         N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616,
         N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626,
         N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636,
         N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646,
         N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656,
         N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666,
         N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676,
         N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686,
         N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696,
         N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706,
         N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716,
         N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726,
         N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736,
         N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746,
         N1747, N1748, net12313, net12314, net12315, net12316, net12317,
         net12318, net12319, net12320, net12321, net12322, net12323, net12324,
         net12325, net12326, net12327, net12328, net12329, net12330, net12331,
         net12332, net12333, net12334, net12335, net12336, net12337, net12338,
         net12339, net12340, net12341, net12342, net12343, net12344, net12345,
         net12346, net12347, net12348, net12349, net12350, net12351, net12352,
         net12353, net12354, net12355, net12356, net12357, net12358, net12359,
         net12360, net12361, net12362, net12363, net12364, net12365, net12366,
         net12367, net12368, net12369, net12370, net12371, net12372, net12373,
         net12374, net12375, net12376, net12377, net12378, net12379, net12380,
         net12381, net12382, net12383, net12384, net12385, net12386, net12387,
         net12388, net12389, net12390, net12391, net12392, net12393, net12394,
         net12395, net12396, net12397, net12398, net12399, net12400, net12401,
         net12402, net12403, net12404, net12405, net12406, net12407, net12408,
         net12409, net12410, net12411, net12412, net12413, net12414, net12415,
         net12416, net12417, net12418, net12419, net12420, net12421, net12422,
         net12423, net12424, net12425, net12426, net12427, net12428, net12429,
         net12430, net12431, net12432, net12433, net12434, net12435, net12436,
         net12437, net12438, net12439, net12440, net12441, net12442, net12443,
         net12444, net12445, net12446, net12447, net12448, net12449, net12450,
         net12451, net12452, net12453, net12454, net12455, net12456, net12457,
         net12458, net12459, net12460, net12461, net12462, net12463, net12464,
         net12465, net12466, net12467, net12468, net12469, net12470, net12471,
         net12472, net12473, net12474, net12475, net12476, net12477, net12478,
         net12479, net12480, net12481, net12482, net12483, net12484, net12485,
         net12486, net12487, net12488, net12489, net12490, net12491, net12492,
         net12493, net12494, net12495, net12496, net12497, net12498, net12499,
         net12500, net12501, net12502, net12503, net12504, net12505, net12506,
         net12507, net12508, net12509, net12510, net12511, net12512, net12513,
         net12514, net12515, net12516, net12517, net12518, net12519, net12520,
         net12521, net12522, net12523, net12524, net12525, net12526, net12527,
         net12528, net12529, net12530, net12531, net12532, net12533, net12534,
         net12535, net12536, net12537, net12538, net12539, net12540, net12541,
         net12542, net12543, net12544, net12545, net12546, net12547, net12548,
         net12549, net12550, net12551, net12552, net12553, net12554, net12555,
         net12556, net12557, net12558, net12559, net12560, net12561, net12562,
         net12563, net12564, net12565, net12566, net12567, net12568, net12569,
         net12570, net12571, net12572, net12573, net12574, net12575, net12576,
         net12577, net12578, net12579, net12580, net12581, net12582, net12583,
         net12584, net12585, net12586, net12587, net12588, net12589, net12590,
         net12591, net12592, net12593, net12594, net12595, net12596, net12597,
         net12598, net12599, net12600, net12601, net12602, net12603, net12604,
         net12605, net12606, net12607, net12608, net12609, net12610, net12611,
         net12612, net12613, net12614, net12615, net12616, net12617, net12618,
         net12619, net12620, net12621, net12622, net12623, net12624, net12625,
         net12626, net12627, net12628, net12629, net12630, net12631, net12632,
         net12633, net12634, net12635, net12636, net12637, net12638, net12639,
         net12640, net12641, net12642, net12643, net12644, net12645, net12646,
         net12647, net12648, net12649, net12650, net12651, net12652, net12653,
         net12654, net12655, net12656, net12657, net12658, net12659, net12660,
         net12661, net12662, net12663, net12664, net12665, net12666, net12667,
         net12668, net12669, net12670, net12671, net12672, net12673, net12674,
         net12675, net12676, net12677, net12678, net12679, net12680, net12681,
         net12682, net12683, net12684, net12685, net12686, net12687, net12688,
         net12689, net12690, net12691, net12692, net12693, net12694, net12695,
         net12696, net12697, net12698, net12699, net12700, net12701, net12702,
         net12703, net12704, net12705, net12706, net12707, net12708, net12709,
         net12710, net12711, net12712, net12713, net12714, net12715, net12716,
         net12717, net12718, net12719, net12720, net12721, net12722, net12723,
         net12724, net12725, net12726, net12727, net12728, net12729, net12730,
         net12731, net12732, net12733, net12734, net12735, net12736, net12737,
         net12738, net12739, net12740, net12741, net12742, net12743, net12744,
         net12745, net12746, net12747, net12748, net12749, net12750, net12751,
         net12752, net12753, net12754, net12755, net12756, net12757, net12758,
         net12759, net12760, net12761, net12762, net12763, net12764, net12765,
         net12766, net12767, net12768, net12769, net12770, net12771, net12772,
         net12773, net12774, net12775, net12776, net12777, net12778, net12779,
         net12780, net12781, net12782, net12783, net12784, net12785, net12786,
         net12787, net12788, net12789, net12790, net12791, net12792, net12793,
         net12794, net12795, net12796, net12797, net12798, net12799, net12800,
         net12801, net12802, net12803, net12804, net12805, net12806, net12807,
         net12808, net12809, net12810, net12811, net12812, net12813, net12814,
         net12815, net12816;
  wire   [54:0] div_frac_in1;
  wire   [54:0] div_frac_in2;
  wire   [52:0] div_norm_inv_in;
  wire   [52:0] div_norm_inv;
  wire   [52:0] div_norm;
  wire   [5:0] div_lead0;
  wire   [5:0] div_shl_cnta;
  wire   [52:0] div_shl_data;
  wire   [105:53] div_shl_tmp;
  wire   [54:0] div_shl_save;
  wire   [52:0] div_frac_add_in2_in;
  wire   [54:0] div_frac_add_in2;
  wire   [52:52] div_frac_out;
  wire   [28:3] d6stg_frac;
  wire   [54:0] div_frac_add;
  wire   [54:0] div_frac_add_in1;
  wire   [54:0] div_frac_add_in1_in;
  wire   [54:0] div_frac_add_in1a;
  wire   [54:0] div_frac_out_in;

  clken_buf ckbuf_div_frac_dp ( .clk(clk), .rclk(rclk), .enb_l(fdiv_clken_l), 
        .tmb_l(se_l) );
  dffe_SIZE55 i_div_frac_in1 ( .din(inq_in1), .en(d1stg_step), .clk(clk), .q(
        div_frac_in1), .se(se), .si({net12762, net12763, net12764, net12765, 
        net12766, net12767, net12768, net12769, net12770, net12771, net12772, 
        net12773, net12774, net12775, net12776, net12777, net12778, net12779, 
        net12780, net12781, net12782, net12783, net12784, net12785, net12786, 
        net12787, net12788, net12789, net12790, net12791, net12792, net12793, 
        net12794, net12795, net12796, net12797, net12798, net12799, net12800, 
        net12801, net12802, net12803, net12804, net12805, net12806, net12807, 
        net12808, net12809, net12810, net12811, net12812, net12813, net12814, 
        net12815, net12816}) );
  dffe_SIZE55 i_div_frac_in2 ( .din(inq_in2), .en(d1stg_step), .clk(clk), .q(
        div_frac_in2), .se(se), .si({net12707, net12708, net12709, net12710, 
        net12711, net12712, net12713, net12714, net12715, net12716, net12717, 
        net12718, net12719, net12720, net12721, net12722, net12723, net12724, 
        net12725, net12726, net12727, net12728, net12729, net12730, net12731, 
        net12732, net12733, net12734, net12735, net12736, net12737, net12738, 
        net12739, net12740, net12741, net12742, net12743, net12744, net12745, 
        net12746, net12747, net12748, net12749, net12750, net12751, net12752, 
        net12753, net12754, net12755, net12756, net12757, net12758, net12759, 
        net12760, net12761}) );
  dff_SIZE53 i_div_norm_inv ( .din(div_norm_inv_in), .clk(clk), .q(
        div_norm_inv), .se(se), .si({net12654, net12655, net12656, net12657, 
        net12658, net12659, net12660, net12661, net12662, net12663, net12664, 
        net12665, net12666, net12667, net12668, net12669, net12670, net12671, 
        net12672, net12673, net12674, net12675, net12676, net12677, net12678, 
        net12679, net12680, net12681, net12682, net12683, net12684, net12685, 
        net12686, net12687, net12688, net12689, net12690, net12691, net12692, 
        net12693, net12694, net12695, net12696, net12697, net12698, net12699, 
        net12700, net12701, net12702, net12703, net12704, net12705, net12706})
         );
  fpu_cnt_lead0_53b i_div_lead0 ( .din(div_norm), .lead0(div_lead0) );
  dff_SIZE12 i_dstg_xtra_regs ( .din({div_lead0, div_lead0}), .clk(clk), .q({
        div_shl_cnta, div_shl_cnt}), .se(se), .si({net12642, net12643, 
        net12644, net12645, net12646, net12647, net12648, net12649, net12650, 
        net12651, net12652, net12653}) );
  dff_SIZE53 i_div_shl_data ( .din(div_norm), .clk(clk), .q(div_shl_data), 
        .se(se), .si({net12589, net12590, net12591, net12592, net12593, 
        net12594, net12595, net12596, net12597, net12598, net12599, net12600, 
        net12601, net12602, net12603, net12604, net12605, net12606, net12607, 
        net12608, net12609, net12610, net12611, net12612, net12613, net12614, 
        net12615, net12616, net12617, net12618, net12619, net12620, net12621, 
        net12622, net12623, net12624, net12625, net12626, net12627, net12628, 
        net12629, net12630, net12631, net12632, net12633, net12634, net12635, 
        net12636, net12637, net12638, net12639, net12640, net12641}) );
  ASH_UNS_UNS_OP sll_312 ( .A(div_shl_data), .SH(div_shl_cnta), .Z(div_shl_tmp) );
  dffe_SIZE55 i_div_shl_save ( .din({1'b0, 1'b0, div_shl_tmp}), .en(d3stg_fdiv), .clk(clk), .q(div_shl_save), .se(se), .si({net12534, net12535, net12536, 
        net12537, net12538, net12539, net12540, net12541, net12542, net12543, 
        net12544, net12545, net12546, net12547, net12548, net12549, net12550, 
        net12551, net12552, net12553, net12554, net12555, net12556, net12557, 
        net12558, net12559, net12560, net12561, net12562, net12563, net12564, 
        net12565, net12566, net12567, net12568, net12569, net12570, net12571, 
        net12572, net12573, net12574, net12575, net12576, net12577, net12578, 
        net12579, net12580, net12581, net12582, net12583, net12584, net12585, 
        net12586, net12587, net12588}) );
  dffe_SIZE55 i_div_frac_add_in2 ( .din({d4stg_fdiv, d4stg_fdiv, 
        div_frac_add_in2_in}), .en(div_frac_add_in2_load), .clk(clk), .q(
        div_frac_add_in2), .se(se), .si({net12479, net12480, net12481, 
        net12482, net12483, net12484, net12485, net12486, net12487, net12488, 
        net12489, net12490, net12491, net12492, net12493, net12494, net12495, 
        net12496, net12497, net12498, net12499, net12500, net12501, net12502, 
        net12503, net12504, net12505, net12506, net12507, net12508, net12509, 
        net12510, net12511, net12512, net12513, net12514, net12515, net12516, 
        net12517, net12518, net12519, net12520, net12521, net12522, net12523, 
        net12524, net12525, net12526, net12527, net12528, net12529, net12530, 
        net12531, net12532, net12533}) );
  dffe_SIZE55 i_div_frac_add_in1 ( .din(div_frac_add_in1_in), .en(
        div_frac_add_in1_load), .clk(clk), .q(div_frac_add_in1), .se(se), .si(
        {net12424, net12425, net12426, net12427, net12428, net12429, net12430, 
        net12431, net12432, net12433, net12434, net12435, net12436, net12437, 
        net12438, net12439, net12440, net12441, net12442, net12443, net12444, 
        net12445, net12446, net12447, net12448, net12449, net12450, net12451, 
        net12452, net12453, net12454, net12455, net12456, net12457, net12458, 
        net12459, net12460, net12461, net12462, net12463, net12464, net12465, 
        net12466, net12467, net12468, net12469, net12470, net12471, net12472, 
        net12473, net12474, net12475, net12476, net12477, net12478}) );
  dffe_SIZE55 i_div_frac_add_in1a ( .din(div_frac_add_in1_in), .en(
        div_frac_add_in1_load), .clk(clk), .q(div_frac_add_in1a), .se(se), 
        .si({net12369, net12370, net12371, net12372, net12373, net12374, 
        net12375, net12376, net12377, net12378, net12379, net12380, net12381, 
        net12382, net12383, net12384, net12385, net12386, net12387, net12388, 
        net12389, net12390, net12391, net12392, net12393, net12394, net12395, 
        net12396, net12397, net12398, net12399, net12400, net12401, net12402, 
        net12403, net12404, net12405, net12406, net12407, net12408, net12409, 
        net12410, net12411, net12412, net12413, net12414, net12415, net12416, 
        net12417, net12418, net12419, net12420, net12421, net12422, net12423})
         );
  dffe_SIZE55 i_div_frac_out ( .din(div_frac_out_in), .en(div_frac_out_load), 
        .clk(clk), .q({div_frac_out_54_53, div_frac_out[52], div_frac_outa}), 
        .se(se), .si({net12314, net12315, net12316, net12317, net12318, 
        net12319, net12320, net12321, net12322, net12323, net12324, net12325, 
        net12326, net12327, net12328, net12329, net12330, net12331, net12332, 
        net12333, net12334, net12335, net12336, net12337, net12338, net12339, 
        net12340, net12341, net12342, net12343, net12344, net12345, net12346, 
        net12347, net12348, net12349, net12350, net12351, net12352, net12353, 
        net12354, net12355, net12356, net12357, net12358, net12359, net12360, 
        net12361, net12362, net12363, net12364, net12365, net12366, net12367, 
        net12368}) );
  ADD_UNS_OP add_407 ( .A(div_frac_add_in1a), .B(div_frac_add_in2), .Z({N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  ADD_UNS_OP add_407_2 ( .A({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, 
        N0}), .B(d5stg_fdivb), .Z(div_frac_add) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_NOT I_1 ( .A(N67), .Z(div_norm_inv_in[52]) );
  GTECH_OR2 C337 ( .A(N66), .B(div_norm_qnan), .Z(N67) );
  GTECH_OR2 C338 ( .A(N65), .B(div_norm_inf), .Z(N66) );
  GTECH_OR2 C339 ( .A(N63), .B(N64), .Z(N65) );
  GTECH_OR2 C340 ( .A(N62), .B(div_norm_frac_in2_sng_norm), .Z(N63) );
  GTECH_OR2 C341 ( .A(N60), .B(N61), .Z(N62) );
  GTECH_OR2 C342 ( .A(N59), .B(div_norm_frac_in2_dbl_norm), .Z(N60) );
  GTECH_OR2 C343 ( .A(N57), .B(N58), .Z(N59) );
  GTECH_OR2 C344 ( .A(N56), .B(div_norm_frac_in1_sng_norm), .Z(N57) );
  GTECH_OR2 C345 ( .A(div_norm_frac_in1_dbl_norm), .B(N55), .Z(N56) );
  GTECH_AND2 C346 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[51]), .Z(
        N55) );
  GTECH_AND2 C347 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[54]), .Z(
        N58) );
  GTECH_AND2 C348 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[51]), .Z(
        N61) );
  GTECH_AND2 C349 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[54]), .Z(
        N64) );
  GTECH_NOT I_2 ( .A(N87), .Z(div_norm_inv_in[51]) );
  GTECH_OR2 C351 ( .A(N86), .B(div_norm_qnan), .Z(N87) );
  GTECH_OR2 C352 ( .A(N84), .B(N85), .Z(N86) );
  GTECH_OR2 C353 ( .A(N81), .B(N83), .Z(N84) );
  GTECH_OR2 C354 ( .A(N79), .B(N80), .Z(N81) );
  GTECH_OR2 C355 ( .A(N76), .B(N78), .Z(N79) );
  GTECH_OR2 C356 ( .A(N74), .B(N75), .Z(N76) );
  GTECH_OR2 C357 ( .A(N71), .B(N73), .Z(N74) );
  GTECH_OR2 C358 ( .A(N69), .B(N70), .Z(N71) );
  GTECH_AND2 C359 ( .A(div_norm_frac_in1_dbl_norm), .B(N68), .Z(N69) );
  GTECH_OR2 C360 ( .A(div_frac_in1[51]), .B(d1stg_snan_dbl_in1), .Z(N68) );
  GTECH_AND2 C361 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[50]), .Z(
        N70) );
  GTECH_AND2 C362 ( .A(div_norm_frac_in1_sng_norm), .B(N72), .Z(N73) );
  GTECH_OR2 C363 ( .A(div_frac_in1[54]), .B(d1stg_snan_sng_in1), .Z(N72) );
  GTECH_AND2 C364 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[53]), .Z(
        N75) );
  GTECH_AND2 C365 ( .A(div_norm_frac_in2_dbl_norm), .B(N77), .Z(N78) );
  GTECH_OR2 C366 ( .A(div_frac_in2[51]), .B(d1stg_snan_dbl_in2), .Z(N77) );
  GTECH_AND2 C367 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[50]), .Z(
        N80) );
  GTECH_AND2 C368 ( .A(div_norm_frac_in2_sng_norm), .B(N82), .Z(N83) );
  GTECH_OR2 C369 ( .A(div_frac_in2[54]), .B(d1stg_snan_sng_in2), .Z(N82) );
  GTECH_AND2 C370 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[53]), .Z(
        N85) );
  GTECH_NOT I_3 ( .A(N103), .Z(div_norm_inv_in[50]) );
  GTECH_OR2 C372 ( .A(N102), .B(div_norm_qnan), .Z(N103) );
  GTECH_OR2 C373 ( .A(N100), .B(N101), .Z(N102) );
  GTECH_OR2 C374 ( .A(N98), .B(N99), .Z(N100) );
  GTECH_OR2 C375 ( .A(N96), .B(N97), .Z(N98) );
  GTECH_OR2 C376 ( .A(N94), .B(N95), .Z(N96) );
  GTECH_OR2 C377 ( .A(N92), .B(N93), .Z(N94) );
  GTECH_OR2 C378 ( .A(N90), .B(N91), .Z(N92) );
  GTECH_OR2 C379 ( .A(N88), .B(N89), .Z(N90) );
  GTECH_AND2 C380 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[50]), .Z(
        N88) );
  GTECH_AND2 C381 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[49]), .Z(
        N89) );
  GTECH_AND2 C382 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[53]), .Z(
        N91) );
  GTECH_AND2 C383 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[52]), .Z(
        N93) );
  GTECH_AND2 C384 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[50]), .Z(
        N95) );
  GTECH_AND2 C385 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[49]), .Z(
        N97) );
  GTECH_AND2 C386 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[53]), .Z(
        N99) );
  GTECH_AND2 C387 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[52]), .Z(
        N101) );
  GTECH_NOT I_4 ( .A(N119), .Z(div_norm_inv_in[49]) );
  GTECH_OR2 C389 ( .A(N118), .B(div_norm_qnan), .Z(N119) );
  GTECH_OR2 C390 ( .A(N116), .B(N117), .Z(N118) );
  GTECH_OR2 C391 ( .A(N114), .B(N115), .Z(N116) );
  GTECH_OR2 C392 ( .A(N112), .B(N113), .Z(N114) );
  GTECH_OR2 C393 ( .A(N110), .B(N111), .Z(N112) );
  GTECH_OR2 C394 ( .A(N108), .B(N109), .Z(N110) );
  GTECH_OR2 C395 ( .A(N106), .B(N107), .Z(N108) );
  GTECH_OR2 C396 ( .A(N104), .B(N105), .Z(N106) );
  GTECH_AND2 C397 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[49]), .Z(
        N104) );
  GTECH_AND2 C398 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[48]), .Z(
        N105) );
  GTECH_AND2 C399 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[52]), .Z(
        N107) );
  GTECH_AND2 C400 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[51]), .Z(
        N109) );
  GTECH_AND2 C401 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[49]), .Z(
        N111) );
  GTECH_AND2 C402 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[48]), .Z(
        N113) );
  GTECH_AND2 C403 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[52]), .Z(
        N115) );
  GTECH_AND2 C404 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[51]), .Z(
        N117) );
  GTECH_NOT I_5 ( .A(N135), .Z(div_norm_inv_in[48]) );
  GTECH_OR2 C406 ( .A(N134), .B(div_norm_qnan), .Z(N135) );
  GTECH_OR2 C407 ( .A(N132), .B(N133), .Z(N134) );
  GTECH_OR2 C408 ( .A(N130), .B(N131), .Z(N132) );
  GTECH_OR2 C409 ( .A(N128), .B(N129), .Z(N130) );
  GTECH_OR2 C410 ( .A(N126), .B(N127), .Z(N128) );
  GTECH_OR2 C411 ( .A(N124), .B(N125), .Z(N126) );
  GTECH_OR2 C412 ( .A(N122), .B(N123), .Z(N124) );
  GTECH_OR2 C413 ( .A(N120), .B(N121), .Z(N122) );
  GTECH_AND2 C414 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[48]), .Z(
        N120) );
  GTECH_AND2 C415 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[47]), .Z(
        N121) );
  GTECH_AND2 C416 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[51]), .Z(
        N123) );
  GTECH_AND2 C417 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[50]), .Z(
        N125) );
  GTECH_AND2 C418 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[48]), .Z(
        N127) );
  GTECH_AND2 C419 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[47]), .Z(
        N129) );
  GTECH_AND2 C420 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[51]), .Z(
        N131) );
  GTECH_AND2 C421 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[50]), .Z(
        N133) );
  GTECH_NOT I_6 ( .A(N151), .Z(div_norm_inv_in[47]) );
  GTECH_OR2 C423 ( .A(N150), .B(div_norm_qnan), .Z(N151) );
  GTECH_OR2 C424 ( .A(N148), .B(N149), .Z(N150) );
  GTECH_OR2 C425 ( .A(N146), .B(N147), .Z(N148) );
  GTECH_OR2 C426 ( .A(N144), .B(N145), .Z(N146) );
  GTECH_OR2 C427 ( .A(N142), .B(N143), .Z(N144) );
  GTECH_OR2 C428 ( .A(N140), .B(N141), .Z(N142) );
  GTECH_OR2 C429 ( .A(N138), .B(N139), .Z(N140) );
  GTECH_OR2 C430 ( .A(N136), .B(N137), .Z(N138) );
  GTECH_AND2 C431 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[47]), .Z(
        N136) );
  GTECH_AND2 C432 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[46]), .Z(
        N137) );
  GTECH_AND2 C433 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[50]), .Z(
        N139) );
  GTECH_AND2 C434 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[49]), .Z(
        N141) );
  GTECH_AND2 C435 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[47]), .Z(
        N143) );
  GTECH_AND2 C436 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[46]), .Z(
        N145) );
  GTECH_AND2 C437 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[50]), .Z(
        N147) );
  GTECH_AND2 C438 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[49]), .Z(
        N149) );
  GTECH_NOT I_7 ( .A(N167), .Z(div_norm_inv_in[46]) );
  GTECH_OR2 C440 ( .A(N166), .B(div_norm_qnan), .Z(N167) );
  GTECH_OR2 C441 ( .A(N164), .B(N165), .Z(N166) );
  GTECH_OR2 C442 ( .A(N162), .B(N163), .Z(N164) );
  GTECH_OR2 C443 ( .A(N160), .B(N161), .Z(N162) );
  GTECH_OR2 C444 ( .A(N158), .B(N159), .Z(N160) );
  GTECH_OR2 C445 ( .A(N156), .B(N157), .Z(N158) );
  GTECH_OR2 C446 ( .A(N154), .B(N155), .Z(N156) );
  GTECH_OR2 C447 ( .A(N152), .B(N153), .Z(N154) );
  GTECH_AND2 C448 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[46]), .Z(
        N152) );
  GTECH_AND2 C449 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[45]), .Z(
        N153) );
  GTECH_AND2 C450 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[49]), .Z(
        N155) );
  GTECH_AND2 C451 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[48]), .Z(
        N157) );
  GTECH_AND2 C452 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[46]), .Z(
        N159) );
  GTECH_AND2 C453 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[45]), .Z(
        N161) );
  GTECH_AND2 C454 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[49]), .Z(
        N163) );
  GTECH_AND2 C455 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[48]), .Z(
        N165) );
  GTECH_NOT I_8 ( .A(N183), .Z(div_norm_inv_in[45]) );
  GTECH_OR2 C457 ( .A(N182), .B(div_norm_qnan), .Z(N183) );
  GTECH_OR2 C458 ( .A(N180), .B(N181), .Z(N182) );
  GTECH_OR2 C459 ( .A(N178), .B(N179), .Z(N180) );
  GTECH_OR2 C460 ( .A(N176), .B(N177), .Z(N178) );
  GTECH_OR2 C461 ( .A(N174), .B(N175), .Z(N176) );
  GTECH_OR2 C462 ( .A(N172), .B(N173), .Z(N174) );
  GTECH_OR2 C463 ( .A(N170), .B(N171), .Z(N172) );
  GTECH_OR2 C464 ( .A(N168), .B(N169), .Z(N170) );
  GTECH_AND2 C465 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[45]), .Z(
        N168) );
  GTECH_AND2 C466 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[44]), .Z(
        N169) );
  GTECH_AND2 C467 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[48]), .Z(
        N171) );
  GTECH_AND2 C468 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[47]), .Z(
        N173) );
  GTECH_AND2 C469 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[45]), .Z(
        N175) );
  GTECH_AND2 C470 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[44]), .Z(
        N177) );
  GTECH_AND2 C471 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[48]), .Z(
        N179) );
  GTECH_AND2 C472 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[47]), .Z(
        N181) );
  GTECH_NOT I_9 ( .A(N199), .Z(div_norm_inv_in[44]) );
  GTECH_OR2 C474 ( .A(N198), .B(div_norm_qnan), .Z(N199) );
  GTECH_OR2 C475 ( .A(N196), .B(N197), .Z(N198) );
  GTECH_OR2 C476 ( .A(N194), .B(N195), .Z(N196) );
  GTECH_OR2 C477 ( .A(N192), .B(N193), .Z(N194) );
  GTECH_OR2 C478 ( .A(N190), .B(N191), .Z(N192) );
  GTECH_OR2 C479 ( .A(N188), .B(N189), .Z(N190) );
  GTECH_OR2 C480 ( .A(N186), .B(N187), .Z(N188) );
  GTECH_OR2 C481 ( .A(N184), .B(N185), .Z(N186) );
  GTECH_AND2 C482 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[44]), .Z(
        N184) );
  GTECH_AND2 C483 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[43]), .Z(
        N185) );
  GTECH_AND2 C484 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[47]), .Z(
        N187) );
  GTECH_AND2 C485 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[46]), .Z(
        N189) );
  GTECH_AND2 C486 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[44]), .Z(
        N191) );
  GTECH_AND2 C487 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[43]), .Z(
        N193) );
  GTECH_AND2 C488 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[47]), .Z(
        N195) );
  GTECH_AND2 C489 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[46]), .Z(
        N197) );
  GTECH_NOT I_10 ( .A(N215), .Z(div_norm_inv_in[43]) );
  GTECH_OR2 C491 ( .A(N214), .B(div_norm_qnan), .Z(N215) );
  GTECH_OR2 C492 ( .A(N212), .B(N213), .Z(N214) );
  GTECH_OR2 C493 ( .A(N210), .B(N211), .Z(N212) );
  GTECH_OR2 C494 ( .A(N208), .B(N209), .Z(N210) );
  GTECH_OR2 C495 ( .A(N206), .B(N207), .Z(N208) );
  GTECH_OR2 C496 ( .A(N204), .B(N205), .Z(N206) );
  GTECH_OR2 C497 ( .A(N202), .B(N203), .Z(N204) );
  GTECH_OR2 C498 ( .A(N200), .B(N201), .Z(N202) );
  GTECH_AND2 C499 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[43]), .Z(
        N200) );
  GTECH_AND2 C500 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[42]), .Z(
        N201) );
  GTECH_AND2 C501 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[46]), .Z(
        N203) );
  GTECH_AND2 C502 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[45]), .Z(
        N205) );
  GTECH_AND2 C503 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[43]), .Z(
        N207) );
  GTECH_AND2 C504 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[42]), .Z(
        N209) );
  GTECH_AND2 C505 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[46]), .Z(
        N211) );
  GTECH_AND2 C506 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[45]), .Z(
        N213) );
  GTECH_NOT I_11 ( .A(N231), .Z(div_norm_inv_in[42]) );
  GTECH_OR2 C508 ( .A(N230), .B(div_norm_qnan), .Z(N231) );
  GTECH_OR2 C509 ( .A(N228), .B(N229), .Z(N230) );
  GTECH_OR2 C510 ( .A(N226), .B(N227), .Z(N228) );
  GTECH_OR2 C511 ( .A(N224), .B(N225), .Z(N226) );
  GTECH_OR2 C512 ( .A(N222), .B(N223), .Z(N224) );
  GTECH_OR2 C513 ( .A(N220), .B(N221), .Z(N222) );
  GTECH_OR2 C514 ( .A(N218), .B(N219), .Z(N220) );
  GTECH_OR2 C515 ( .A(N216), .B(N217), .Z(N218) );
  GTECH_AND2 C516 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[42]), .Z(
        N216) );
  GTECH_AND2 C517 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[41]), .Z(
        N217) );
  GTECH_AND2 C518 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[45]), .Z(
        N219) );
  GTECH_AND2 C519 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[44]), .Z(
        N221) );
  GTECH_AND2 C520 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[42]), .Z(
        N223) );
  GTECH_AND2 C521 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[41]), .Z(
        N225) );
  GTECH_AND2 C522 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[45]), .Z(
        N227) );
  GTECH_AND2 C523 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[44]), .Z(
        N229) );
  GTECH_NOT I_12 ( .A(N247), .Z(div_norm_inv_in[41]) );
  GTECH_OR2 C525 ( .A(N246), .B(div_norm_qnan), .Z(N247) );
  GTECH_OR2 C526 ( .A(N244), .B(N245), .Z(N246) );
  GTECH_OR2 C527 ( .A(N242), .B(N243), .Z(N244) );
  GTECH_OR2 C528 ( .A(N240), .B(N241), .Z(N242) );
  GTECH_OR2 C529 ( .A(N238), .B(N239), .Z(N240) );
  GTECH_OR2 C530 ( .A(N236), .B(N237), .Z(N238) );
  GTECH_OR2 C531 ( .A(N234), .B(N235), .Z(N236) );
  GTECH_OR2 C532 ( .A(N232), .B(N233), .Z(N234) );
  GTECH_AND2 C533 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[41]), .Z(
        N232) );
  GTECH_AND2 C534 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[40]), .Z(
        N233) );
  GTECH_AND2 C535 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[44]), .Z(
        N235) );
  GTECH_AND2 C536 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[43]), .Z(
        N237) );
  GTECH_AND2 C537 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[41]), .Z(
        N239) );
  GTECH_AND2 C538 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[40]), .Z(
        N241) );
  GTECH_AND2 C539 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[44]), .Z(
        N243) );
  GTECH_AND2 C540 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[43]), .Z(
        N245) );
  GTECH_NOT I_13 ( .A(N263), .Z(div_norm_inv_in[40]) );
  GTECH_OR2 C542 ( .A(N262), .B(div_norm_qnan), .Z(N263) );
  GTECH_OR2 C543 ( .A(N260), .B(N261), .Z(N262) );
  GTECH_OR2 C544 ( .A(N258), .B(N259), .Z(N260) );
  GTECH_OR2 C545 ( .A(N256), .B(N257), .Z(N258) );
  GTECH_OR2 C546 ( .A(N254), .B(N255), .Z(N256) );
  GTECH_OR2 C547 ( .A(N252), .B(N253), .Z(N254) );
  GTECH_OR2 C548 ( .A(N250), .B(N251), .Z(N252) );
  GTECH_OR2 C549 ( .A(N248), .B(N249), .Z(N250) );
  GTECH_AND2 C550 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[40]), .Z(
        N248) );
  GTECH_AND2 C551 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[39]), .Z(
        N249) );
  GTECH_AND2 C552 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[43]), .Z(
        N251) );
  GTECH_AND2 C553 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[42]), .Z(
        N253) );
  GTECH_AND2 C554 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[40]), .Z(
        N255) );
  GTECH_AND2 C555 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[39]), .Z(
        N257) );
  GTECH_AND2 C556 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[43]), .Z(
        N259) );
  GTECH_AND2 C557 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[42]), .Z(
        N261) );
  GTECH_NOT I_14 ( .A(N279), .Z(div_norm_inv_in[39]) );
  GTECH_OR2 C559 ( .A(N278), .B(div_norm_qnan), .Z(N279) );
  GTECH_OR2 C560 ( .A(N276), .B(N277), .Z(N278) );
  GTECH_OR2 C561 ( .A(N274), .B(N275), .Z(N276) );
  GTECH_OR2 C562 ( .A(N272), .B(N273), .Z(N274) );
  GTECH_OR2 C563 ( .A(N270), .B(N271), .Z(N272) );
  GTECH_OR2 C564 ( .A(N268), .B(N269), .Z(N270) );
  GTECH_OR2 C565 ( .A(N266), .B(N267), .Z(N268) );
  GTECH_OR2 C566 ( .A(N264), .B(N265), .Z(N266) );
  GTECH_AND2 C567 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[39]), .Z(
        N264) );
  GTECH_AND2 C568 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[38]), .Z(
        N265) );
  GTECH_AND2 C569 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[42]), .Z(
        N267) );
  GTECH_AND2 C570 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[41]), .Z(
        N269) );
  GTECH_AND2 C571 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[39]), .Z(
        N271) );
  GTECH_AND2 C572 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[38]), .Z(
        N273) );
  GTECH_AND2 C573 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[42]), .Z(
        N275) );
  GTECH_AND2 C574 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[41]), .Z(
        N277) );
  GTECH_NOT I_15 ( .A(N295), .Z(div_norm_inv_in[38]) );
  GTECH_OR2 C576 ( .A(N294), .B(div_norm_qnan), .Z(N295) );
  GTECH_OR2 C577 ( .A(N292), .B(N293), .Z(N294) );
  GTECH_OR2 C578 ( .A(N290), .B(N291), .Z(N292) );
  GTECH_OR2 C579 ( .A(N288), .B(N289), .Z(N290) );
  GTECH_OR2 C580 ( .A(N286), .B(N287), .Z(N288) );
  GTECH_OR2 C581 ( .A(N284), .B(N285), .Z(N286) );
  GTECH_OR2 C582 ( .A(N282), .B(N283), .Z(N284) );
  GTECH_OR2 C583 ( .A(N280), .B(N281), .Z(N282) );
  GTECH_AND2 C584 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[38]), .Z(
        N280) );
  GTECH_AND2 C585 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[37]), .Z(
        N281) );
  GTECH_AND2 C586 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[41]), .Z(
        N283) );
  GTECH_AND2 C587 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[40]), .Z(
        N285) );
  GTECH_AND2 C588 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[38]), .Z(
        N287) );
  GTECH_AND2 C589 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[37]), .Z(
        N289) );
  GTECH_AND2 C590 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[41]), .Z(
        N291) );
  GTECH_AND2 C591 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[40]), .Z(
        N293) );
  GTECH_NOT I_16 ( .A(N311), .Z(div_norm_inv_in[37]) );
  GTECH_OR2 C593 ( .A(N310), .B(div_norm_qnan), .Z(N311) );
  GTECH_OR2 C594 ( .A(N308), .B(N309), .Z(N310) );
  GTECH_OR2 C595 ( .A(N306), .B(N307), .Z(N308) );
  GTECH_OR2 C596 ( .A(N304), .B(N305), .Z(N306) );
  GTECH_OR2 C597 ( .A(N302), .B(N303), .Z(N304) );
  GTECH_OR2 C598 ( .A(N300), .B(N301), .Z(N302) );
  GTECH_OR2 C599 ( .A(N298), .B(N299), .Z(N300) );
  GTECH_OR2 C600 ( .A(N296), .B(N297), .Z(N298) );
  GTECH_AND2 C601 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[37]), .Z(
        N296) );
  GTECH_AND2 C602 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[36]), .Z(
        N297) );
  GTECH_AND2 C603 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[40]), .Z(
        N299) );
  GTECH_AND2 C604 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[39]), .Z(
        N301) );
  GTECH_AND2 C605 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[37]), .Z(
        N303) );
  GTECH_AND2 C606 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[36]), .Z(
        N305) );
  GTECH_AND2 C607 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[40]), .Z(
        N307) );
  GTECH_AND2 C608 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[39]), .Z(
        N309) );
  GTECH_NOT I_17 ( .A(N327), .Z(div_norm_inv_in[36]) );
  GTECH_OR2 C610 ( .A(N326), .B(div_norm_qnan), .Z(N327) );
  GTECH_OR2 C611 ( .A(N324), .B(N325), .Z(N326) );
  GTECH_OR2 C612 ( .A(N322), .B(N323), .Z(N324) );
  GTECH_OR2 C613 ( .A(N320), .B(N321), .Z(N322) );
  GTECH_OR2 C614 ( .A(N318), .B(N319), .Z(N320) );
  GTECH_OR2 C615 ( .A(N316), .B(N317), .Z(N318) );
  GTECH_OR2 C616 ( .A(N314), .B(N315), .Z(N316) );
  GTECH_OR2 C617 ( .A(N312), .B(N313), .Z(N314) );
  GTECH_AND2 C618 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[36]), .Z(
        N312) );
  GTECH_AND2 C619 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[35]), .Z(
        N313) );
  GTECH_AND2 C620 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[39]), .Z(
        N315) );
  GTECH_AND2 C621 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[38]), .Z(
        N317) );
  GTECH_AND2 C622 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[36]), .Z(
        N319) );
  GTECH_AND2 C623 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[35]), .Z(
        N321) );
  GTECH_AND2 C624 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[39]), .Z(
        N323) );
  GTECH_AND2 C625 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[38]), .Z(
        N325) );
  GTECH_NOT I_18 ( .A(N343), .Z(div_norm_inv_in[35]) );
  GTECH_OR2 C627 ( .A(N342), .B(div_norm_qnan), .Z(N343) );
  GTECH_OR2 C628 ( .A(N340), .B(N341), .Z(N342) );
  GTECH_OR2 C629 ( .A(N338), .B(N339), .Z(N340) );
  GTECH_OR2 C630 ( .A(N336), .B(N337), .Z(N338) );
  GTECH_OR2 C631 ( .A(N334), .B(N335), .Z(N336) );
  GTECH_OR2 C632 ( .A(N332), .B(N333), .Z(N334) );
  GTECH_OR2 C633 ( .A(N330), .B(N331), .Z(N332) );
  GTECH_OR2 C634 ( .A(N328), .B(N329), .Z(N330) );
  GTECH_AND2 C635 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[35]), .Z(
        N328) );
  GTECH_AND2 C636 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[34]), .Z(
        N329) );
  GTECH_AND2 C637 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[38]), .Z(
        N331) );
  GTECH_AND2 C638 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[37]), .Z(
        N333) );
  GTECH_AND2 C639 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[35]), .Z(
        N335) );
  GTECH_AND2 C640 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[34]), .Z(
        N337) );
  GTECH_AND2 C641 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[38]), .Z(
        N339) );
  GTECH_AND2 C642 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[37]), .Z(
        N341) );
  GTECH_NOT I_19 ( .A(N359), .Z(div_norm_inv_in[34]) );
  GTECH_OR2 C644 ( .A(N358), .B(div_norm_qnan), .Z(N359) );
  GTECH_OR2 C645 ( .A(N356), .B(N357), .Z(N358) );
  GTECH_OR2 C646 ( .A(N354), .B(N355), .Z(N356) );
  GTECH_OR2 C647 ( .A(N352), .B(N353), .Z(N354) );
  GTECH_OR2 C648 ( .A(N350), .B(N351), .Z(N352) );
  GTECH_OR2 C649 ( .A(N348), .B(N349), .Z(N350) );
  GTECH_OR2 C650 ( .A(N346), .B(N347), .Z(N348) );
  GTECH_OR2 C651 ( .A(N344), .B(N345), .Z(N346) );
  GTECH_AND2 C652 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[34]), .Z(
        N344) );
  GTECH_AND2 C653 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[33]), .Z(
        N345) );
  GTECH_AND2 C654 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[37]), .Z(
        N347) );
  GTECH_AND2 C655 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[36]), .Z(
        N349) );
  GTECH_AND2 C656 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[34]), .Z(
        N351) );
  GTECH_AND2 C657 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[33]), .Z(
        N353) );
  GTECH_AND2 C658 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[37]), .Z(
        N355) );
  GTECH_AND2 C659 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[36]), .Z(
        N357) );
  GTECH_NOT I_20 ( .A(N375), .Z(div_norm_inv_in[33]) );
  GTECH_OR2 C661 ( .A(N374), .B(div_norm_qnan), .Z(N375) );
  GTECH_OR2 C662 ( .A(N372), .B(N373), .Z(N374) );
  GTECH_OR2 C663 ( .A(N370), .B(N371), .Z(N372) );
  GTECH_OR2 C664 ( .A(N368), .B(N369), .Z(N370) );
  GTECH_OR2 C665 ( .A(N366), .B(N367), .Z(N368) );
  GTECH_OR2 C666 ( .A(N364), .B(N365), .Z(N366) );
  GTECH_OR2 C667 ( .A(N362), .B(N363), .Z(N364) );
  GTECH_OR2 C668 ( .A(N360), .B(N361), .Z(N362) );
  GTECH_AND2 C669 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[33]), .Z(
        N360) );
  GTECH_AND2 C670 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[32]), .Z(
        N361) );
  GTECH_AND2 C671 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[36]), .Z(
        N363) );
  GTECH_AND2 C672 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[35]), .Z(
        N365) );
  GTECH_AND2 C673 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[33]), .Z(
        N367) );
  GTECH_AND2 C674 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[32]), .Z(
        N369) );
  GTECH_AND2 C675 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[36]), .Z(
        N371) );
  GTECH_AND2 C676 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[35]), .Z(
        N373) );
  GTECH_NOT I_21 ( .A(N391), .Z(div_norm_inv_in[32]) );
  GTECH_OR2 C678 ( .A(N390), .B(div_norm_qnan), .Z(N391) );
  GTECH_OR2 C679 ( .A(N388), .B(N389), .Z(N390) );
  GTECH_OR2 C680 ( .A(N386), .B(N387), .Z(N388) );
  GTECH_OR2 C681 ( .A(N384), .B(N385), .Z(N386) );
  GTECH_OR2 C682 ( .A(N382), .B(N383), .Z(N384) );
  GTECH_OR2 C683 ( .A(N380), .B(N381), .Z(N382) );
  GTECH_OR2 C684 ( .A(N378), .B(N379), .Z(N380) );
  GTECH_OR2 C685 ( .A(N376), .B(N377), .Z(N378) );
  GTECH_AND2 C686 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[32]), .Z(
        N376) );
  GTECH_AND2 C687 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[31]), .Z(
        N377) );
  GTECH_AND2 C688 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[35]), .Z(
        N379) );
  GTECH_AND2 C689 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[34]), .Z(
        N381) );
  GTECH_AND2 C690 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[32]), .Z(
        N383) );
  GTECH_AND2 C691 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[31]), .Z(
        N385) );
  GTECH_AND2 C692 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[35]), .Z(
        N387) );
  GTECH_AND2 C693 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[34]), .Z(
        N389) );
  GTECH_NOT I_22 ( .A(N407), .Z(div_norm_inv_in[31]) );
  GTECH_OR2 C695 ( .A(N406), .B(div_norm_qnan), .Z(N407) );
  GTECH_OR2 C696 ( .A(N404), .B(N405), .Z(N406) );
  GTECH_OR2 C697 ( .A(N402), .B(N403), .Z(N404) );
  GTECH_OR2 C698 ( .A(N400), .B(N401), .Z(N402) );
  GTECH_OR2 C699 ( .A(N398), .B(N399), .Z(N400) );
  GTECH_OR2 C700 ( .A(N396), .B(N397), .Z(N398) );
  GTECH_OR2 C701 ( .A(N394), .B(N395), .Z(N396) );
  GTECH_OR2 C702 ( .A(N392), .B(N393), .Z(N394) );
  GTECH_AND2 C703 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[31]), .Z(
        N392) );
  GTECH_AND2 C704 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[30]), .Z(
        N393) );
  GTECH_AND2 C705 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[34]), .Z(
        N395) );
  GTECH_AND2 C706 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[33]), .Z(
        N397) );
  GTECH_AND2 C707 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[31]), .Z(
        N399) );
  GTECH_AND2 C708 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[30]), .Z(
        N401) );
  GTECH_AND2 C709 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[34]), .Z(
        N403) );
  GTECH_AND2 C710 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[33]), .Z(
        N405) );
  GTECH_NOT I_23 ( .A(N423), .Z(div_norm_inv_in[30]) );
  GTECH_OR2 C712 ( .A(N422), .B(div_norm_qnan), .Z(N423) );
  GTECH_OR2 C713 ( .A(N420), .B(N421), .Z(N422) );
  GTECH_OR2 C714 ( .A(N418), .B(N419), .Z(N420) );
  GTECH_OR2 C715 ( .A(N416), .B(N417), .Z(N418) );
  GTECH_OR2 C716 ( .A(N414), .B(N415), .Z(N416) );
  GTECH_OR2 C717 ( .A(N412), .B(N413), .Z(N414) );
  GTECH_OR2 C718 ( .A(N410), .B(N411), .Z(N412) );
  GTECH_OR2 C719 ( .A(N408), .B(N409), .Z(N410) );
  GTECH_AND2 C720 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[30]), .Z(
        N408) );
  GTECH_AND2 C721 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[29]), .Z(
        N409) );
  GTECH_AND2 C722 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[33]), .Z(
        N411) );
  GTECH_AND2 C723 ( .A(div_norm_frac_in1_sng_dnrm), .B(div_frac_in1[32]), .Z(
        N413) );
  GTECH_AND2 C724 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[30]), .Z(
        N415) );
  GTECH_AND2 C725 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[29]), .Z(
        N417) );
  GTECH_AND2 C726 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[33]), .Z(
        N419) );
  GTECH_AND2 C727 ( .A(div_norm_frac_in2_sng_dnrm), .B(div_frac_in2[32]), .Z(
        N421) );
  GTECH_NOT I_24 ( .A(N435), .Z(div_norm_inv_in[29]) );
  GTECH_OR2 C729 ( .A(N434), .B(div_norm_qnan), .Z(N435) );
  GTECH_OR2 C730 ( .A(N432), .B(N433), .Z(N434) );
  GTECH_OR2 C731 ( .A(N430), .B(N431), .Z(N432) );
  GTECH_OR2 C732 ( .A(N428), .B(N429), .Z(N430) );
  GTECH_OR2 C733 ( .A(N426), .B(N427), .Z(N428) );
  GTECH_OR2 C734 ( .A(N424), .B(N425), .Z(N426) );
  GTECH_AND2 C735 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[29]), .Z(
        N424) );
  GTECH_AND2 C736 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[28]), .Z(
        N425) );
  GTECH_AND2 C737 ( .A(div_norm_frac_in1_sng_norm), .B(div_frac_in1[32]), .Z(
        N427) );
  GTECH_AND2 C738 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[29]), .Z(
        N429) );
  GTECH_AND2 C739 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[28]), .Z(
        N431) );
  GTECH_AND2 C740 ( .A(div_norm_frac_in2_sng_norm), .B(div_frac_in2[32]), .Z(
        N433) );
  GTECH_NOT I_25 ( .A(N444), .Z(div_norm_inv_in[28]) );
  GTECH_OR2 C742 ( .A(N442), .B(N443), .Z(N444) );
  GTECH_OR2 C743 ( .A(N440), .B(N441), .Z(N442) );
  GTECH_OR2 C744 ( .A(N438), .B(N439), .Z(N440) );
  GTECH_OR2 C745 ( .A(N436), .B(N437), .Z(N438) );
  GTECH_AND2 C746 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[28]), .Z(
        N436) );
  GTECH_AND2 C747 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[27]), .Z(
        N437) );
  GTECH_AND2 C748 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[28]), .Z(
        N439) );
  GTECH_AND2 C749 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[27]), .Z(
        N441) );
  GTECH_AND2 C750 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N443) );
  GTECH_NOT I_26 ( .A(N453), .Z(div_norm_inv_in[27]) );
  GTECH_OR2 C752 ( .A(N451), .B(N452), .Z(N453) );
  GTECH_OR2 C753 ( .A(N449), .B(N450), .Z(N451) );
  GTECH_OR2 C754 ( .A(N447), .B(N448), .Z(N449) );
  GTECH_OR2 C755 ( .A(N445), .B(N446), .Z(N447) );
  GTECH_AND2 C756 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[27]), .Z(
        N445) );
  GTECH_AND2 C757 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[26]), .Z(
        N446) );
  GTECH_AND2 C758 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[27]), .Z(
        N448) );
  GTECH_AND2 C759 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[26]), .Z(
        N450) );
  GTECH_AND2 C760 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N452) );
  GTECH_NOT I_27 ( .A(N462), .Z(div_norm_inv_in[26]) );
  GTECH_OR2 C762 ( .A(N460), .B(N461), .Z(N462) );
  GTECH_OR2 C763 ( .A(N458), .B(N459), .Z(N460) );
  GTECH_OR2 C764 ( .A(N456), .B(N457), .Z(N458) );
  GTECH_OR2 C765 ( .A(N454), .B(N455), .Z(N456) );
  GTECH_AND2 C766 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[26]), .Z(
        N454) );
  GTECH_AND2 C767 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[25]), .Z(
        N455) );
  GTECH_AND2 C768 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[26]), .Z(
        N457) );
  GTECH_AND2 C769 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[25]), .Z(
        N459) );
  GTECH_AND2 C770 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N461) );
  GTECH_NOT I_28 ( .A(N471), .Z(div_norm_inv_in[25]) );
  GTECH_OR2 C772 ( .A(N469), .B(N470), .Z(N471) );
  GTECH_OR2 C773 ( .A(N467), .B(N468), .Z(N469) );
  GTECH_OR2 C774 ( .A(N465), .B(N466), .Z(N467) );
  GTECH_OR2 C775 ( .A(N463), .B(N464), .Z(N465) );
  GTECH_AND2 C776 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[25]), .Z(
        N463) );
  GTECH_AND2 C777 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[24]), .Z(
        N464) );
  GTECH_AND2 C778 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[25]), .Z(
        N466) );
  GTECH_AND2 C779 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[24]), .Z(
        N468) );
  GTECH_AND2 C780 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N470) );
  GTECH_NOT I_29 ( .A(N480), .Z(div_norm_inv_in[24]) );
  GTECH_OR2 C782 ( .A(N478), .B(N479), .Z(N480) );
  GTECH_OR2 C783 ( .A(N476), .B(N477), .Z(N478) );
  GTECH_OR2 C784 ( .A(N474), .B(N475), .Z(N476) );
  GTECH_OR2 C785 ( .A(N472), .B(N473), .Z(N474) );
  GTECH_AND2 C786 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[24]), .Z(
        N472) );
  GTECH_AND2 C787 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[23]), .Z(
        N473) );
  GTECH_AND2 C788 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[24]), .Z(
        N475) );
  GTECH_AND2 C789 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[23]), .Z(
        N477) );
  GTECH_AND2 C790 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N479) );
  GTECH_NOT I_30 ( .A(N489), .Z(div_norm_inv_in[23]) );
  GTECH_OR2 C792 ( .A(N487), .B(N488), .Z(N489) );
  GTECH_OR2 C793 ( .A(N485), .B(N486), .Z(N487) );
  GTECH_OR2 C794 ( .A(N483), .B(N484), .Z(N485) );
  GTECH_OR2 C795 ( .A(N481), .B(N482), .Z(N483) );
  GTECH_AND2 C796 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[23]), .Z(
        N481) );
  GTECH_AND2 C797 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[22]), .Z(
        N482) );
  GTECH_AND2 C798 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[23]), .Z(
        N484) );
  GTECH_AND2 C799 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[22]), .Z(
        N486) );
  GTECH_AND2 C800 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N488) );
  GTECH_NOT I_31 ( .A(N498), .Z(div_norm_inv_in[22]) );
  GTECH_OR2 C802 ( .A(N496), .B(N497), .Z(N498) );
  GTECH_OR2 C803 ( .A(N494), .B(N495), .Z(N496) );
  GTECH_OR2 C804 ( .A(N492), .B(N493), .Z(N494) );
  GTECH_OR2 C805 ( .A(N490), .B(N491), .Z(N492) );
  GTECH_AND2 C806 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[22]), .Z(
        N490) );
  GTECH_AND2 C807 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[21]), .Z(
        N491) );
  GTECH_AND2 C808 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[22]), .Z(
        N493) );
  GTECH_AND2 C809 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[21]), .Z(
        N495) );
  GTECH_AND2 C810 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N497) );
  GTECH_NOT I_32 ( .A(N507), .Z(div_norm_inv_in[21]) );
  GTECH_OR2 C812 ( .A(N505), .B(N506), .Z(N507) );
  GTECH_OR2 C813 ( .A(N503), .B(N504), .Z(N505) );
  GTECH_OR2 C814 ( .A(N501), .B(N502), .Z(N503) );
  GTECH_OR2 C815 ( .A(N499), .B(N500), .Z(N501) );
  GTECH_AND2 C816 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[21]), .Z(
        N499) );
  GTECH_AND2 C817 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[20]), .Z(
        N500) );
  GTECH_AND2 C818 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[21]), .Z(
        N502) );
  GTECH_AND2 C819 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[20]), .Z(
        N504) );
  GTECH_AND2 C820 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N506) );
  GTECH_NOT I_33 ( .A(N516), .Z(div_norm_inv_in[20]) );
  GTECH_OR2 C822 ( .A(N514), .B(N515), .Z(N516) );
  GTECH_OR2 C823 ( .A(N512), .B(N513), .Z(N514) );
  GTECH_OR2 C824 ( .A(N510), .B(N511), .Z(N512) );
  GTECH_OR2 C825 ( .A(N508), .B(N509), .Z(N510) );
  GTECH_AND2 C826 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[20]), .Z(
        N508) );
  GTECH_AND2 C827 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[19]), .Z(
        N509) );
  GTECH_AND2 C828 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[20]), .Z(
        N511) );
  GTECH_AND2 C829 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[19]), .Z(
        N513) );
  GTECH_AND2 C830 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N515) );
  GTECH_NOT I_34 ( .A(N525), .Z(div_norm_inv_in[19]) );
  GTECH_OR2 C832 ( .A(N523), .B(N524), .Z(N525) );
  GTECH_OR2 C833 ( .A(N521), .B(N522), .Z(N523) );
  GTECH_OR2 C834 ( .A(N519), .B(N520), .Z(N521) );
  GTECH_OR2 C835 ( .A(N517), .B(N518), .Z(N519) );
  GTECH_AND2 C836 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[19]), .Z(
        N517) );
  GTECH_AND2 C837 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[18]), .Z(
        N518) );
  GTECH_AND2 C838 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[19]), .Z(
        N520) );
  GTECH_AND2 C839 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[18]), .Z(
        N522) );
  GTECH_AND2 C840 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N524) );
  GTECH_NOT I_35 ( .A(N534), .Z(div_norm_inv_in[18]) );
  GTECH_OR2 C842 ( .A(N532), .B(N533), .Z(N534) );
  GTECH_OR2 C843 ( .A(N530), .B(N531), .Z(N532) );
  GTECH_OR2 C844 ( .A(N528), .B(N529), .Z(N530) );
  GTECH_OR2 C845 ( .A(N526), .B(N527), .Z(N528) );
  GTECH_AND2 C846 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[18]), .Z(
        N526) );
  GTECH_AND2 C847 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[17]), .Z(
        N527) );
  GTECH_AND2 C848 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[18]), .Z(
        N529) );
  GTECH_AND2 C849 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[17]), .Z(
        N531) );
  GTECH_AND2 C850 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N533) );
  GTECH_NOT I_36 ( .A(N543), .Z(div_norm_inv_in[17]) );
  GTECH_OR2 C852 ( .A(N541), .B(N542), .Z(N543) );
  GTECH_OR2 C853 ( .A(N539), .B(N540), .Z(N541) );
  GTECH_OR2 C854 ( .A(N537), .B(N538), .Z(N539) );
  GTECH_OR2 C855 ( .A(N535), .B(N536), .Z(N537) );
  GTECH_AND2 C856 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[17]), .Z(
        N535) );
  GTECH_AND2 C857 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[16]), .Z(
        N536) );
  GTECH_AND2 C858 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[17]), .Z(
        N538) );
  GTECH_AND2 C859 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[16]), .Z(
        N540) );
  GTECH_AND2 C860 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N542) );
  GTECH_NOT I_37 ( .A(N552), .Z(div_norm_inv_in[16]) );
  GTECH_OR2 C862 ( .A(N550), .B(N551), .Z(N552) );
  GTECH_OR2 C863 ( .A(N548), .B(N549), .Z(N550) );
  GTECH_OR2 C864 ( .A(N546), .B(N547), .Z(N548) );
  GTECH_OR2 C865 ( .A(N544), .B(N545), .Z(N546) );
  GTECH_AND2 C866 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[16]), .Z(
        N544) );
  GTECH_AND2 C867 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[15]), .Z(
        N545) );
  GTECH_AND2 C868 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[16]), .Z(
        N547) );
  GTECH_AND2 C869 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[15]), .Z(
        N549) );
  GTECH_AND2 C870 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N551) );
  GTECH_NOT I_38 ( .A(N561), .Z(div_norm_inv_in[15]) );
  GTECH_OR2 C872 ( .A(N559), .B(N560), .Z(N561) );
  GTECH_OR2 C873 ( .A(N557), .B(N558), .Z(N559) );
  GTECH_OR2 C874 ( .A(N555), .B(N556), .Z(N557) );
  GTECH_OR2 C875 ( .A(N553), .B(N554), .Z(N555) );
  GTECH_AND2 C876 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[15]), .Z(
        N553) );
  GTECH_AND2 C877 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[14]), .Z(
        N554) );
  GTECH_AND2 C878 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[15]), .Z(
        N556) );
  GTECH_AND2 C879 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[14]), .Z(
        N558) );
  GTECH_AND2 C880 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N560) );
  GTECH_NOT I_39 ( .A(N570), .Z(div_norm_inv_in[14]) );
  GTECH_OR2 C882 ( .A(N568), .B(N569), .Z(N570) );
  GTECH_OR2 C883 ( .A(N566), .B(N567), .Z(N568) );
  GTECH_OR2 C884 ( .A(N564), .B(N565), .Z(N566) );
  GTECH_OR2 C885 ( .A(N562), .B(N563), .Z(N564) );
  GTECH_AND2 C886 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[14]), .Z(
        N562) );
  GTECH_AND2 C887 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[13]), .Z(
        N563) );
  GTECH_AND2 C888 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[14]), .Z(
        N565) );
  GTECH_AND2 C889 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[13]), .Z(
        N567) );
  GTECH_AND2 C890 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N569) );
  GTECH_NOT I_40 ( .A(N579), .Z(div_norm_inv_in[13]) );
  GTECH_OR2 C892 ( .A(N577), .B(N578), .Z(N579) );
  GTECH_OR2 C893 ( .A(N575), .B(N576), .Z(N577) );
  GTECH_OR2 C894 ( .A(N573), .B(N574), .Z(N575) );
  GTECH_OR2 C895 ( .A(N571), .B(N572), .Z(N573) );
  GTECH_AND2 C896 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[13]), .Z(
        N571) );
  GTECH_AND2 C897 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[12]), .Z(
        N572) );
  GTECH_AND2 C898 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[13]), .Z(
        N574) );
  GTECH_AND2 C899 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[12]), .Z(
        N576) );
  GTECH_AND2 C900 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N578) );
  GTECH_NOT I_41 ( .A(N588), .Z(div_norm_inv_in[12]) );
  GTECH_OR2 C902 ( .A(N586), .B(N587), .Z(N588) );
  GTECH_OR2 C903 ( .A(N584), .B(N585), .Z(N586) );
  GTECH_OR2 C904 ( .A(N582), .B(N583), .Z(N584) );
  GTECH_OR2 C905 ( .A(N580), .B(N581), .Z(N582) );
  GTECH_AND2 C906 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[12]), .Z(
        N580) );
  GTECH_AND2 C907 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[11]), .Z(
        N581) );
  GTECH_AND2 C908 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[12]), .Z(
        N583) );
  GTECH_AND2 C909 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[11]), .Z(
        N585) );
  GTECH_AND2 C910 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N587) );
  GTECH_NOT I_42 ( .A(N597), .Z(div_norm_inv_in[11]) );
  GTECH_OR2 C912 ( .A(N595), .B(N596), .Z(N597) );
  GTECH_OR2 C913 ( .A(N593), .B(N594), .Z(N595) );
  GTECH_OR2 C914 ( .A(N591), .B(N592), .Z(N593) );
  GTECH_OR2 C915 ( .A(N589), .B(N590), .Z(N591) );
  GTECH_AND2 C916 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[11]), .Z(
        N589) );
  GTECH_AND2 C917 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[10]), .Z(
        N590) );
  GTECH_AND2 C918 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[11]), .Z(
        N592) );
  GTECH_AND2 C919 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[10]), .Z(
        N594) );
  GTECH_AND2 C920 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N596) );
  GTECH_NOT I_43 ( .A(N606), .Z(div_norm_inv_in[10]) );
  GTECH_OR2 C922 ( .A(N604), .B(N605), .Z(N606) );
  GTECH_OR2 C923 ( .A(N602), .B(N603), .Z(N604) );
  GTECH_OR2 C924 ( .A(N600), .B(N601), .Z(N602) );
  GTECH_OR2 C925 ( .A(N598), .B(N599), .Z(N600) );
  GTECH_AND2 C926 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[10]), .Z(
        N598) );
  GTECH_AND2 C927 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[9]), .Z(
        N599) );
  GTECH_AND2 C928 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[10]), .Z(
        N601) );
  GTECH_AND2 C929 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[9]), .Z(
        N603) );
  GTECH_AND2 C930 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N605) );
  GTECH_NOT I_44 ( .A(N615), .Z(div_norm_inv_in[9]) );
  GTECH_OR2 C932 ( .A(N613), .B(N614), .Z(N615) );
  GTECH_OR2 C933 ( .A(N611), .B(N612), .Z(N613) );
  GTECH_OR2 C934 ( .A(N609), .B(N610), .Z(N611) );
  GTECH_OR2 C935 ( .A(N607), .B(N608), .Z(N609) );
  GTECH_AND2 C936 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[9]), .Z(
        N607) );
  GTECH_AND2 C937 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[8]), .Z(
        N608) );
  GTECH_AND2 C938 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[9]), .Z(
        N610) );
  GTECH_AND2 C939 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[8]), .Z(
        N612) );
  GTECH_AND2 C940 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N614) );
  GTECH_NOT I_45 ( .A(N624), .Z(div_norm_inv_in[8]) );
  GTECH_OR2 C942 ( .A(N622), .B(N623), .Z(N624) );
  GTECH_OR2 C943 ( .A(N620), .B(N621), .Z(N622) );
  GTECH_OR2 C944 ( .A(N618), .B(N619), .Z(N620) );
  GTECH_OR2 C945 ( .A(N616), .B(N617), .Z(N618) );
  GTECH_AND2 C946 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[8]), .Z(
        N616) );
  GTECH_AND2 C947 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[7]), .Z(
        N617) );
  GTECH_AND2 C948 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[8]), .Z(
        N619) );
  GTECH_AND2 C949 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[7]), .Z(
        N621) );
  GTECH_AND2 C950 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N623) );
  GTECH_NOT I_46 ( .A(N633), .Z(div_norm_inv_in[7]) );
  GTECH_OR2 C952 ( .A(N631), .B(N632), .Z(N633) );
  GTECH_OR2 C953 ( .A(N629), .B(N630), .Z(N631) );
  GTECH_OR2 C954 ( .A(N627), .B(N628), .Z(N629) );
  GTECH_OR2 C955 ( .A(N625), .B(N626), .Z(N627) );
  GTECH_AND2 C956 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[7]), .Z(
        N625) );
  GTECH_AND2 C957 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[6]), .Z(
        N626) );
  GTECH_AND2 C958 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[7]), .Z(
        N628) );
  GTECH_AND2 C959 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[6]), .Z(
        N630) );
  GTECH_AND2 C960 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N632) );
  GTECH_NOT I_47 ( .A(N642), .Z(div_norm_inv_in[6]) );
  GTECH_OR2 C962 ( .A(N640), .B(N641), .Z(N642) );
  GTECH_OR2 C963 ( .A(N638), .B(N639), .Z(N640) );
  GTECH_OR2 C964 ( .A(N636), .B(N637), .Z(N638) );
  GTECH_OR2 C965 ( .A(N634), .B(N635), .Z(N636) );
  GTECH_AND2 C966 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[6]), .Z(
        N634) );
  GTECH_AND2 C967 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[5]), .Z(
        N635) );
  GTECH_AND2 C968 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[6]), .Z(
        N637) );
  GTECH_AND2 C969 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[5]), .Z(
        N639) );
  GTECH_AND2 C970 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N641) );
  GTECH_NOT I_48 ( .A(N651), .Z(div_norm_inv_in[5]) );
  GTECH_OR2 C972 ( .A(N649), .B(N650), .Z(N651) );
  GTECH_OR2 C973 ( .A(N647), .B(N648), .Z(N649) );
  GTECH_OR2 C974 ( .A(N645), .B(N646), .Z(N647) );
  GTECH_OR2 C975 ( .A(N643), .B(N644), .Z(N645) );
  GTECH_AND2 C976 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[5]), .Z(
        N643) );
  GTECH_AND2 C977 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[4]), .Z(
        N644) );
  GTECH_AND2 C978 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[5]), .Z(
        N646) );
  GTECH_AND2 C979 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[4]), .Z(
        N648) );
  GTECH_AND2 C980 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N650) );
  GTECH_NOT I_49 ( .A(N660), .Z(div_norm_inv_in[4]) );
  GTECH_OR2 C982 ( .A(N658), .B(N659), .Z(N660) );
  GTECH_OR2 C983 ( .A(N656), .B(N657), .Z(N658) );
  GTECH_OR2 C984 ( .A(N654), .B(N655), .Z(N656) );
  GTECH_OR2 C985 ( .A(N652), .B(N653), .Z(N654) );
  GTECH_AND2 C986 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[4]), .Z(
        N652) );
  GTECH_AND2 C987 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[3]), .Z(
        N653) );
  GTECH_AND2 C988 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[4]), .Z(
        N655) );
  GTECH_AND2 C989 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[3]), .Z(
        N657) );
  GTECH_AND2 C990 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N659) );
  GTECH_NOT I_50 ( .A(N669), .Z(div_norm_inv_in[3]) );
  GTECH_OR2 C992 ( .A(N667), .B(N668), .Z(N669) );
  GTECH_OR2 C993 ( .A(N665), .B(N666), .Z(N667) );
  GTECH_OR2 C994 ( .A(N663), .B(N664), .Z(N665) );
  GTECH_OR2 C995 ( .A(N661), .B(N662), .Z(N663) );
  GTECH_AND2 C996 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[3]), .Z(
        N661) );
  GTECH_AND2 C997 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[2]), .Z(
        N662) );
  GTECH_AND2 C998 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[3]), .Z(
        N664) );
  GTECH_AND2 C999 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[2]), .Z(
        N666) );
  GTECH_AND2 C1000 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N668) );
  GTECH_NOT I_51 ( .A(N678), .Z(div_norm_inv_in[2]) );
  GTECH_OR2 C1002 ( .A(N676), .B(N677), .Z(N678) );
  GTECH_OR2 C1003 ( .A(N674), .B(N675), .Z(N676) );
  GTECH_OR2 C1004 ( .A(N672), .B(N673), .Z(N674) );
  GTECH_OR2 C1005 ( .A(N670), .B(N671), .Z(N672) );
  GTECH_AND2 C1006 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[2]), .Z(
        N670) );
  GTECH_AND2 C1007 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[1]), .Z(
        N671) );
  GTECH_AND2 C1008 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[2]), .Z(
        N673) );
  GTECH_AND2 C1009 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[1]), .Z(
        N675) );
  GTECH_AND2 C1010 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N677) );
  GTECH_NOT I_52 ( .A(N687), .Z(div_norm_inv_in[1]) );
  GTECH_OR2 C1012 ( .A(N685), .B(N686), .Z(N687) );
  GTECH_OR2 C1013 ( .A(N683), .B(N684), .Z(N685) );
  GTECH_OR2 C1014 ( .A(N681), .B(N682), .Z(N683) );
  GTECH_OR2 C1015 ( .A(N679), .B(N680), .Z(N681) );
  GTECH_AND2 C1016 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[1]), .Z(
        N679) );
  GTECH_AND2 C1017 ( .A(div_norm_frac_in1_dbl_dnrm), .B(div_frac_in1[0]), .Z(
        N680) );
  GTECH_AND2 C1018 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[1]), .Z(
        N682) );
  GTECH_AND2 C1019 ( .A(div_norm_frac_in2_dbl_dnrm), .B(div_frac_in2[0]), .Z(
        N684) );
  GTECH_AND2 C1020 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N686) );
  GTECH_NOT I_53 ( .A(N692), .Z(div_norm_inv_in[0]) );
  GTECH_OR2 C1022 ( .A(N690), .B(N691), .Z(N692) );
  GTECH_OR2 C1023 ( .A(N688), .B(N689), .Z(N690) );
  GTECH_AND2 C1024 ( .A(div_norm_frac_in1_dbl_norm), .B(div_frac_in1[0]), .Z(
        N688) );
  GTECH_AND2 C1025 ( .A(div_norm_frac_in2_dbl_norm), .B(div_frac_in2[0]), .Z(
        N689) );
  GTECH_AND2 C1026 ( .A(div_norm_qnan), .B(d1stg_dblop), .Z(N691) );
  GTECH_NOT I_54 ( .A(div_norm_inv[52]), .Z(div_norm[52]) );
  GTECH_NOT I_55 ( .A(div_norm_inv[51]), .Z(div_norm[51]) );
  GTECH_NOT I_56 ( .A(div_norm_inv[50]), .Z(div_norm[50]) );
  GTECH_NOT I_57 ( .A(div_norm_inv[49]), .Z(div_norm[49]) );
  GTECH_NOT I_58 ( .A(div_norm_inv[48]), .Z(div_norm[48]) );
  GTECH_NOT I_59 ( .A(div_norm_inv[47]), .Z(div_norm[47]) );
  GTECH_NOT I_60 ( .A(div_norm_inv[46]), .Z(div_norm[46]) );
  GTECH_NOT I_61 ( .A(div_norm_inv[45]), .Z(div_norm[45]) );
  GTECH_NOT I_62 ( .A(div_norm_inv[44]), .Z(div_norm[44]) );
  GTECH_NOT I_63 ( .A(div_norm_inv[43]), .Z(div_norm[43]) );
  GTECH_NOT I_64 ( .A(div_norm_inv[42]), .Z(div_norm[42]) );
  GTECH_NOT I_65 ( .A(div_norm_inv[41]), .Z(div_norm[41]) );
  GTECH_NOT I_66 ( .A(div_norm_inv[40]), .Z(div_norm[40]) );
  GTECH_NOT I_67 ( .A(div_norm_inv[39]), .Z(div_norm[39]) );
  GTECH_NOT I_68 ( .A(div_norm_inv[38]), .Z(div_norm[38]) );
  GTECH_NOT I_69 ( .A(div_norm_inv[37]), .Z(div_norm[37]) );
  GTECH_NOT I_70 ( .A(div_norm_inv[36]), .Z(div_norm[36]) );
  GTECH_NOT I_71 ( .A(div_norm_inv[35]), .Z(div_norm[35]) );
  GTECH_NOT I_72 ( .A(div_norm_inv[34]), .Z(div_norm[34]) );
  GTECH_NOT I_73 ( .A(div_norm_inv[33]), .Z(div_norm[33]) );
  GTECH_NOT I_74 ( .A(div_norm_inv[32]), .Z(div_norm[32]) );
  GTECH_NOT I_75 ( .A(div_norm_inv[31]), .Z(div_norm[31]) );
  GTECH_NOT I_76 ( .A(div_norm_inv[30]), .Z(div_norm[30]) );
  GTECH_NOT I_77 ( .A(div_norm_inv[29]), .Z(div_norm[29]) );
  GTECH_NOT I_78 ( .A(div_norm_inv[28]), .Z(div_norm[28]) );
  GTECH_NOT I_79 ( .A(div_norm_inv[27]), .Z(div_norm[27]) );
  GTECH_NOT I_80 ( .A(div_norm_inv[26]), .Z(div_norm[26]) );
  GTECH_NOT I_81 ( .A(div_norm_inv[25]), .Z(div_norm[25]) );
  GTECH_NOT I_82 ( .A(div_norm_inv[24]), .Z(div_norm[24]) );
  GTECH_NOT I_83 ( .A(div_norm_inv[23]), .Z(div_norm[23]) );
  GTECH_NOT I_84 ( .A(div_norm_inv[22]), .Z(div_norm[22]) );
  GTECH_NOT I_85 ( .A(div_norm_inv[21]), .Z(div_norm[21]) );
  GTECH_NOT I_86 ( .A(div_norm_inv[20]), .Z(div_norm[20]) );
  GTECH_NOT I_87 ( .A(div_norm_inv[19]), .Z(div_norm[19]) );
  GTECH_NOT I_88 ( .A(div_norm_inv[18]), .Z(div_norm[18]) );
  GTECH_NOT I_89 ( .A(div_norm_inv[17]), .Z(div_norm[17]) );
  GTECH_NOT I_90 ( .A(div_norm_inv[16]), .Z(div_norm[16]) );
  GTECH_NOT I_91 ( .A(div_norm_inv[15]), .Z(div_norm[15]) );
  GTECH_NOT I_92 ( .A(div_norm_inv[14]), .Z(div_norm[14]) );
  GTECH_NOT I_93 ( .A(div_norm_inv[13]), .Z(div_norm[13]) );
  GTECH_NOT I_94 ( .A(div_norm_inv[12]), .Z(div_norm[12]) );
  GTECH_NOT I_95 ( .A(div_norm_inv[11]), .Z(div_norm[11]) );
  GTECH_NOT I_96 ( .A(div_norm_inv[10]), .Z(div_norm[10]) );
  GTECH_NOT I_97 ( .A(div_norm_inv[9]), .Z(div_norm[9]) );
  GTECH_NOT I_98 ( .A(div_norm_inv[8]), .Z(div_norm[8]) );
  GTECH_NOT I_99 ( .A(div_norm_inv[7]), .Z(div_norm[7]) );
  GTECH_NOT I_100 ( .A(div_norm_inv[6]), .Z(div_norm[6]) );
  GTECH_NOT I_101 ( .A(div_norm_inv[5]), .Z(div_norm[5]) );
  GTECH_NOT I_102 ( .A(div_norm_inv[4]), .Z(div_norm[4]) );
  GTECH_NOT I_103 ( .A(div_norm_inv[3]), .Z(div_norm[3]) );
  GTECH_NOT I_104 ( .A(div_norm_inv[2]), .Z(div_norm[2]) );
  GTECH_NOT I_105 ( .A(div_norm_inv[1]), .Z(div_norm[1]) );
  GTECH_NOT I_106 ( .A(div_norm_inv[0]), .Z(div_norm[0]) );
  GTECH_AND2 C1080 ( .A(d4stg_fdiv), .B(N693), .Z(div_frac_add_in2_in[52]) );
  GTECH_NOT I_107 ( .A(div_shl_tmp[105]), .Z(N693) );
  GTECH_AND2 C1082 ( .A(d4stg_fdiv), .B(N694), .Z(div_frac_add_in2_in[51]) );
  GTECH_NOT I_108 ( .A(div_shl_tmp[104]), .Z(N694) );
  GTECH_AND2 C1084 ( .A(d4stg_fdiv), .B(N695), .Z(div_frac_add_in2_in[50]) );
  GTECH_NOT I_109 ( .A(div_shl_tmp[103]), .Z(N695) );
  GTECH_AND2 C1086 ( .A(d4stg_fdiv), .B(N696), .Z(div_frac_add_in2_in[49]) );
  GTECH_NOT I_110 ( .A(div_shl_tmp[102]), .Z(N696) );
  GTECH_AND2 C1088 ( .A(d4stg_fdiv), .B(N697), .Z(div_frac_add_in2_in[48]) );
  GTECH_NOT I_111 ( .A(div_shl_tmp[101]), .Z(N697) );
  GTECH_AND2 C1090 ( .A(d4stg_fdiv), .B(N698), .Z(div_frac_add_in2_in[47]) );
  GTECH_NOT I_112 ( .A(div_shl_tmp[100]), .Z(N698) );
  GTECH_AND2 C1092 ( .A(d4stg_fdiv), .B(N699), .Z(div_frac_add_in2_in[46]) );
  GTECH_NOT I_113 ( .A(div_shl_tmp[99]), .Z(N699) );
  GTECH_AND2 C1094 ( .A(d4stg_fdiv), .B(N700), .Z(div_frac_add_in2_in[45]) );
  GTECH_NOT I_114 ( .A(div_shl_tmp[98]), .Z(N700) );
  GTECH_AND2 C1096 ( .A(d4stg_fdiv), .B(N701), .Z(div_frac_add_in2_in[44]) );
  GTECH_NOT I_115 ( .A(div_shl_tmp[97]), .Z(N701) );
  GTECH_AND2 C1098 ( .A(d4stg_fdiv), .B(N702), .Z(div_frac_add_in2_in[43]) );
  GTECH_NOT I_116 ( .A(div_shl_tmp[96]), .Z(N702) );
  GTECH_AND2 C1100 ( .A(d4stg_fdiv), .B(N703), .Z(div_frac_add_in2_in[42]) );
  GTECH_NOT I_117 ( .A(div_shl_tmp[95]), .Z(N703) );
  GTECH_AND2 C1102 ( .A(d4stg_fdiv), .B(N704), .Z(div_frac_add_in2_in[41]) );
  GTECH_NOT I_118 ( .A(div_shl_tmp[94]), .Z(N704) );
  GTECH_AND2 C1104 ( .A(d4stg_fdiv), .B(N705), .Z(div_frac_add_in2_in[40]) );
  GTECH_NOT I_119 ( .A(div_shl_tmp[93]), .Z(N705) );
  GTECH_AND2 C1106 ( .A(d4stg_fdiv), .B(N706), .Z(div_frac_add_in2_in[39]) );
  GTECH_NOT I_120 ( .A(div_shl_tmp[92]), .Z(N706) );
  GTECH_AND2 C1108 ( .A(d4stg_fdiv), .B(N707), .Z(div_frac_add_in2_in[38]) );
  GTECH_NOT I_121 ( .A(div_shl_tmp[91]), .Z(N707) );
  GTECH_AND2 C1110 ( .A(d4stg_fdiv), .B(N708), .Z(div_frac_add_in2_in[37]) );
  GTECH_NOT I_122 ( .A(div_shl_tmp[90]), .Z(N708) );
  GTECH_AND2 C1112 ( .A(d4stg_fdiv), .B(N709), .Z(div_frac_add_in2_in[36]) );
  GTECH_NOT I_123 ( .A(div_shl_tmp[89]), .Z(N709) );
  GTECH_AND2 C1114 ( .A(d4stg_fdiv), .B(N710), .Z(div_frac_add_in2_in[35]) );
  GTECH_NOT I_124 ( .A(div_shl_tmp[88]), .Z(N710) );
  GTECH_AND2 C1116 ( .A(d4stg_fdiv), .B(N711), .Z(div_frac_add_in2_in[34]) );
  GTECH_NOT I_125 ( .A(div_shl_tmp[87]), .Z(N711) );
  GTECH_AND2 C1118 ( .A(d4stg_fdiv), .B(N712), .Z(div_frac_add_in2_in[33]) );
  GTECH_NOT I_126 ( .A(div_shl_tmp[86]), .Z(N712) );
  GTECH_AND2 C1120 ( .A(d4stg_fdiv), .B(N713), .Z(div_frac_add_in2_in[32]) );
  GTECH_NOT I_127 ( .A(div_shl_tmp[85]), .Z(N713) );
  GTECH_AND2 C1122 ( .A(d4stg_fdiv), .B(N714), .Z(div_frac_add_in2_in[31]) );
  GTECH_NOT I_128 ( .A(div_shl_tmp[84]), .Z(N714) );
  GTECH_AND2 C1124 ( .A(d4stg_fdiv), .B(N715), .Z(div_frac_add_in2_in[30]) );
  GTECH_NOT I_129 ( .A(div_shl_tmp[83]), .Z(N715) );
  GTECH_OR2 C1126 ( .A(N717), .B(N718), .Z(div_frac_add_in2_in[29]) );
  GTECH_AND2 C1127 ( .A(d4stg_fdiv), .B(N716), .Z(N717) );
  GTECH_NOT I_130 ( .A(div_shl_tmp[82]), .Z(N716) );
  GTECH_AND2 C1129 ( .A(d6stg_fdiv), .B(d6stg_fdivs), .Z(N718) );
  GTECH_AND2 C1130 ( .A(d4stg_fdiv), .B(N719), .Z(div_frac_add_in2_in[28]) );
  GTECH_NOT I_131 ( .A(div_shl_tmp[81]), .Z(N719) );
  GTECH_AND2 C1132 ( .A(d4stg_fdiv), .B(N720), .Z(div_frac_add_in2_in[27]) );
  GTECH_NOT I_132 ( .A(div_shl_tmp[80]), .Z(N720) );
  GTECH_AND2 C1134 ( .A(d4stg_fdiv), .B(N721), .Z(div_frac_add_in2_in[26]) );
  GTECH_NOT I_133 ( .A(div_shl_tmp[79]), .Z(N721) );
  GTECH_AND2 C1136 ( .A(d4stg_fdiv), .B(N722), .Z(div_frac_add_in2_in[25]) );
  GTECH_NOT I_134 ( .A(div_shl_tmp[78]), .Z(N722) );
  GTECH_AND2 C1138 ( .A(d4stg_fdiv), .B(N723), .Z(div_frac_add_in2_in[24]) );
  GTECH_NOT I_135 ( .A(div_shl_tmp[77]), .Z(N723) );
  GTECH_AND2 C1140 ( .A(d4stg_fdiv), .B(N724), .Z(div_frac_add_in2_in[23]) );
  GTECH_NOT I_136 ( .A(div_shl_tmp[76]), .Z(N724) );
  GTECH_AND2 C1142 ( .A(d4stg_fdiv), .B(N725), .Z(div_frac_add_in2_in[22]) );
  GTECH_NOT I_137 ( .A(div_shl_tmp[75]), .Z(N725) );
  GTECH_AND2 C1144 ( .A(d4stg_fdiv), .B(N726), .Z(div_frac_add_in2_in[21]) );
  GTECH_NOT I_138 ( .A(div_shl_tmp[74]), .Z(N726) );
  GTECH_AND2 C1146 ( .A(d4stg_fdiv), .B(N727), .Z(div_frac_add_in2_in[20]) );
  GTECH_NOT I_139 ( .A(div_shl_tmp[73]), .Z(N727) );
  GTECH_AND2 C1148 ( .A(d4stg_fdiv), .B(N728), .Z(div_frac_add_in2_in[19]) );
  GTECH_NOT I_140 ( .A(div_shl_tmp[72]), .Z(N728) );
  GTECH_AND2 C1150 ( .A(d4stg_fdiv), .B(N729), .Z(div_frac_add_in2_in[18]) );
  GTECH_NOT I_141 ( .A(div_shl_tmp[71]), .Z(N729) );
  GTECH_AND2 C1152 ( .A(d4stg_fdiv), .B(N730), .Z(div_frac_add_in2_in[17]) );
  GTECH_NOT I_142 ( .A(div_shl_tmp[70]), .Z(N730) );
  GTECH_AND2 C1154 ( .A(d4stg_fdiv), .B(N731), .Z(div_frac_add_in2_in[16]) );
  GTECH_NOT I_143 ( .A(div_shl_tmp[69]), .Z(N731) );
  GTECH_AND2 C1156 ( .A(d4stg_fdiv), .B(N732), .Z(div_frac_add_in2_in[15]) );
  GTECH_NOT I_144 ( .A(div_shl_tmp[68]), .Z(N732) );
  GTECH_AND2 C1158 ( .A(d4stg_fdiv), .B(N733), .Z(div_frac_add_in2_in[14]) );
  GTECH_NOT I_145 ( .A(div_shl_tmp[67]), .Z(N733) );
  GTECH_AND2 C1160 ( .A(d4stg_fdiv), .B(N734), .Z(div_frac_add_in2_in[13]) );
  GTECH_NOT I_146 ( .A(div_shl_tmp[66]), .Z(N734) );
  GTECH_AND2 C1162 ( .A(d4stg_fdiv), .B(N735), .Z(div_frac_add_in2_in[12]) );
  GTECH_NOT I_147 ( .A(div_shl_tmp[65]), .Z(N735) );
  GTECH_AND2 C1164 ( .A(d4stg_fdiv), .B(N736), .Z(div_frac_add_in2_in[11]) );
  GTECH_NOT I_148 ( .A(div_shl_tmp[64]), .Z(N736) );
  GTECH_AND2 C1166 ( .A(d4stg_fdiv), .B(N737), .Z(div_frac_add_in2_in[10]) );
  GTECH_NOT I_149 ( .A(div_shl_tmp[63]), .Z(N737) );
  GTECH_AND2 C1168 ( .A(d4stg_fdiv), .B(N738), .Z(div_frac_add_in2_in[9]) );
  GTECH_NOT I_150 ( .A(div_shl_tmp[62]), .Z(N738) );
  GTECH_AND2 C1170 ( .A(d4stg_fdiv), .B(N739), .Z(div_frac_add_in2_in[8]) );
  GTECH_NOT I_151 ( .A(div_shl_tmp[61]), .Z(N739) );
  GTECH_AND2 C1172 ( .A(d4stg_fdiv), .B(N740), .Z(div_frac_add_in2_in[7]) );
  GTECH_NOT I_152 ( .A(div_shl_tmp[60]), .Z(N740) );
  GTECH_AND2 C1174 ( .A(d4stg_fdiv), .B(N741), .Z(div_frac_add_in2_in[6]) );
  GTECH_NOT I_153 ( .A(div_shl_tmp[59]), .Z(N741) );
  GTECH_AND2 C1176 ( .A(d4stg_fdiv), .B(N742), .Z(div_frac_add_in2_in[5]) );
  GTECH_NOT I_154 ( .A(div_shl_tmp[58]), .Z(N742) );
  GTECH_AND2 C1178 ( .A(d4stg_fdiv), .B(N743), .Z(div_frac_add_in2_in[4]) );
  GTECH_NOT I_155 ( .A(div_shl_tmp[57]), .Z(N743) );
  GTECH_AND2 C1180 ( .A(d4stg_fdiv), .B(N744), .Z(div_frac_add_in2_in[3]) );
  GTECH_NOT I_156 ( .A(div_shl_tmp[56]), .Z(N744) );
  GTECH_AND2 C1182 ( .A(d4stg_fdiv), .B(N745), .Z(div_frac_add_in2_in[2]) );
  GTECH_NOT I_157 ( .A(div_shl_tmp[55]), .Z(N745) );
  GTECH_AND2 C1184 ( .A(d4stg_fdiv), .B(N746), .Z(div_frac_add_in2_in[1]) );
  GTECH_NOT I_158 ( .A(div_shl_tmp[54]), .Z(N746) );
  GTECH_OR2 C1186 ( .A(N748), .B(N749), .Z(div_frac_add_in2_in[0]) );
  GTECH_AND2 C1187 ( .A(d4stg_fdiv), .B(N747), .Z(N748) );
  GTECH_NOT I_159 ( .A(div_shl_tmp[53]), .Z(N747) );
  GTECH_AND2 C1189 ( .A(d6stg_fdiv), .B(d6stg_fdivd), .Z(N749) );
  GTECH_OR2 C1190 ( .A(N750), .B(N751), .Z(d6stg_frac_53) );
  GTECH_AND2 C1191 ( .A(d6stg_frac_out_shl1), .B(div_frac_out[52]), .Z(N750)
         );
  GTECH_AND2 C1192 ( .A(d6stg_frac_out_nosh), .B(div_frac_out_54_53[0]), .Z(
        N751) );
  GTECH_OR2 C1193 ( .A(N752), .B(N753), .Z(d6stg_frac_52) );
  GTECH_AND2 C1194 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[51]), .Z(N752)
         );
  GTECH_AND2 C1195 ( .A(d6stg_frac_out_nosh), .B(div_frac_out[52]), .Z(N753)
         );
  GTECH_OR2 C1196 ( .A(N754), .B(N755), .Z(d6stg_frac_51) );
  GTECH_AND2 C1197 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[50]), .Z(N754)
         );
  GTECH_AND2 C1198 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[51]), .Z(N755)
         );
  GTECH_OR2 C1199 ( .A(N756), .B(N757), .Z(d6stg_frac_50) );
  GTECH_AND2 C1200 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[49]), .Z(N756)
         );
  GTECH_AND2 C1201 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[50]), .Z(N757)
         );
  GTECH_OR2 C1202 ( .A(N758), .B(N759), .Z(d6stg_frac_49) );
  GTECH_AND2 C1203 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[48]), .Z(N758)
         );
  GTECH_AND2 C1204 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[49]), .Z(N759)
         );
  GTECH_OR2 C1205 ( .A(N760), .B(N761), .Z(d6stg_frac_48) );
  GTECH_AND2 C1206 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[47]), .Z(N760)
         );
  GTECH_AND2 C1207 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[48]), .Z(N761)
         );
  GTECH_OR2 C1208 ( .A(N762), .B(N763), .Z(d6stg_frac_47) );
  GTECH_AND2 C1209 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[46]), .Z(N762)
         );
  GTECH_AND2 C1210 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[47]), .Z(N763)
         );
  GTECH_OR2 C1211 ( .A(N764), .B(N765), .Z(d6stg_frac_46) );
  GTECH_AND2 C1212 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[45]), .Z(N764)
         );
  GTECH_AND2 C1213 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[46]), .Z(N765)
         );
  GTECH_OR2 C1214 ( .A(N766), .B(N767), .Z(d6stg_frac_45) );
  GTECH_AND2 C1215 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[44]), .Z(N766)
         );
  GTECH_AND2 C1216 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[45]), .Z(N767)
         );
  GTECH_OR2 C1217 ( .A(N768), .B(N769), .Z(d6stg_frac_44) );
  GTECH_AND2 C1218 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[43]), .Z(N768)
         );
  GTECH_AND2 C1219 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[44]), .Z(N769)
         );
  GTECH_OR2 C1220 ( .A(N770), .B(N771), .Z(d6stg_frac_43) );
  GTECH_AND2 C1221 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[42]), .Z(N770)
         );
  GTECH_AND2 C1222 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[43]), .Z(N771)
         );
  GTECH_OR2 C1223 ( .A(N772), .B(N773), .Z(d6stg_frac_42) );
  GTECH_AND2 C1224 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[41]), .Z(N772)
         );
  GTECH_AND2 C1225 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[42]), .Z(N773)
         );
  GTECH_OR2 C1226 ( .A(N774), .B(N775), .Z(d6stg_frac_41) );
  GTECH_AND2 C1227 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[40]), .Z(N774)
         );
  GTECH_AND2 C1228 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[41]), .Z(N775)
         );
  GTECH_OR2 C1229 ( .A(N776), .B(N777), .Z(d6stg_frac_40) );
  GTECH_AND2 C1230 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[39]), .Z(N776)
         );
  GTECH_AND2 C1231 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[40]), .Z(N777)
         );
  GTECH_OR2 C1232 ( .A(N778), .B(N779), .Z(d6stg_frac_39) );
  GTECH_AND2 C1233 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[38]), .Z(N778)
         );
  GTECH_AND2 C1234 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[39]), .Z(N779)
         );
  GTECH_OR2 C1235 ( .A(N780), .B(N781), .Z(d6stg_frac_38) );
  GTECH_AND2 C1236 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[37]), .Z(N780)
         );
  GTECH_AND2 C1237 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[38]), .Z(N781)
         );
  GTECH_OR2 C1238 ( .A(N782), .B(N783), .Z(d6stg_frac_37) );
  GTECH_AND2 C1239 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[36]), .Z(N782)
         );
  GTECH_AND2 C1240 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[37]), .Z(N783)
         );
  GTECH_OR2 C1241 ( .A(N784), .B(N785), .Z(d6stg_frac_36) );
  GTECH_AND2 C1242 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[35]), .Z(N784)
         );
  GTECH_AND2 C1243 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[36]), .Z(N785)
         );
  GTECH_OR2 C1244 ( .A(N786), .B(N787), .Z(d6stg_frac_35) );
  GTECH_AND2 C1245 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[34]), .Z(N786)
         );
  GTECH_AND2 C1246 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[35]), .Z(N787)
         );
  GTECH_OR2 C1247 ( .A(N788), .B(N789), .Z(d6stg_frac_34) );
  GTECH_AND2 C1248 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[33]), .Z(N788)
         );
  GTECH_AND2 C1249 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[34]), .Z(N789)
         );
  GTECH_OR2 C1250 ( .A(N790), .B(N791), .Z(d6stg_frac_33) );
  GTECH_AND2 C1251 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[32]), .Z(N790)
         );
  GTECH_AND2 C1252 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[33]), .Z(N791)
         );
  GTECH_OR2 C1253 ( .A(N792), .B(N793), .Z(d6stg_frac_32) );
  GTECH_AND2 C1254 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[31]), .Z(N792)
         );
  GTECH_AND2 C1255 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[32]), .Z(N793)
         );
  GTECH_OR2 C1256 ( .A(N794), .B(N795), .Z(d6stg_frac_31) );
  GTECH_AND2 C1257 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[30]), .Z(N794)
         );
  GTECH_AND2 C1258 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[31]), .Z(N795)
         );
  GTECH_OR2 C1259 ( .A(N796), .B(N797), .Z(d6stg_frac_30) );
  GTECH_AND2 C1260 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[29]), .Z(N796)
         );
  GTECH_AND2 C1261 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[30]), .Z(N797)
         );
  GTECH_OR2 C1262 ( .A(N798), .B(N799), .Z(d6stg_frac_29) );
  GTECH_AND2 C1263 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[28]), .Z(N798)
         );
  GTECH_AND2 C1264 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[29]), .Z(N799)
         );
  GTECH_OR2 C1265 ( .A(N800), .B(N801), .Z(d6stg_frac[28]) );
  GTECH_AND2 C1266 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[27]), .Z(N800)
         );
  GTECH_AND2 C1267 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[28]), .Z(N801)
         );
  GTECH_OR2 C1268 ( .A(N802), .B(N803), .Z(d6stg_frac[27]) );
  GTECH_AND2 C1269 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[26]), .Z(N802)
         );
  GTECH_AND2 C1270 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[27]), .Z(N803)
         );
  GTECH_OR2 C1271 ( .A(N804), .B(N805), .Z(d6stg_frac[26]) );
  GTECH_AND2 C1272 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[25]), .Z(N804)
         );
  GTECH_AND2 C1273 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[26]), .Z(N805)
         );
  GTECH_OR2 C1274 ( .A(N806), .B(N807), .Z(d6stg_frac[25]) );
  GTECH_AND2 C1275 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[24]), .Z(N806)
         );
  GTECH_AND2 C1276 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[25]), .Z(N807)
         );
  GTECH_OR2 C1277 ( .A(N808), .B(N809), .Z(d6stg_frac[24]) );
  GTECH_AND2 C1278 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[23]), .Z(N808)
         );
  GTECH_AND2 C1279 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[24]), .Z(N809)
         );
  GTECH_OR2 C1280 ( .A(N810), .B(N811), .Z(d6stg_frac[23]) );
  GTECH_AND2 C1281 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[22]), .Z(N810)
         );
  GTECH_AND2 C1282 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[23]), .Z(N811)
         );
  GTECH_OR2 C1283 ( .A(N812), .B(N813), .Z(d6stg_frac[22]) );
  GTECH_AND2 C1284 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[21]), .Z(N812)
         );
  GTECH_AND2 C1285 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[22]), .Z(N813)
         );
  GTECH_OR2 C1286 ( .A(N814), .B(N815), .Z(d6stg_frac[21]) );
  GTECH_AND2 C1287 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[20]), .Z(N814)
         );
  GTECH_AND2 C1288 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[21]), .Z(N815)
         );
  GTECH_OR2 C1289 ( .A(N816), .B(N817), .Z(d6stg_frac[20]) );
  GTECH_AND2 C1290 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[19]), .Z(N816)
         );
  GTECH_AND2 C1291 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[20]), .Z(N817)
         );
  GTECH_OR2 C1292 ( .A(N818), .B(N819), .Z(d6stg_frac[19]) );
  GTECH_AND2 C1293 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[18]), .Z(N818)
         );
  GTECH_AND2 C1294 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[19]), .Z(N819)
         );
  GTECH_OR2 C1295 ( .A(N820), .B(N821), .Z(d6stg_frac[18]) );
  GTECH_AND2 C1296 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[17]), .Z(N820)
         );
  GTECH_AND2 C1297 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[18]), .Z(N821)
         );
  GTECH_OR2 C1298 ( .A(N822), .B(N823), .Z(d6stg_frac[17]) );
  GTECH_AND2 C1299 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[16]), .Z(N822)
         );
  GTECH_AND2 C1300 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[17]), .Z(N823)
         );
  GTECH_OR2 C1301 ( .A(N824), .B(N825), .Z(d6stg_frac[16]) );
  GTECH_AND2 C1302 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[15]), .Z(N824)
         );
  GTECH_AND2 C1303 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[16]), .Z(N825)
         );
  GTECH_OR2 C1304 ( .A(N826), .B(N827), .Z(d6stg_frac[15]) );
  GTECH_AND2 C1305 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[14]), .Z(N826)
         );
  GTECH_AND2 C1306 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[15]), .Z(N827)
         );
  GTECH_OR2 C1307 ( .A(N828), .B(N829), .Z(d6stg_frac[14]) );
  GTECH_AND2 C1308 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[13]), .Z(N828)
         );
  GTECH_AND2 C1309 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[14]), .Z(N829)
         );
  GTECH_OR2 C1310 ( .A(N830), .B(N831), .Z(d6stg_frac[13]) );
  GTECH_AND2 C1311 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[12]), .Z(N830)
         );
  GTECH_AND2 C1312 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[13]), .Z(N831)
         );
  GTECH_OR2 C1313 ( .A(N832), .B(N833), .Z(d6stg_frac[12]) );
  GTECH_AND2 C1314 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[11]), .Z(N832)
         );
  GTECH_AND2 C1315 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[12]), .Z(N833)
         );
  GTECH_OR2 C1316 ( .A(N834), .B(N835), .Z(d6stg_frac[11]) );
  GTECH_AND2 C1317 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[10]), .Z(N834)
         );
  GTECH_AND2 C1318 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[11]), .Z(N835)
         );
  GTECH_OR2 C1319 ( .A(N836), .B(N837), .Z(d6stg_frac[10]) );
  GTECH_AND2 C1320 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[9]), .Z(N836)
         );
  GTECH_AND2 C1321 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[10]), .Z(N837)
         );
  GTECH_OR2 C1322 ( .A(N838), .B(N839), .Z(d6stg_frac[9]) );
  GTECH_AND2 C1323 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[8]), .Z(N838)
         );
  GTECH_AND2 C1324 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[9]), .Z(N839)
         );
  GTECH_OR2 C1325 ( .A(N840), .B(N841), .Z(d6stg_frac[8]) );
  GTECH_AND2 C1326 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[7]), .Z(N840)
         );
  GTECH_AND2 C1327 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[8]), .Z(N841)
         );
  GTECH_OR2 C1328 ( .A(N842), .B(N843), .Z(d6stg_frac[7]) );
  GTECH_AND2 C1329 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[6]), .Z(N842)
         );
  GTECH_AND2 C1330 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[7]), .Z(N843)
         );
  GTECH_OR2 C1331 ( .A(N844), .B(N845), .Z(d6stg_frac[6]) );
  GTECH_AND2 C1332 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[5]), .Z(N844)
         );
  GTECH_AND2 C1333 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[6]), .Z(N845)
         );
  GTECH_OR2 C1334 ( .A(N846), .B(N847), .Z(d6stg_frac[5]) );
  GTECH_AND2 C1335 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[4]), .Z(N846)
         );
  GTECH_AND2 C1336 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[5]), .Z(N847)
         );
  GTECH_OR2 C1337 ( .A(N848), .B(N849), .Z(d6stg_frac[4]) );
  GTECH_AND2 C1338 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[3]), .Z(N848)
         );
  GTECH_AND2 C1339 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[4]), .Z(N849)
         );
  GTECH_OR2 C1340 ( .A(N850), .B(N851), .Z(d6stg_frac[3]) );
  GTECH_AND2 C1341 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[2]), .Z(N850)
         );
  GTECH_AND2 C1342 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[3]), .Z(N851)
         );
  GTECH_OR2 C1343 ( .A(N852), .B(N853), .Z(d6stg_frac_2) );
  GTECH_AND2 C1344 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[1]), .Z(N852)
         );
  GTECH_AND2 C1345 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[2]), .Z(N853)
         );
  GTECH_OR2 C1346 ( .A(N854), .B(N855), .Z(d6stg_frac_1) );
  GTECH_AND2 C1347 ( .A(d6stg_frac_out_shl1), .B(div_frac_outa[0]), .Z(N854)
         );
  GTECH_AND2 C1348 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[1]), .Z(N855)
         );
  GTECH_AND2 C1349 ( .A(d6stg_frac_out_nosh), .B(div_frac_outa[0]), .Z(
        d6stg_frac_0) );
  GTECH_OR2 C1350 ( .A(N860), .B(N862), .Z(div_frac_add_in1_in[54]) );
  GTECH_OR2 C1351 ( .A(N856), .B(N859), .Z(N860) );
  GTECH_AND2 C1352 ( .A(d4stg_fdiv), .B(div_shl_save[54]), .Z(N856) );
  GTECH_AND2 C1353 ( .A(N858), .B(div_frac_add[53]), .Z(N859) );
  GTECH_AND2 C1354 ( .A(div_frac_add_in1_add), .B(N857), .Z(N858) );
  GTECH_NOT I_160 ( .A(div_frac_add[54]), .Z(N857) );
  GTECH_AND2 C1356 ( .A(N861), .B(div_frac_add_in1[53]), .Z(N862) );
  GTECH_AND2 C1357 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N861)
         );
  GTECH_OR2 C1358 ( .A(N866), .B(N868), .Z(div_frac_add_in1_in[53]) );
  GTECH_OR2 C1359 ( .A(N863), .B(N865), .Z(N866) );
  GTECH_AND2 C1360 ( .A(d4stg_fdiv), .B(div_shl_save[53]), .Z(N863) );
  GTECH_AND2 C1361 ( .A(N864), .B(div_frac_add[52]), .Z(N865) );
  GTECH_AND2 C1362 ( .A(div_frac_add_in1_add), .B(N857), .Z(N864) );
  GTECH_AND2 C1364 ( .A(N867), .B(div_frac_add_in1[52]), .Z(N868) );
  GTECH_AND2 C1365 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N867)
         );
  GTECH_OR2 C1366 ( .A(N872), .B(N874), .Z(div_frac_add_in1_in[52]) );
  GTECH_OR2 C1367 ( .A(N869), .B(N871), .Z(N872) );
  GTECH_AND2 C1368 ( .A(d4stg_fdiv), .B(div_shl_save[52]), .Z(N869) );
  GTECH_AND2 C1369 ( .A(N870), .B(div_frac_add[51]), .Z(N871) );
  GTECH_AND2 C1370 ( .A(div_frac_add_in1_add), .B(N857), .Z(N870) );
  GTECH_AND2 C1372 ( .A(N873), .B(div_frac_add_in1[51]), .Z(N874) );
  GTECH_AND2 C1373 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N873)
         );
  GTECH_OR2 C1374 ( .A(N881), .B(N882), .Z(div_frac_add_in1_in[51]) );
  GTECH_OR2 C1375 ( .A(N878), .B(N880), .Z(N881) );
  GTECH_OR2 C1376 ( .A(N875), .B(N877), .Z(N878) );
  GTECH_AND2 C1377 ( .A(d4stg_fdiv), .B(div_shl_save[51]), .Z(N875) );
  GTECH_AND2 C1378 ( .A(N876), .B(div_frac_add[50]), .Z(N877) );
  GTECH_AND2 C1379 ( .A(div_frac_add_in1_add), .B(N857), .Z(N876) );
  GTECH_AND2 C1381 ( .A(N879), .B(div_frac_add_in1[50]), .Z(N880) );
  GTECH_AND2 C1382 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N879)
         );
  GTECH_AND2 C1383 ( .A(d6stg_fdiv), .B(d6stg_frac_53), .Z(N882) );
  GTECH_OR2 C1384 ( .A(N889), .B(N890), .Z(div_frac_add_in1_in[50]) );
  GTECH_OR2 C1385 ( .A(N886), .B(N888), .Z(N889) );
  GTECH_OR2 C1386 ( .A(N883), .B(N885), .Z(N886) );
  GTECH_AND2 C1387 ( .A(d4stg_fdiv), .B(div_shl_save[50]), .Z(N883) );
  GTECH_AND2 C1388 ( .A(N884), .B(div_frac_add[49]), .Z(N885) );
  GTECH_AND2 C1389 ( .A(div_frac_add_in1_add), .B(N857), .Z(N884) );
  GTECH_AND2 C1391 ( .A(N887), .B(div_frac_add_in1[49]), .Z(N888) );
  GTECH_AND2 C1392 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N887)
         );
  GTECH_AND2 C1393 ( .A(d6stg_fdiv), .B(d6stg_frac_52), .Z(N890) );
  GTECH_OR2 C1394 ( .A(N897), .B(N898), .Z(div_frac_add_in1_in[49]) );
  GTECH_OR2 C1395 ( .A(N894), .B(N896), .Z(N897) );
  GTECH_OR2 C1396 ( .A(N891), .B(N893), .Z(N894) );
  GTECH_AND2 C1397 ( .A(d4stg_fdiv), .B(div_shl_save[49]), .Z(N891) );
  GTECH_AND2 C1398 ( .A(N892), .B(div_frac_add[48]), .Z(N893) );
  GTECH_AND2 C1399 ( .A(div_frac_add_in1_add), .B(N857), .Z(N892) );
  GTECH_AND2 C1401 ( .A(N895), .B(div_frac_add_in1[48]), .Z(N896) );
  GTECH_AND2 C1402 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N895)
         );
  GTECH_AND2 C1403 ( .A(d6stg_fdiv), .B(d6stg_frac_51), .Z(N898) );
  GTECH_OR2 C1404 ( .A(N905), .B(N906), .Z(div_frac_add_in1_in[48]) );
  GTECH_OR2 C1405 ( .A(N902), .B(N904), .Z(N905) );
  GTECH_OR2 C1406 ( .A(N899), .B(N901), .Z(N902) );
  GTECH_AND2 C1407 ( .A(d4stg_fdiv), .B(div_shl_save[48]), .Z(N899) );
  GTECH_AND2 C1408 ( .A(N900), .B(div_frac_add[47]), .Z(N901) );
  GTECH_AND2 C1409 ( .A(div_frac_add_in1_add), .B(N857), .Z(N900) );
  GTECH_AND2 C1411 ( .A(N903), .B(div_frac_add_in1[47]), .Z(N904) );
  GTECH_AND2 C1412 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N903)
         );
  GTECH_AND2 C1413 ( .A(d6stg_fdiv), .B(d6stg_frac_50), .Z(N906) );
  GTECH_OR2 C1414 ( .A(N913), .B(N914), .Z(div_frac_add_in1_in[47]) );
  GTECH_OR2 C1415 ( .A(N910), .B(N912), .Z(N913) );
  GTECH_OR2 C1416 ( .A(N907), .B(N909), .Z(N910) );
  GTECH_AND2 C1417 ( .A(d4stg_fdiv), .B(div_shl_save[47]), .Z(N907) );
  GTECH_AND2 C1418 ( .A(N908), .B(div_frac_add[46]), .Z(N909) );
  GTECH_AND2 C1419 ( .A(div_frac_add_in1_add), .B(N857), .Z(N908) );
  GTECH_AND2 C1421 ( .A(N911), .B(div_frac_add_in1[46]), .Z(N912) );
  GTECH_AND2 C1422 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N911)
         );
  GTECH_AND2 C1423 ( .A(d6stg_fdiv), .B(d6stg_frac_49), .Z(N914) );
  GTECH_OR2 C1424 ( .A(N921), .B(N922), .Z(div_frac_add_in1_in[46]) );
  GTECH_OR2 C1425 ( .A(N918), .B(N920), .Z(N921) );
  GTECH_OR2 C1426 ( .A(N915), .B(N917), .Z(N918) );
  GTECH_AND2 C1427 ( .A(d4stg_fdiv), .B(div_shl_save[46]), .Z(N915) );
  GTECH_AND2 C1428 ( .A(N916), .B(div_frac_add[45]), .Z(N917) );
  GTECH_AND2 C1429 ( .A(div_frac_add_in1_add), .B(N857), .Z(N916) );
  GTECH_AND2 C1431 ( .A(N919), .B(div_frac_add_in1[45]), .Z(N920) );
  GTECH_AND2 C1432 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N919)
         );
  GTECH_AND2 C1433 ( .A(d6stg_fdiv), .B(d6stg_frac_48), .Z(N922) );
  GTECH_OR2 C1434 ( .A(N929), .B(N930), .Z(div_frac_add_in1_in[45]) );
  GTECH_OR2 C1435 ( .A(N926), .B(N928), .Z(N929) );
  GTECH_OR2 C1436 ( .A(N923), .B(N925), .Z(N926) );
  GTECH_AND2 C1437 ( .A(d4stg_fdiv), .B(div_shl_save[45]), .Z(N923) );
  GTECH_AND2 C1438 ( .A(N924), .B(div_frac_add[44]), .Z(N925) );
  GTECH_AND2 C1439 ( .A(div_frac_add_in1_add), .B(N857), .Z(N924) );
  GTECH_AND2 C1441 ( .A(N927), .B(div_frac_add_in1[44]), .Z(N928) );
  GTECH_AND2 C1442 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N927)
         );
  GTECH_AND2 C1443 ( .A(d6stg_fdiv), .B(d6stg_frac_47), .Z(N930) );
  GTECH_OR2 C1444 ( .A(N937), .B(N938), .Z(div_frac_add_in1_in[44]) );
  GTECH_OR2 C1445 ( .A(N934), .B(N936), .Z(N937) );
  GTECH_OR2 C1446 ( .A(N931), .B(N933), .Z(N934) );
  GTECH_AND2 C1447 ( .A(d4stg_fdiv), .B(div_shl_save[44]), .Z(N931) );
  GTECH_AND2 C1448 ( .A(N932), .B(div_frac_add[43]), .Z(N933) );
  GTECH_AND2 C1449 ( .A(div_frac_add_in1_add), .B(N857), .Z(N932) );
  GTECH_AND2 C1451 ( .A(N935), .B(div_frac_add_in1[43]), .Z(N936) );
  GTECH_AND2 C1452 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N935)
         );
  GTECH_AND2 C1453 ( .A(d6stg_fdiv), .B(d6stg_frac_46), .Z(N938) );
  GTECH_OR2 C1454 ( .A(N945), .B(N946), .Z(div_frac_add_in1_in[43]) );
  GTECH_OR2 C1455 ( .A(N942), .B(N944), .Z(N945) );
  GTECH_OR2 C1456 ( .A(N939), .B(N941), .Z(N942) );
  GTECH_AND2 C1457 ( .A(d4stg_fdiv), .B(div_shl_save[43]), .Z(N939) );
  GTECH_AND2 C1458 ( .A(N940), .B(div_frac_add[42]), .Z(N941) );
  GTECH_AND2 C1459 ( .A(div_frac_add_in1_add), .B(N857), .Z(N940) );
  GTECH_AND2 C1461 ( .A(N943), .B(div_frac_add_in1[42]), .Z(N944) );
  GTECH_AND2 C1462 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N943)
         );
  GTECH_AND2 C1463 ( .A(d6stg_fdiv), .B(d6stg_frac_45), .Z(N946) );
  GTECH_OR2 C1464 ( .A(N953), .B(N954), .Z(div_frac_add_in1_in[42]) );
  GTECH_OR2 C1465 ( .A(N950), .B(N952), .Z(N953) );
  GTECH_OR2 C1466 ( .A(N947), .B(N949), .Z(N950) );
  GTECH_AND2 C1467 ( .A(d4stg_fdiv), .B(div_shl_save[42]), .Z(N947) );
  GTECH_AND2 C1468 ( .A(N948), .B(div_frac_add[41]), .Z(N949) );
  GTECH_AND2 C1469 ( .A(div_frac_add_in1_add), .B(N857), .Z(N948) );
  GTECH_AND2 C1471 ( .A(N951), .B(div_frac_add_in1[41]), .Z(N952) );
  GTECH_AND2 C1472 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N951)
         );
  GTECH_AND2 C1473 ( .A(d6stg_fdiv), .B(d6stg_frac_44), .Z(N954) );
  GTECH_OR2 C1474 ( .A(N961), .B(N962), .Z(div_frac_add_in1_in[41]) );
  GTECH_OR2 C1475 ( .A(N958), .B(N960), .Z(N961) );
  GTECH_OR2 C1476 ( .A(N955), .B(N957), .Z(N958) );
  GTECH_AND2 C1477 ( .A(d4stg_fdiv), .B(div_shl_save[41]), .Z(N955) );
  GTECH_AND2 C1478 ( .A(N956), .B(div_frac_add[40]), .Z(N957) );
  GTECH_AND2 C1479 ( .A(div_frac_add_in1_add), .B(N857), .Z(N956) );
  GTECH_AND2 C1481 ( .A(N959), .B(div_frac_add_in1[40]), .Z(N960) );
  GTECH_AND2 C1482 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N959)
         );
  GTECH_AND2 C1483 ( .A(d6stg_fdiv), .B(d6stg_frac_43), .Z(N962) );
  GTECH_OR2 C1484 ( .A(N969), .B(N970), .Z(div_frac_add_in1_in[40]) );
  GTECH_OR2 C1485 ( .A(N966), .B(N968), .Z(N969) );
  GTECH_OR2 C1486 ( .A(N963), .B(N965), .Z(N966) );
  GTECH_AND2 C1487 ( .A(d4stg_fdiv), .B(div_shl_save[40]), .Z(N963) );
  GTECH_AND2 C1488 ( .A(N964), .B(div_frac_add[39]), .Z(N965) );
  GTECH_AND2 C1489 ( .A(div_frac_add_in1_add), .B(N857), .Z(N964) );
  GTECH_AND2 C1491 ( .A(N967), .B(div_frac_add_in1[39]), .Z(N968) );
  GTECH_AND2 C1492 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N967)
         );
  GTECH_AND2 C1493 ( .A(d6stg_fdiv), .B(d6stg_frac_42), .Z(N970) );
  GTECH_OR2 C1494 ( .A(N977), .B(N978), .Z(div_frac_add_in1_in[39]) );
  GTECH_OR2 C1495 ( .A(N974), .B(N976), .Z(N977) );
  GTECH_OR2 C1496 ( .A(N971), .B(N973), .Z(N974) );
  GTECH_AND2 C1497 ( .A(d4stg_fdiv), .B(div_shl_save[39]), .Z(N971) );
  GTECH_AND2 C1498 ( .A(N972), .B(div_frac_add[38]), .Z(N973) );
  GTECH_AND2 C1499 ( .A(div_frac_add_in1_add), .B(N857), .Z(N972) );
  GTECH_AND2 C1501 ( .A(N975), .B(div_frac_add_in1[38]), .Z(N976) );
  GTECH_AND2 C1502 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N975)
         );
  GTECH_AND2 C1503 ( .A(d6stg_fdiv), .B(d6stg_frac_41), .Z(N978) );
  GTECH_OR2 C1504 ( .A(N985), .B(N986), .Z(div_frac_add_in1_in[38]) );
  GTECH_OR2 C1505 ( .A(N982), .B(N984), .Z(N985) );
  GTECH_OR2 C1506 ( .A(N979), .B(N981), .Z(N982) );
  GTECH_AND2 C1507 ( .A(d4stg_fdiv), .B(div_shl_save[38]), .Z(N979) );
  GTECH_AND2 C1508 ( .A(N980), .B(div_frac_add[37]), .Z(N981) );
  GTECH_AND2 C1509 ( .A(div_frac_add_in1_add), .B(N857), .Z(N980) );
  GTECH_AND2 C1511 ( .A(N983), .B(div_frac_add_in1[37]), .Z(N984) );
  GTECH_AND2 C1512 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N983)
         );
  GTECH_AND2 C1513 ( .A(d6stg_fdiv), .B(d6stg_frac_40), .Z(N986) );
  GTECH_OR2 C1514 ( .A(N993), .B(N994), .Z(div_frac_add_in1_in[37]) );
  GTECH_OR2 C1515 ( .A(N990), .B(N992), .Z(N993) );
  GTECH_OR2 C1516 ( .A(N987), .B(N989), .Z(N990) );
  GTECH_AND2 C1517 ( .A(d4stg_fdiv), .B(div_shl_save[37]), .Z(N987) );
  GTECH_AND2 C1518 ( .A(N988), .B(div_frac_add[36]), .Z(N989) );
  GTECH_AND2 C1519 ( .A(div_frac_add_in1_add), .B(N857), .Z(N988) );
  GTECH_AND2 C1521 ( .A(N991), .B(div_frac_add_in1[36]), .Z(N992) );
  GTECH_AND2 C1522 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N991)
         );
  GTECH_AND2 C1523 ( .A(d6stg_fdiv), .B(d6stg_frac_39), .Z(N994) );
  GTECH_OR2 C1524 ( .A(N1001), .B(N1002), .Z(div_frac_add_in1_in[36]) );
  GTECH_OR2 C1525 ( .A(N998), .B(N1000), .Z(N1001) );
  GTECH_OR2 C1526 ( .A(N995), .B(N997), .Z(N998) );
  GTECH_AND2 C1527 ( .A(d4stg_fdiv), .B(div_shl_save[36]), .Z(N995) );
  GTECH_AND2 C1528 ( .A(N996), .B(div_frac_add[35]), .Z(N997) );
  GTECH_AND2 C1529 ( .A(div_frac_add_in1_add), .B(N857), .Z(N996) );
  GTECH_AND2 C1531 ( .A(N999), .B(div_frac_add_in1[35]), .Z(N1000) );
  GTECH_AND2 C1532 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N999)
         );
  GTECH_AND2 C1533 ( .A(d6stg_fdiv), .B(d6stg_frac_38), .Z(N1002) );
  GTECH_OR2 C1534 ( .A(N1009), .B(N1010), .Z(div_frac_add_in1_in[35]) );
  GTECH_OR2 C1535 ( .A(N1006), .B(N1008), .Z(N1009) );
  GTECH_OR2 C1536 ( .A(N1003), .B(N1005), .Z(N1006) );
  GTECH_AND2 C1537 ( .A(d4stg_fdiv), .B(div_shl_save[35]), .Z(N1003) );
  GTECH_AND2 C1538 ( .A(N1004), .B(div_frac_add[34]), .Z(N1005) );
  GTECH_AND2 C1539 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1004) );
  GTECH_AND2 C1541 ( .A(N1007), .B(div_frac_add_in1[34]), .Z(N1008) );
  GTECH_AND2 C1542 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1007)
         );
  GTECH_AND2 C1543 ( .A(d6stg_fdiv), .B(d6stg_frac_37), .Z(N1010) );
  GTECH_OR2 C1544 ( .A(N1017), .B(N1018), .Z(div_frac_add_in1_in[34]) );
  GTECH_OR2 C1545 ( .A(N1014), .B(N1016), .Z(N1017) );
  GTECH_OR2 C1546 ( .A(N1011), .B(N1013), .Z(N1014) );
  GTECH_AND2 C1547 ( .A(d4stg_fdiv), .B(div_shl_save[34]), .Z(N1011) );
  GTECH_AND2 C1548 ( .A(N1012), .B(div_frac_add[33]), .Z(N1013) );
  GTECH_AND2 C1549 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1012) );
  GTECH_AND2 C1551 ( .A(N1015), .B(div_frac_add_in1[33]), .Z(N1016) );
  GTECH_AND2 C1552 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1015)
         );
  GTECH_AND2 C1553 ( .A(d6stg_fdiv), .B(d6stg_frac_36), .Z(N1018) );
  GTECH_OR2 C1554 ( .A(N1025), .B(N1026), .Z(div_frac_add_in1_in[33]) );
  GTECH_OR2 C1555 ( .A(N1022), .B(N1024), .Z(N1025) );
  GTECH_OR2 C1556 ( .A(N1019), .B(N1021), .Z(N1022) );
  GTECH_AND2 C1557 ( .A(d4stg_fdiv), .B(div_shl_save[33]), .Z(N1019) );
  GTECH_AND2 C1558 ( .A(N1020), .B(div_frac_add[32]), .Z(N1021) );
  GTECH_AND2 C1559 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1020) );
  GTECH_AND2 C1561 ( .A(N1023), .B(div_frac_add_in1[32]), .Z(N1024) );
  GTECH_AND2 C1562 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1023)
         );
  GTECH_AND2 C1563 ( .A(d6stg_fdiv), .B(d6stg_frac_35), .Z(N1026) );
  GTECH_OR2 C1564 ( .A(N1033), .B(N1034), .Z(div_frac_add_in1_in[32]) );
  GTECH_OR2 C1565 ( .A(N1030), .B(N1032), .Z(N1033) );
  GTECH_OR2 C1566 ( .A(N1027), .B(N1029), .Z(N1030) );
  GTECH_AND2 C1567 ( .A(d4stg_fdiv), .B(div_shl_save[32]), .Z(N1027) );
  GTECH_AND2 C1568 ( .A(N1028), .B(div_frac_add[31]), .Z(N1029) );
  GTECH_AND2 C1569 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1028) );
  GTECH_AND2 C1571 ( .A(N1031), .B(div_frac_add_in1[31]), .Z(N1032) );
  GTECH_AND2 C1572 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1031)
         );
  GTECH_AND2 C1573 ( .A(d6stg_fdiv), .B(d6stg_frac_34), .Z(N1034) );
  GTECH_OR2 C1574 ( .A(N1041), .B(N1042), .Z(div_frac_add_in1_in[31]) );
  GTECH_OR2 C1575 ( .A(N1038), .B(N1040), .Z(N1041) );
  GTECH_OR2 C1576 ( .A(N1035), .B(N1037), .Z(N1038) );
  GTECH_AND2 C1577 ( .A(d4stg_fdiv), .B(div_shl_save[31]), .Z(N1035) );
  GTECH_AND2 C1578 ( .A(N1036), .B(div_frac_add[30]), .Z(N1037) );
  GTECH_AND2 C1579 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1036) );
  GTECH_AND2 C1581 ( .A(N1039), .B(div_frac_add_in1[30]), .Z(N1040) );
  GTECH_AND2 C1582 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1039)
         );
  GTECH_AND2 C1583 ( .A(d6stg_fdiv), .B(d6stg_frac_33), .Z(N1042) );
  GTECH_OR2 C1584 ( .A(N1049), .B(N1050), .Z(div_frac_add_in1_in[30]) );
  GTECH_OR2 C1585 ( .A(N1046), .B(N1048), .Z(N1049) );
  GTECH_OR2 C1586 ( .A(N1043), .B(N1045), .Z(N1046) );
  GTECH_AND2 C1587 ( .A(d4stg_fdiv), .B(div_shl_save[30]), .Z(N1043) );
  GTECH_AND2 C1588 ( .A(N1044), .B(div_frac_add[29]), .Z(N1045) );
  GTECH_AND2 C1589 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1044) );
  GTECH_AND2 C1591 ( .A(N1047), .B(div_frac_add_in1[29]), .Z(N1048) );
  GTECH_AND2 C1592 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1047)
         );
  GTECH_AND2 C1593 ( .A(d6stg_fdiv), .B(d6stg_frac_32), .Z(N1050) );
  GTECH_OR2 C1594 ( .A(N1057), .B(N1058), .Z(div_frac_add_in1_in[29]) );
  GTECH_OR2 C1595 ( .A(N1054), .B(N1056), .Z(N1057) );
  GTECH_OR2 C1596 ( .A(N1051), .B(N1053), .Z(N1054) );
  GTECH_AND2 C1597 ( .A(d4stg_fdiv), .B(div_shl_save[29]), .Z(N1051) );
  GTECH_AND2 C1598 ( .A(N1052), .B(div_frac_add[28]), .Z(N1053) );
  GTECH_AND2 C1599 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1052) );
  GTECH_AND2 C1601 ( .A(N1055), .B(div_frac_add_in1[28]), .Z(N1056) );
  GTECH_AND2 C1602 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1055)
         );
  GTECH_AND2 C1603 ( .A(d6stg_fdiv), .B(d6stg_frac_31), .Z(N1058) );
  GTECH_OR2 C1604 ( .A(N1065), .B(N1067), .Z(div_frac_add_in1_in[28]) );
  GTECH_OR2 C1605 ( .A(N1062), .B(N1064), .Z(N1065) );
  GTECH_OR2 C1606 ( .A(N1059), .B(N1061), .Z(N1062) );
  GTECH_AND2 C1607 ( .A(d4stg_fdiv), .B(div_shl_save[28]), .Z(N1059) );
  GTECH_AND2 C1608 ( .A(N1060), .B(div_frac_add[27]), .Z(N1061) );
  GTECH_AND2 C1609 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1060) );
  GTECH_AND2 C1611 ( .A(N1063), .B(div_frac_add_in1[27]), .Z(N1064) );
  GTECH_AND2 C1612 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1063)
         );
  GTECH_AND2 C1613 ( .A(d6stg_fdiv), .B(N1066), .Z(N1067) );
  GTECH_AND2 C1614 ( .A(d6stg_frac_30), .B(d6stg_fdivd), .Z(N1066) );
  GTECH_OR2 C1615 ( .A(N1074), .B(N1076), .Z(div_frac_add_in1_in[27]) );
  GTECH_OR2 C1616 ( .A(N1071), .B(N1073), .Z(N1074) );
  GTECH_OR2 C1617 ( .A(N1068), .B(N1070), .Z(N1071) );
  GTECH_AND2 C1618 ( .A(d4stg_fdiv), .B(div_shl_save[27]), .Z(N1068) );
  GTECH_AND2 C1619 ( .A(N1069), .B(div_frac_add[26]), .Z(N1070) );
  GTECH_AND2 C1620 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1069) );
  GTECH_AND2 C1622 ( .A(N1072), .B(div_frac_add_in1[26]), .Z(N1073) );
  GTECH_AND2 C1623 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1072)
         );
  GTECH_AND2 C1624 ( .A(d6stg_fdiv), .B(N1075), .Z(N1076) );
  GTECH_AND2 C1625 ( .A(d6stg_frac_29), .B(d6stg_fdivd), .Z(N1075) );
  GTECH_OR2 C1626 ( .A(N1083), .B(N1085), .Z(div_frac_add_in1_in[26]) );
  GTECH_OR2 C1627 ( .A(N1080), .B(N1082), .Z(N1083) );
  GTECH_OR2 C1628 ( .A(N1077), .B(N1079), .Z(N1080) );
  GTECH_AND2 C1629 ( .A(d4stg_fdiv), .B(div_shl_save[26]), .Z(N1077) );
  GTECH_AND2 C1630 ( .A(N1078), .B(div_frac_add[25]), .Z(N1079) );
  GTECH_AND2 C1631 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1078) );
  GTECH_AND2 C1633 ( .A(N1081), .B(div_frac_add_in1[25]), .Z(N1082) );
  GTECH_AND2 C1634 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1081)
         );
  GTECH_AND2 C1635 ( .A(d6stg_fdiv), .B(N1084), .Z(N1085) );
  GTECH_AND2 C1636 ( .A(d6stg_frac[28]), .B(d6stg_fdivd), .Z(N1084) );
  GTECH_OR2 C1637 ( .A(N1092), .B(N1094), .Z(div_frac_add_in1_in[25]) );
  GTECH_OR2 C1638 ( .A(N1089), .B(N1091), .Z(N1092) );
  GTECH_OR2 C1639 ( .A(N1086), .B(N1088), .Z(N1089) );
  GTECH_AND2 C1640 ( .A(d4stg_fdiv), .B(div_shl_save[25]), .Z(N1086) );
  GTECH_AND2 C1641 ( .A(N1087), .B(div_frac_add[24]), .Z(N1088) );
  GTECH_AND2 C1642 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1087) );
  GTECH_AND2 C1644 ( .A(N1090), .B(div_frac_add_in1[24]), .Z(N1091) );
  GTECH_AND2 C1645 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1090)
         );
  GTECH_AND2 C1646 ( .A(d6stg_fdiv), .B(N1093), .Z(N1094) );
  GTECH_AND2 C1647 ( .A(d6stg_frac[27]), .B(d6stg_fdivd), .Z(N1093) );
  GTECH_OR2 C1648 ( .A(N1101), .B(N1103), .Z(div_frac_add_in1_in[24]) );
  GTECH_OR2 C1649 ( .A(N1098), .B(N1100), .Z(N1101) );
  GTECH_OR2 C1650 ( .A(N1095), .B(N1097), .Z(N1098) );
  GTECH_AND2 C1651 ( .A(d4stg_fdiv), .B(div_shl_save[24]), .Z(N1095) );
  GTECH_AND2 C1652 ( .A(N1096), .B(div_frac_add[23]), .Z(N1097) );
  GTECH_AND2 C1653 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1096) );
  GTECH_AND2 C1655 ( .A(N1099), .B(div_frac_add_in1[23]), .Z(N1100) );
  GTECH_AND2 C1656 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1099)
         );
  GTECH_AND2 C1657 ( .A(d6stg_fdiv), .B(N1102), .Z(N1103) );
  GTECH_AND2 C1658 ( .A(d6stg_frac[26]), .B(d6stg_fdivd), .Z(N1102) );
  GTECH_OR2 C1659 ( .A(N1110), .B(N1112), .Z(div_frac_add_in1_in[23]) );
  GTECH_OR2 C1660 ( .A(N1107), .B(N1109), .Z(N1110) );
  GTECH_OR2 C1661 ( .A(N1104), .B(N1106), .Z(N1107) );
  GTECH_AND2 C1662 ( .A(d4stg_fdiv), .B(div_shl_save[23]), .Z(N1104) );
  GTECH_AND2 C1663 ( .A(N1105), .B(div_frac_add[22]), .Z(N1106) );
  GTECH_AND2 C1664 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1105) );
  GTECH_AND2 C1666 ( .A(N1108), .B(div_frac_add_in1[22]), .Z(N1109) );
  GTECH_AND2 C1667 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1108)
         );
  GTECH_AND2 C1668 ( .A(d6stg_fdiv), .B(N1111), .Z(N1112) );
  GTECH_AND2 C1669 ( .A(d6stg_frac[25]), .B(d6stg_fdivd), .Z(N1111) );
  GTECH_OR2 C1670 ( .A(N1119), .B(N1121), .Z(div_frac_add_in1_in[22]) );
  GTECH_OR2 C1671 ( .A(N1116), .B(N1118), .Z(N1119) );
  GTECH_OR2 C1672 ( .A(N1113), .B(N1115), .Z(N1116) );
  GTECH_AND2 C1673 ( .A(d4stg_fdiv), .B(div_shl_save[22]), .Z(N1113) );
  GTECH_AND2 C1674 ( .A(N1114), .B(div_frac_add[21]), .Z(N1115) );
  GTECH_AND2 C1675 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1114) );
  GTECH_AND2 C1677 ( .A(N1117), .B(div_frac_add_in1[21]), .Z(N1118) );
  GTECH_AND2 C1678 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1117)
         );
  GTECH_AND2 C1679 ( .A(d6stg_fdiv), .B(N1120), .Z(N1121) );
  GTECH_AND2 C1680 ( .A(d6stg_frac[24]), .B(d6stg_fdivd), .Z(N1120) );
  GTECH_OR2 C1681 ( .A(N1128), .B(N1130), .Z(div_frac_add_in1_in[21]) );
  GTECH_OR2 C1682 ( .A(N1125), .B(N1127), .Z(N1128) );
  GTECH_OR2 C1683 ( .A(N1122), .B(N1124), .Z(N1125) );
  GTECH_AND2 C1684 ( .A(d4stg_fdiv), .B(div_shl_save[21]), .Z(N1122) );
  GTECH_AND2 C1685 ( .A(N1123), .B(div_frac_add[20]), .Z(N1124) );
  GTECH_AND2 C1686 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1123) );
  GTECH_AND2 C1688 ( .A(N1126), .B(div_frac_add_in1[20]), .Z(N1127) );
  GTECH_AND2 C1689 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1126)
         );
  GTECH_AND2 C1690 ( .A(d6stg_fdiv), .B(N1129), .Z(N1130) );
  GTECH_AND2 C1691 ( .A(d6stg_frac[23]), .B(d6stg_fdivd), .Z(N1129) );
  GTECH_OR2 C1692 ( .A(N1137), .B(N1139), .Z(div_frac_add_in1_in[20]) );
  GTECH_OR2 C1693 ( .A(N1134), .B(N1136), .Z(N1137) );
  GTECH_OR2 C1694 ( .A(N1131), .B(N1133), .Z(N1134) );
  GTECH_AND2 C1695 ( .A(d4stg_fdiv), .B(div_shl_save[20]), .Z(N1131) );
  GTECH_AND2 C1696 ( .A(N1132), .B(div_frac_add[19]), .Z(N1133) );
  GTECH_AND2 C1697 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1132) );
  GTECH_AND2 C1699 ( .A(N1135), .B(div_frac_add_in1[19]), .Z(N1136) );
  GTECH_AND2 C1700 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1135)
         );
  GTECH_AND2 C1701 ( .A(d6stg_fdiv), .B(N1138), .Z(N1139) );
  GTECH_AND2 C1702 ( .A(d6stg_frac[22]), .B(d6stg_fdivd), .Z(N1138) );
  GTECH_OR2 C1703 ( .A(N1146), .B(N1148), .Z(div_frac_add_in1_in[19]) );
  GTECH_OR2 C1704 ( .A(N1143), .B(N1145), .Z(N1146) );
  GTECH_OR2 C1705 ( .A(N1140), .B(N1142), .Z(N1143) );
  GTECH_AND2 C1706 ( .A(d4stg_fdiv), .B(div_shl_save[19]), .Z(N1140) );
  GTECH_AND2 C1707 ( .A(N1141), .B(div_frac_add[18]), .Z(N1142) );
  GTECH_AND2 C1708 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1141) );
  GTECH_AND2 C1710 ( .A(N1144), .B(div_frac_add_in1[18]), .Z(N1145) );
  GTECH_AND2 C1711 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1144)
         );
  GTECH_AND2 C1712 ( .A(d6stg_fdiv), .B(N1147), .Z(N1148) );
  GTECH_AND2 C1713 ( .A(d6stg_frac[21]), .B(d6stg_fdivd), .Z(N1147) );
  GTECH_OR2 C1714 ( .A(N1155), .B(N1157), .Z(div_frac_add_in1_in[18]) );
  GTECH_OR2 C1715 ( .A(N1152), .B(N1154), .Z(N1155) );
  GTECH_OR2 C1716 ( .A(N1149), .B(N1151), .Z(N1152) );
  GTECH_AND2 C1717 ( .A(d4stg_fdiv), .B(div_shl_save[18]), .Z(N1149) );
  GTECH_AND2 C1718 ( .A(N1150), .B(div_frac_add[17]), .Z(N1151) );
  GTECH_AND2 C1719 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1150) );
  GTECH_AND2 C1721 ( .A(N1153), .B(div_frac_add_in1[17]), .Z(N1154) );
  GTECH_AND2 C1722 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1153)
         );
  GTECH_AND2 C1723 ( .A(d6stg_fdiv), .B(N1156), .Z(N1157) );
  GTECH_AND2 C1724 ( .A(d6stg_frac[20]), .B(d6stg_fdivd), .Z(N1156) );
  GTECH_OR2 C1725 ( .A(N1164), .B(N1166), .Z(div_frac_add_in1_in[17]) );
  GTECH_OR2 C1726 ( .A(N1161), .B(N1163), .Z(N1164) );
  GTECH_OR2 C1727 ( .A(N1158), .B(N1160), .Z(N1161) );
  GTECH_AND2 C1728 ( .A(d4stg_fdiv), .B(div_shl_save[17]), .Z(N1158) );
  GTECH_AND2 C1729 ( .A(N1159), .B(div_frac_add[16]), .Z(N1160) );
  GTECH_AND2 C1730 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1159) );
  GTECH_AND2 C1732 ( .A(N1162), .B(div_frac_add_in1[16]), .Z(N1163) );
  GTECH_AND2 C1733 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1162)
         );
  GTECH_AND2 C1734 ( .A(d6stg_fdiv), .B(N1165), .Z(N1166) );
  GTECH_AND2 C1735 ( .A(d6stg_frac[19]), .B(d6stg_fdivd), .Z(N1165) );
  GTECH_OR2 C1736 ( .A(N1173), .B(N1175), .Z(div_frac_add_in1_in[16]) );
  GTECH_OR2 C1737 ( .A(N1170), .B(N1172), .Z(N1173) );
  GTECH_OR2 C1738 ( .A(N1167), .B(N1169), .Z(N1170) );
  GTECH_AND2 C1739 ( .A(d4stg_fdiv), .B(div_shl_save[16]), .Z(N1167) );
  GTECH_AND2 C1740 ( .A(N1168), .B(div_frac_add[15]), .Z(N1169) );
  GTECH_AND2 C1741 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1168) );
  GTECH_AND2 C1743 ( .A(N1171), .B(div_frac_add_in1[15]), .Z(N1172) );
  GTECH_AND2 C1744 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1171)
         );
  GTECH_AND2 C1745 ( .A(d6stg_fdiv), .B(N1174), .Z(N1175) );
  GTECH_AND2 C1746 ( .A(d6stg_frac[18]), .B(d6stg_fdivd), .Z(N1174) );
  GTECH_OR2 C1747 ( .A(N1182), .B(N1184), .Z(div_frac_add_in1_in[15]) );
  GTECH_OR2 C1748 ( .A(N1179), .B(N1181), .Z(N1182) );
  GTECH_OR2 C1749 ( .A(N1176), .B(N1178), .Z(N1179) );
  GTECH_AND2 C1750 ( .A(d4stg_fdiv), .B(div_shl_save[15]), .Z(N1176) );
  GTECH_AND2 C1751 ( .A(N1177), .B(div_frac_add[14]), .Z(N1178) );
  GTECH_AND2 C1752 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1177) );
  GTECH_AND2 C1754 ( .A(N1180), .B(div_frac_add_in1[14]), .Z(N1181) );
  GTECH_AND2 C1755 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1180)
         );
  GTECH_AND2 C1756 ( .A(d6stg_fdiv), .B(N1183), .Z(N1184) );
  GTECH_AND2 C1757 ( .A(d6stg_frac[17]), .B(d6stg_fdivd), .Z(N1183) );
  GTECH_OR2 C1758 ( .A(N1191), .B(N1193), .Z(div_frac_add_in1_in[14]) );
  GTECH_OR2 C1759 ( .A(N1188), .B(N1190), .Z(N1191) );
  GTECH_OR2 C1760 ( .A(N1185), .B(N1187), .Z(N1188) );
  GTECH_AND2 C1761 ( .A(d4stg_fdiv), .B(div_shl_save[14]), .Z(N1185) );
  GTECH_AND2 C1762 ( .A(N1186), .B(div_frac_add[13]), .Z(N1187) );
  GTECH_AND2 C1763 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1186) );
  GTECH_AND2 C1765 ( .A(N1189), .B(div_frac_add_in1[13]), .Z(N1190) );
  GTECH_AND2 C1766 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1189)
         );
  GTECH_AND2 C1767 ( .A(d6stg_fdiv), .B(N1192), .Z(N1193) );
  GTECH_AND2 C1768 ( .A(d6stg_frac[16]), .B(d6stg_fdivd), .Z(N1192) );
  GTECH_OR2 C1769 ( .A(N1200), .B(N1202), .Z(div_frac_add_in1_in[13]) );
  GTECH_OR2 C1770 ( .A(N1197), .B(N1199), .Z(N1200) );
  GTECH_OR2 C1771 ( .A(N1194), .B(N1196), .Z(N1197) );
  GTECH_AND2 C1772 ( .A(d4stg_fdiv), .B(div_shl_save[13]), .Z(N1194) );
  GTECH_AND2 C1773 ( .A(N1195), .B(div_frac_add[12]), .Z(N1196) );
  GTECH_AND2 C1774 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1195) );
  GTECH_AND2 C1776 ( .A(N1198), .B(div_frac_add_in1[12]), .Z(N1199) );
  GTECH_AND2 C1777 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1198)
         );
  GTECH_AND2 C1778 ( .A(d6stg_fdiv), .B(N1201), .Z(N1202) );
  GTECH_AND2 C1779 ( .A(d6stg_frac[15]), .B(d6stg_fdivd), .Z(N1201) );
  GTECH_OR2 C1780 ( .A(N1209), .B(N1211), .Z(div_frac_add_in1_in[12]) );
  GTECH_OR2 C1781 ( .A(N1206), .B(N1208), .Z(N1209) );
  GTECH_OR2 C1782 ( .A(N1203), .B(N1205), .Z(N1206) );
  GTECH_AND2 C1783 ( .A(d4stg_fdiv), .B(div_shl_save[12]), .Z(N1203) );
  GTECH_AND2 C1784 ( .A(N1204), .B(div_frac_add[11]), .Z(N1205) );
  GTECH_AND2 C1785 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1204) );
  GTECH_AND2 C1787 ( .A(N1207), .B(div_frac_add_in1[11]), .Z(N1208) );
  GTECH_AND2 C1788 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1207)
         );
  GTECH_AND2 C1789 ( .A(d6stg_fdiv), .B(N1210), .Z(N1211) );
  GTECH_AND2 C1790 ( .A(d6stg_frac[14]), .B(d6stg_fdivd), .Z(N1210) );
  GTECH_OR2 C1791 ( .A(N1218), .B(N1220), .Z(div_frac_add_in1_in[11]) );
  GTECH_OR2 C1792 ( .A(N1215), .B(N1217), .Z(N1218) );
  GTECH_OR2 C1793 ( .A(N1212), .B(N1214), .Z(N1215) );
  GTECH_AND2 C1794 ( .A(d4stg_fdiv), .B(div_shl_save[11]), .Z(N1212) );
  GTECH_AND2 C1795 ( .A(N1213), .B(div_frac_add[10]), .Z(N1214) );
  GTECH_AND2 C1796 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1213) );
  GTECH_AND2 C1798 ( .A(N1216), .B(div_frac_add_in1[10]), .Z(N1217) );
  GTECH_AND2 C1799 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1216)
         );
  GTECH_AND2 C1800 ( .A(d6stg_fdiv), .B(N1219), .Z(N1220) );
  GTECH_AND2 C1801 ( .A(d6stg_frac[13]), .B(d6stg_fdivd), .Z(N1219) );
  GTECH_OR2 C1802 ( .A(N1227), .B(N1229), .Z(div_frac_add_in1_in[10]) );
  GTECH_OR2 C1803 ( .A(N1224), .B(N1226), .Z(N1227) );
  GTECH_OR2 C1804 ( .A(N1221), .B(N1223), .Z(N1224) );
  GTECH_AND2 C1805 ( .A(d4stg_fdiv), .B(div_shl_save[10]), .Z(N1221) );
  GTECH_AND2 C1806 ( .A(N1222), .B(div_frac_add[9]), .Z(N1223) );
  GTECH_AND2 C1807 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1222) );
  GTECH_AND2 C1809 ( .A(N1225), .B(div_frac_add_in1[9]), .Z(N1226) );
  GTECH_AND2 C1810 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1225)
         );
  GTECH_AND2 C1811 ( .A(d6stg_fdiv), .B(N1228), .Z(N1229) );
  GTECH_AND2 C1812 ( .A(d6stg_frac[12]), .B(d6stg_fdivd), .Z(N1228) );
  GTECH_OR2 C1813 ( .A(N1236), .B(N1238), .Z(div_frac_add_in1_in[9]) );
  GTECH_OR2 C1814 ( .A(N1233), .B(N1235), .Z(N1236) );
  GTECH_OR2 C1815 ( .A(N1230), .B(N1232), .Z(N1233) );
  GTECH_AND2 C1816 ( .A(d4stg_fdiv), .B(div_shl_save[9]), .Z(N1230) );
  GTECH_AND2 C1817 ( .A(N1231), .B(div_frac_add[8]), .Z(N1232) );
  GTECH_AND2 C1818 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1231) );
  GTECH_AND2 C1820 ( .A(N1234), .B(div_frac_add_in1[8]), .Z(N1235) );
  GTECH_AND2 C1821 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1234)
         );
  GTECH_AND2 C1822 ( .A(d6stg_fdiv), .B(N1237), .Z(N1238) );
  GTECH_AND2 C1823 ( .A(d6stg_frac[11]), .B(d6stg_fdivd), .Z(N1237) );
  GTECH_OR2 C1824 ( .A(N1245), .B(N1247), .Z(div_frac_add_in1_in[8]) );
  GTECH_OR2 C1825 ( .A(N1242), .B(N1244), .Z(N1245) );
  GTECH_OR2 C1826 ( .A(N1239), .B(N1241), .Z(N1242) );
  GTECH_AND2 C1827 ( .A(d4stg_fdiv), .B(div_shl_save[8]), .Z(N1239) );
  GTECH_AND2 C1828 ( .A(N1240), .B(div_frac_add[7]), .Z(N1241) );
  GTECH_AND2 C1829 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1240) );
  GTECH_AND2 C1831 ( .A(N1243), .B(div_frac_add_in1[7]), .Z(N1244) );
  GTECH_AND2 C1832 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1243)
         );
  GTECH_AND2 C1833 ( .A(d6stg_fdiv), .B(N1246), .Z(N1247) );
  GTECH_AND2 C1834 ( .A(d6stg_frac[10]), .B(d6stg_fdivd), .Z(N1246) );
  GTECH_OR2 C1835 ( .A(N1254), .B(N1256), .Z(div_frac_add_in1_in[7]) );
  GTECH_OR2 C1836 ( .A(N1251), .B(N1253), .Z(N1254) );
  GTECH_OR2 C1837 ( .A(N1248), .B(N1250), .Z(N1251) );
  GTECH_AND2 C1838 ( .A(d4stg_fdiv), .B(div_shl_save[7]), .Z(N1248) );
  GTECH_AND2 C1839 ( .A(N1249), .B(div_frac_add[6]), .Z(N1250) );
  GTECH_AND2 C1840 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1249) );
  GTECH_AND2 C1842 ( .A(N1252), .B(div_frac_add_in1[6]), .Z(N1253) );
  GTECH_AND2 C1843 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1252)
         );
  GTECH_AND2 C1844 ( .A(d6stg_fdiv), .B(N1255), .Z(N1256) );
  GTECH_AND2 C1845 ( .A(d6stg_frac[9]), .B(d6stg_fdivd), .Z(N1255) );
  GTECH_OR2 C1846 ( .A(N1263), .B(N1265), .Z(div_frac_add_in1_in[6]) );
  GTECH_OR2 C1847 ( .A(N1260), .B(N1262), .Z(N1263) );
  GTECH_OR2 C1848 ( .A(N1257), .B(N1259), .Z(N1260) );
  GTECH_AND2 C1849 ( .A(d4stg_fdiv), .B(div_shl_save[6]), .Z(N1257) );
  GTECH_AND2 C1850 ( .A(N1258), .B(div_frac_add[5]), .Z(N1259) );
  GTECH_AND2 C1851 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1258) );
  GTECH_AND2 C1853 ( .A(N1261), .B(div_frac_add_in1[5]), .Z(N1262) );
  GTECH_AND2 C1854 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1261)
         );
  GTECH_AND2 C1855 ( .A(d6stg_fdiv), .B(N1264), .Z(N1265) );
  GTECH_AND2 C1856 ( .A(d6stg_frac[8]), .B(d6stg_fdivd), .Z(N1264) );
  GTECH_OR2 C1857 ( .A(N1272), .B(N1274), .Z(div_frac_add_in1_in[5]) );
  GTECH_OR2 C1858 ( .A(N1269), .B(N1271), .Z(N1272) );
  GTECH_OR2 C1859 ( .A(N1266), .B(N1268), .Z(N1269) );
  GTECH_AND2 C1860 ( .A(d4stg_fdiv), .B(div_shl_save[5]), .Z(N1266) );
  GTECH_AND2 C1861 ( .A(N1267), .B(div_frac_add[4]), .Z(N1268) );
  GTECH_AND2 C1862 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1267) );
  GTECH_AND2 C1864 ( .A(N1270), .B(div_frac_add_in1[4]), .Z(N1271) );
  GTECH_AND2 C1865 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1270)
         );
  GTECH_AND2 C1866 ( .A(d6stg_fdiv), .B(N1273), .Z(N1274) );
  GTECH_AND2 C1867 ( .A(d6stg_frac[7]), .B(d6stg_fdivd), .Z(N1273) );
  GTECH_OR2 C1868 ( .A(N1281), .B(N1283), .Z(div_frac_add_in1_in[4]) );
  GTECH_OR2 C1869 ( .A(N1278), .B(N1280), .Z(N1281) );
  GTECH_OR2 C1870 ( .A(N1275), .B(N1277), .Z(N1278) );
  GTECH_AND2 C1871 ( .A(d4stg_fdiv), .B(div_shl_save[4]), .Z(N1275) );
  GTECH_AND2 C1872 ( .A(N1276), .B(div_frac_add[3]), .Z(N1277) );
  GTECH_AND2 C1873 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1276) );
  GTECH_AND2 C1875 ( .A(N1279), .B(div_frac_add_in1[3]), .Z(N1280) );
  GTECH_AND2 C1876 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1279)
         );
  GTECH_AND2 C1877 ( .A(d6stg_fdiv), .B(N1282), .Z(N1283) );
  GTECH_AND2 C1878 ( .A(d6stg_frac[6]), .B(d6stg_fdivd), .Z(N1282) );
  GTECH_OR2 C1879 ( .A(N1290), .B(N1292), .Z(div_frac_add_in1_in[3]) );
  GTECH_OR2 C1880 ( .A(N1287), .B(N1289), .Z(N1290) );
  GTECH_OR2 C1881 ( .A(N1284), .B(N1286), .Z(N1287) );
  GTECH_AND2 C1882 ( .A(d4stg_fdiv), .B(div_shl_save[3]), .Z(N1284) );
  GTECH_AND2 C1883 ( .A(N1285), .B(div_frac_add[2]), .Z(N1286) );
  GTECH_AND2 C1884 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1285) );
  GTECH_AND2 C1886 ( .A(N1288), .B(div_frac_add_in1[2]), .Z(N1289) );
  GTECH_AND2 C1887 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1288)
         );
  GTECH_AND2 C1888 ( .A(d6stg_fdiv), .B(N1291), .Z(N1292) );
  GTECH_AND2 C1889 ( .A(d6stg_frac[5]), .B(d6stg_fdivd), .Z(N1291) );
  GTECH_OR2 C1890 ( .A(N1299), .B(N1301), .Z(div_frac_add_in1_in[2]) );
  GTECH_OR2 C1891 ( .A(N1296), .B(N1298), .Z(N1299) );
  GTECH_OR2 C1892 ( .A(N1293), .B(N1295), .Z(N1296) );
  GTECH_AND2 C1893 ( .A(d4stg_fdiv), .B(div_shl_save[2]), .Z(N1293) );
  GTECH_AND2 C1894 ( .A(N1294), .B(div_frac_add[1]), .Z(N1295) );
  GTECH_AND2 C1895 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1294) );
  GTECH_AND2 C1897 ( .A(N1297), .B(div_frac_add_in1[1]), .Z(N1298) );
  GTECH_AND2 C1898 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1297)
         );
  GTECH_AND2 C1899 ( .A(d6stg_fdiv), .B(N1300), .Z(N1301) );
  GTECH_AND2 C1900 ( .A(d6stg_frac[4]), .B(d6stg_fdivd), .Z(N1300) );
  GTECH_OR2 C1901 ( .A(N1308), .B(N1310), .Z(div_frac_add_in1_in[1]) );
  GTECH_OR2 C1902 ( .A(N1305), .B(N1307), .Z(N1308) );
  GTECH_OR2 C1903 ( .A(N1302), .B(N1304), .Z(N1305) );
  GTECH_AND2 C1904 ( .A(d4stg_fdiv), .B(div_shl_save[1]), .Z(N1302) );
  GTECH_AND2 C1905 ( .A(N1303), .B(div_frac_add[0]), .Z(N1304) );
  GTECH_AND2 C1906 ( .A(div_frac_add_in1_add), .B(N857), .Z(N1303) );
  GTECH_AND2 C1908 ( .A(N1306), .B(div_frac_add_in1[0]), .Z(N1307) );
  GTECH_AND2 C1909 ( .A(div_frac_add_in1_add), .B(div_frac_add[54]), .Z(N1306)
         );
  GTECH_AND2 C1910 ( .A(d6stg_fdiv), .B(N1309), .Z(N1310) );
  GTECH_AND2 C1911 ( .A(d6stg_frac[3]), .B(d6stg_fdivd), .Z(N1309) );
  GTECH_OR2 C1912 ( .A(N1311), .B(N1313), .Z(div_frac_add_in1_in[0]) );
  GTECH_AND2 C1913 ( .A(d4stg_fdiv), .B(div_shl_save[0]), .Z(N1311) );
  GTECH_AND2 C1914 ( .A(d6stg_fdiv), .B(N1312), .Z(N1313) );
  GTECH_AND2 C1915 ( .A(d6stg_frac_2), .B(d6stg_fdivd), .Z(N1312) );
  GTECH_OR2 C1916 ( .A(N1366), .B(div_frac_add_in1[0]), .Z(
        div_frac_add_in1_neq_0) );
  GTECH_OR2 C1917 ( .A(N1365), .B(div_frac_add_in1[1]), .Z(N1366) );
  GTECH_OR2 C1918 ( .A(N1364), .B(div_frac_add_in1[2]), .Z(N1365) );
  GTECH_OR2 C1919 ( .A(N1363), .B(div_frac_add_in1[3]), .Z(N1364) );
  GTECH_OR2 C1920 ( .A(N1362), .B(div_frac_add_in1[4]), .Z(N1363) );
  GTECH_OR2 C1921 ( .A(N1361), .B(div_frac_add_in1[5]), .Z(N1362) );
  GTECH_OR2 C1922 ( .A(N1360), .B(div_frac_add_in1[6]), .Z(N1361) );
  GTECH_OR2 C1923 ( .A(N1359), .B(div_frac_add_in1[7]), .Z(N1360) );
  GTECH_OR2 C1924 ( .A(N1358), .B(div_frac_add_in1[8]), .Z(N1359) );
  GTECH_OR2 C1925 ( .A(N1357), .B(div_frac_add_in1[9]), .Z(N1358) );
  GTECH_OR2 C1926 ( .A(N1356), .B(div_frac_add_in1[10]), .Z(N1357) );
  GTECH_OR2 C1927 ( .A(N1355), .B(div_frac_add_in1[11]), .Z(N1356) );
  GTECH_OR2 C1928 ( .A(N1354), .B(div_frac_add_in1[12]), .Z(N1355) );
  GTECH_OR2 C1929 ( .A(N1353), .B(div_frac_add_in1[13]), .Z(N1354) );
  GTECH_OR2 C1930 ( .A(N1352), .B(div_frac_add_in1[14]), .Z(N1353) );
  GTECH_OR2 C1931 ( .A(N1351), .B(div_frac_add_in1[15]), .Z(N1352) );
  GTECH_OR2 C1932 ( .A(N1350), .B(div_frac_add_in1[16]), .Z(N1351) );
  GTECH_OR2 C1933 ( .A(N1349), .B(div_frac_add_in1[17]), .Z(N1350) );
  GTECH_OR2 C1934 ( .A(N1348), .B(div_frac_add_in1[18]), .Z(N1349) );
  GTECH_OR2 C1935 ( .A(N1347), .B(div_frac_add_in1[19]), .Z(N1348) );
  GTECH_OR2 C1936 ( .A(N1346), .B(div_frac_add_in1[20]), .Z(N1347) );
  GTECH_OR2 C1937 ( .A(N1345), .B(div_frac_add_in1[21]), .Z(N1346) );
  GTECH_OR2 C1938 ( .A(N1344), .B(div_frac_add_in1[22]), .Z(N1345) );
  GTECH_OR2 C1939 ( .A(N1343), .B(div_frac_add_in1[23]), .Z(N1344) );
  GTECH_OR2 C1940 ( .A(N1342), .B(div_frac_add_in1[24]), .Z(N1343) );
  GTECH_OR2 C1941 ( .A(N1341), .B(div_frac_add_in1[25]), .Z(N1342) );
  GTECH_OR2 C1942 ( .A(N1340), .B(div_frac_add_in1[26]), .Z(N1341) );
  GTECH_OR2 C1943 ( .A(N1339), .B(div_frac_add_in1[27]), .Z(N1340) );
  GTECH_OR2 C1944 ( .A(N1338), .B(div_frac_add_in1[28]), .Z(N1339) );
  GTECH_OR2 C1945 ( .A(N1337), .B(div_frac_add_in1[29]), .Z(N1338) );
  GTECH_OR2 C1946 ( .A(N1336), .B(div_frac_add_in1[30]), .Z(N1337) );
  GTECH_OR2 C1947 ( .A(N1335), .B(div_frac_add_in1[31]), .Z(N1336) );
  GTECH_OR2 C1948 ( .A(N1334), .B(div_frac_add_in1[32]), .Z(N1335) );
  GTECH_OR2 C1949 ( .A(N1333), .B(div_frac_add_in1[33]), .Z(N1334) );
  GTECH_OR2 C1950 ( .A(N1332), .B(div_frac_add_in1[34]), .Z(N1333) );
  GTECH_OR2 C1951 ( .A(N1331), .B(div_frac_add_in1[35]), .Z(N1332) );
  GTECH_OR2 C1952 ( .A(N1330), .B(div_frac_add_in1[36]), .Z(N1331) );
  GTECH_OR2 C1953 ( .A(N1329), .B(div_frac_add_in1[37]), .Z(N1330) );
  GTECH_OR2 C1954 ( .A(N1328), .B(div_frac_add_in1[38]), .Z(N1329) );
  GTECH_OR2 C1955 ( .A(N1327), .B(div_frac_add_in1[39]), .Z(N1328) );
  GTECH_OR2 C1956 ( .A(N1326), .B(div_frac_add_in1[40]), .Z(N1327) );
  GTECH_OR2 C1957 ( .A(N1325), .B(div_frac_add_in1[41]), .Z(N1326) );
  GTECH_OR2 C1958 ( .A(N1324), .B(div_frac_add_in1[42]), .Z(N1325) );
  GTECH_OR2 C1959 ( .A(N1323), .B(div_frac_add_in1[43]), .Z(N1324) );
  GTECH_OR2 C1960 ( .A(N1322), .B(div_frac_add_in1[44]), .Z(N1323) );
  GTECH_OR2 C1961 ( .A(N1321), .B(div_frac_add_in1[45]), .Z(N1322) );
  GTECH_OR2 C1962 ( .A(N1320), .B(div_frac_add_in1[46]), .Z(N1321) );
  GTECH_OR2 C1963 ( .A(N1319), .B(div_frac_add_in1[47]), .Z(N1320) );
  GTECH_OR2 C1964 ( .A(N1318), .B(div_frac_add_in1[48]), .Z(N1319) );
  GTECH_OR2 C1965 ( .A(N1317), .B(div_frac_add_in1[49]), .Z(N1318) );
  GTECH_OR2 C1966 ( .A(N1316), .B(div_frac_add_in1[50]), .Z(N1317) );
  GTECH_OR2 C1967 ( .A(N1315), .B(div_frac_add_in1[51]), .Z(N1316) );
  GTECH_OR2 C1968 ( .A(N1314), .B(div_frac_add_in1[52]), .Z(N1315) );
  GTECH_OR2 C1969 ( .A(div_frac_add_in1[54]), .B(div_frac_add_in1[53]), .Z(
        N1314) );
  GTECH_NOT I_161 ( .A(div_frac_add[52]), .Z(div_frac_add_52_inv) );
  GTECH_NOT I_162 ( .A(div_frac_add[52]), .Z(div_frac_add_52_inva) );
  GTECH_OR2 C1973 ( .A(N1373), .B(N1374), .Z(div_frac_out_in[54]) );
  GTECH_OR2 C1974 ( .A(N1371), .B(N1372), .Z(N1373) );
  GTECH_OR2 C1975 ( .A(N1369), .B(N1370), .Z(N1371) );
  GTECH_OR2 C1976 ( .A(N1367), .B(N1368), .Z(N1369) );
  GTECH_AND2 C1977 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[54]), .Z(
        N1367) );
  GTECH_AND2 C1978 ( .A(div_frac_out_add), .B(div_frac_add[54]), .Z(N1368) );
  GTECH_AND2 C1979 ( .A(div_frac_out_shl1_dbl), .B(div_frac_out_54_53[0]), .Z(
        N1370) );
  GTECH_AND2 C1980 ( .A(div_frac_out_shl1_sng), .B(div_frac_out_54_53[0]), .Z(
        N1372) );
  GTECH_AND2 C1981 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1374) );
  GTECH_OR2 C1982 ( .A(N1381), .B(N1382), .Z(div_frac_out_in[53]) );
  GTECH_OR2 C1983 ( .A(N1379), .B(N1380), .Z(N1381) );
  GTECH_OR2 C1984 ( .A(N1377), .B(N1378), .Z(N1379) );
  GTECH_OR2 C1985 ( .A(N1375), .B(N1376), .Z(N1377) );
  GTECH_AND2 C1986 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[53]), .Z(
        N1375) );
  GTECH_AND2 C1987 ( .A(div_frac_out_add), .B(div_frac_add[53]), .Z(N1376) );
  GTECH_AND2 C1988 ( .A(div_frac_out_shl1_dbl), .B(div_frac_out[52]), .Z(N1378) );
  GTECH_AND2 C1989 ( .A(div_frac_out_shl1_sng), .B(div_frac_out[52]), .Z(N1380) );
  GTECH_AND2 C1990 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1382) );
  GTECH_OR2 C1991 ( .A(N1389), .B(N1390), .Z(div_frac_out_in[52]) );
  GTECH_OR2 C1992 ( .A(N1387), .B(N1388), .Z(N1389) );
  GTECH_OR2 C1993 ( .A(N1385), .B(N1386), .Z(N1387) );
  GTECH_OR2 C1994 ( .A(N1383), .B(N1384), .Z(N1385) );
  GTECH_AND2 C1995 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[52]), .Z(
        N1383) );
  GTECH_AND2 C1996 ( .A(div_frac_out_add), .B(div_frac_add[52]), .Z(N1384) );
  GTECH_AND2 C1997 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[51]), .Z(
        N1386) );
  GTECH_AND2 C1998 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[51]), .Z(
        N1388) );
  GTECH_AND2 C1999 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1390) );
  GTECH_OR2 C2000 ( .A(N1397), .B(N1398), .Z(div_frac_out_in[51]) );
  GTECH_OR2 C2001 ( .A(N1395), .B(N1396), .Z(N1397) );
  GTECH_OR2 C2002 ( .A(N1393), .B(N1394), .Z(N1395) );
  GTECH_OR2 C2003 ( .A(N1391), .B(N1392), .Z(N1393) );
  GTECH_AND2 C2004 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[51]), .Z(
        N1391) );
  GTECH_AND2 C2005 ( .A(div_frac_out_add), .B(div_frac_add[51]), .Z(N1392) );
  GTECH_AND2 C2006 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[50]), .Z(
        N1394) );
  GTECH_AND2 C2007 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[50]), .Z(
        N1396) );
  GTECH_AND2 C2008 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1398) );
  GTECH_OR2 C2009 ( .A(N1405), .B(N1406), .Z(div_frac_out_in[50]) );
  GTECH_OR2 C2010 ( .A(N1403), .B(N1404), .Z(N1405) );
  GTECH_OR2 C2011 ( .A(N1401), .B(N1402), .Z(N1403) );
  GTECH_OR2 C2012 ( .A(N1399), .B(N1400), .Z(N1401) );
  GTECH_AND2 C2013 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[50]), .Z(
        N1399) );
  GTECH_AND2 C2014 ( .A(div_frac_out_add), .B(div_frac_add[50]), .Z(N1400) );
  GTECH_AND2 C2015 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[49]), .Z(
        N1402) );
  GTECH_AND2 C2016 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[49]), .Z(
        N1404) );
  GTECH_AND2 C2017 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1406) );
  GTECH_OR2 C2018 ( .A(N1413), .B(N1414), .Z(div_frac_out_in[49]) );
  GTECH_OR2 C2019 ( .A(N1411), .B(N1412), .Z(N1413) );
  GTECH_OR2 C2020 ( .A(N1409), .B(N1410), .Z(N1411) );
  GTECH_OR2 C2021 ( .A(N1407), .B(N1408), .Z(N1409) );
  GTECH_AND2 C2022 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[49]), .Z(
        N1407) );
  GTECH_AND2 C2023 ( .A(div_frac_out_add), .B(div_frac_add[49]), .Z(N1408) );
  GTECH_AND2 C2024 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[48]), .Z(
        N1410) );
  GTECH_AND2 C2025 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[48]), .Z(
        N1412) );
  GTECH_AND2 C2026 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1414) );
  GTECH_OR2 C2027 ( .A(N1421), .B(N1422), .Z(div_frac_out_in[48]) );
  GTECH_OR2 C2028 ( .A(N1419), .B(N1420), .Z(N1421) );
  GTECH_OR2 C2029 ( .A(N1417), .B(N1418), .Z(N1419) );
  GTECH_OR2 C2030 ( .A(N1415), .B(N1416), .Z(N1417) );
  GTECH_AND2 C2031 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[48]), .Z(
        N1415) );
  GTECH_AND2 C2032 ( .A(div_frac_out_add), .B(div_frac_add[48]), .Z(N1416) );
  GTECH_AND2 C2033 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[47]), .Z(
        N1418) );
  GTECH_AND2 C2034 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[47]), .Z(
        N1420) );
  GTECH_AND2 C2035 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1422) );
  GTECH_OR2 C2036 ( .A(N1429), .B(N1430), .Z(div_frac_out_in[47]) );
  GTECH_OR2 C2037 ( .A(N1427), .B(N1428), .Z(N1429) );
  GTECH_OR2 C2038 ( .A(N1425), .B(N1426), .Z(N1427) );
  GTECH_OR2 C2039 ( .A(N1423), .B(N1424), .Z(N1425) );
  GTECH_AND2 C2040 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[47]), .Z(
        N1423) );
  GTECH_AND2 C2041 ( .A(div_frac_out_add), .B(div_frac_add[47]), .Z(N1424) );
  GTECH_AND2 C2042 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[46]), .Z(
        N1426) );
  GTECH_AND2 C2043 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[46]), .Z(
        N1428) );
  GTECH_AND2 C2044 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1430) );
  GTECH_OR2 C2045 ( .A(N1437), .B(N1438), .Z(div_frac_out_in[46]) );
  GTECH_OR2 C2046 ( .A(N1435), .B(N1436), .Z(N1437) );
  GTECH_OR2 C2047 ( .A(N1433), .B(N1434), .Z(N1435) );
  GTECH_OR2 C2048 ( .A(N1431), .B(N1432), .Z(N1433) );
  GTECH_AND2 C2049 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[46]), .Z(
        N1431) );
  GTECH_AND2 C2050 ( .A(div_frac_out_add), .B(div_frac_add[46]), .Z(N1432) );
  GTECH_AND2 C2051 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[45]), .Z(
        N1434) );
  GTECH_AND2 C2052 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[45]), .Z(
        N1436) );
  GTECH_AND2 C2053 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1438) );
  GTECH_OR2 C2054 ( .A(N1445), .B(N1446), .Z(div_frac_out_in[45]) );
  GTECH_OR2 C2055 ( .A(N1443), .B(N1444), .Z(N1445) );
  GTECH_OR2 C2056 ( .A(N1441), .B(N1442), .Z(N1443) );
  GTECH_OR2 C2057 ( .A(N1439), .B(N1440), .Z(N1441) );
  GTECH_AND2 C2058 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[45]), .Z(
        N1439) );
  GTECH_AND2 C2059 ( .A(div_frac_out_add), .B(div_frac_add[45]), .Z(N1440) );
  GTECH_AND2 C2060 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[44]), .Z(
        N1442) );
  GTECH_AND2 C2061 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[44]), .Z(
        N1444) );
  GTECH_AND2 C2062 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1446) );
  GTECH_OR2 C2063 ( .A(N1453), .B(N1454), .Z(div_frac_out_in[44]) );
  GTECH_OR2 C2064 ( .A(N1451), .B(N1452), .Z(N1453) );
  GTECH_OR2 C2065 ( .A(N1449), .B(N1450), .Z(N1451) );
  GTECH_OR2 C2066 ( .A(N1447), .B(N1448), .Z(N1449) );
  GTECH_AND2 C2067 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[44]), .Z(
        N1447) );
  GTECH_AND2 C2068 ( .A(div_frac_out_add), .B(div_frac_add[44]), .Z(N1448) );
  GTECH_AND2 C2069 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[43]), .Z(
        N1450) );
  GTECH_AND2 C2070 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[43]), .Z(
        N1452) );
  GTECH_AND2 C2071 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1454) );
  GTECH_OR2 C2072 ( .A(N1461), .B(N1462), .Z(div_frac_out_in[43]) );
  GTECH_OR2 C2073 ( .A(N1459), .B(N1460), .Z(N1461) );
  GTECH_OR2 C2074 ( .A(N1457), .B(N1458), .Z(N1459) );
  GTECH_OR2 C2075 ( .A(N1455), .B(N1456), .Z(N1457) );
  GTECH_AND2 C2076 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[43]), .Z(
        N1455) );
  GTECH_AND2 C2077 ( .A(div_frac_out_add), .B(div_frac_add[43]), .Z(N1456) );
  GTECH_AND2 C2078 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[42]), .Z(
        N1458) );
  GTECH_AND2 C2079 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[42]), .Z(
        N1460) );
  GTECH_AND2 C2080 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1462) );
  GTECH_OR2 C2081 ( .A(N1469), .B(N1470), .Z(div_frac_out_in[42]) );
  GTECH_OR2 C2082 ( .A(N1467), .B(N1468), .Z(N1469) );
  GTECH_OR2 C2083 ( .A(N1465), .B(N1466), .Z(N1467) );
  GTECH_OR2 C2084 ( .A(N1463), .B(N1464), .Z(N1465) );
  GTECH_AND2 C2085 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[42]), .Z(
        N1463) );
  GTECH_AND2 C2086 ( .A(div_frac_out_add), .B(div_frac_add[42]), .Z(N1464) );
  GTECH_AND2 C2087 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[41]), .Z(
        N1466) );
  GTECH_AND2 C2088 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[41]), .Z(
        N1468) );
  GTECH_AND2 C2089 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1470) );
  GTECH_OR2 C2090 ( .A(N1477), .B(N1478), .Z(div_frac_out_in[41]) );
  GTECH_OR2 C2091 ( .A(N1475), .B(N1476), .Z(N1477) );
  GTECH_OR2 C2092 ( .A(N1473), .B(N1474), .Z(N1475) );
  GTECH_OR2 C2093 ( .A(N1471), .B(N1472), .Z(N1473) );
  GTECH_AND2 C2094 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[41]), .Z(
        N1471) );
  GTECH_AND2 C2095 ( .A(div_frac_out_add), .B(div_frac_add[41]), .Z(N1472) );
  GTECH_AND2 C2096 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[40]), .Z(
        N1474) );
  GTECH_AND2 C2097 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[40]), .Z(
        N1476) );
  GTECH_AND2 C2098 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1478) );
  GTECH_OR2 C2099 ( .A(N1485), .B(N1486), .Z(div_frac_out_in[40]) );
  GTECH_OR2 C2100 ( .A(N1483), .B(N1484), .Z(N1485) );
  GTECH_OR2 C2101 ( .A(N1481), .B(N1482), .Z(N1483) );
  GTECH_OR2 C2102 ( .A(N1479), .B(N1480), .Z(N1481) );
  GTECH_AND2 C2103 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[40]), .Z(
        N1479) );
  GTECH_AND2 C2104 ( .A(div_frac_out_add), .B(div_frac_add[40]), .Z(N1480) );
  GTECH_AND2 C2105 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[39]), .Z(
        N1482) );
  GTECH_AND2 C2106 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[39]), .Z(
        N1484) );
  GTECH_AND2 C2107 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1486) );
  GTECH_OR2 C2108 ( .A(N1493), .B(N1494), .Z(div_frac_out_in[39]) );
  GTECH_OR2 C2109 ( .A(N1491), .B(N1492), .Z(N1493) );
  GTECH_OR2 C2110 ( .A(N1489), .B(N1490), .Z(N1491) );
  GTECH_OR2 C2111 ( .A(N1487), .B(N1488), .Z(N1489) );
  GTECH_AND2 C2112 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[39]), .Z(
        N1487) );
  GTECH_AND2 C2113 ( .A(div_frac_out_add), .B(div_frac_add[39]), .Z(N1488) );
  GTECH_AND2 C2114 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[38]), .Z(
        N1490) );
  GTECH_AND2 C2115 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[38]), .Z(
        N1492) );
  GTECH_AND2 C2116 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1494) );
  GTECH_OR2 C2117 ( .A(N1501), .B(N1502), .Z(div_frac_out_in[38]) );
  GTECH_OR2 C2118 ( .A(N1499), .B(N1500), .Z(N1501) );
  GTECH_OR2 C2119 ( .A(N1497), .B(N1498), .Z(N1499) );
  GTECH_OR2 C2120 ( .A(N1495), .B(N1496), .Z(N1497) );
  GTECH_AND2 C2121 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[38]), .Z(
        N1495) );
  GTECH_AND2 C2122 ( .A(div_frac_out_add), .B(div_frac_add[38]), .Z(N1496) );
  GTECH_AND2 C2123 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[37]), .Z(
        N1498) );
  GTECH_AND2 C2124 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[37]), .Z(
        N1500) );
  GTECH_AND2 C2125 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1502) );
  GTECH_OR2 C2126 ( .A(N1509), .B(N1510), .Z(div_frac_out_in[37]) );
  GTECH_OR2 C2127 ( .A(N1507), .B(N1508), .Z(N1509) );
  GTECH_OR2 C2128 ( .A(N1505), .B(N1506), .Z(N1507) );
  GTECH_OR2 C2129 ( .A(N1503), .B(N1504), .Z(N1505) );
  GTECH_AND2 C2130 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[37]), .Z(
        N1503) );
  GTECH_AND2 C2131 ( .A(div_frac_out_add), .B(div_frac_add[37]), .Z(N1504) );
  GTECH_AND2 C2132 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[36]), .Z(
        N1506) );
  GTECH_AND2 C2133 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[36]), .Z(
        N1508) );
  GTECH_AND2 C2134 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1510) );
  GTECH_OR2 C2135 ( .A(N1517), .B(N1518), .Z(div_frac_out_in[36]) );
  GTECH_OR2 C2136 ( .A(N1515), .B(N1516), .Z(N1517) );
  GTECH_OR2 C2137 ( .A(N1513), .B(N1514), .Z(N1515) );
  GTECH_OR2 C2138 ( .A(N1511), .B(N1512), .Z(N1513) );
  GTECH_AND2 C2139 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[36]), .Z(
        N1511) );
  GTECH_AND2 C2140 ( .A(div_frac_out_add), .B(div_frac_add[36]), .Z(N1512) );
  GTECH_AND2 C2141 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[35]), .Z(
        N1514) );
  GTECH_AND2 C2142 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[35]), .Z(
        N1516) );
  GTECH_AND2 C2143 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1518) );
  GTECH_OR2 C2144 ( .A(N1525), .B(N1526), .Z(div_frac_out_in[35]) );
  GTECH_OR2 C2145 ( .A(N1523), .B(N1524), .Z(N1525) );
  GTECH_OR2 C2146 ( .A(N1521), .B(N1522), .Z(N1523) );
  GTECH_OR2 C2147 ( .A(N1519), .B(N1520), .Z(N1521) );
  GTECH_AND2 C2148 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[35]), .Z(
        N1519) );
  GTECH_AND2 C2149 ( .A(div_frac_out_add), .B(div_frac_add[35]), .Z(N1520) );
  GTECH_AND2 C2150 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[34]), .Z(
        N1522) );
  GTECH_AND2 C2151 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[34]), .Z(
        N1524) );
  GTECH_AND2 C2152 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1526) );
  GTECH_OR2 C2153 ( .A(N1533), .B(N1534), .Z(div_frac_out_in[34]) );
  GTECH_OR2 C2154 ( .A(N1531), .B(N1532), .Z(N1533) );
  GTECH_OR2 C2155 ( .A(N1529), .B(N1530), .Z(N1531) );
  GTECH_OR2 C2156 ( .A(N1527), .B(N1528), .Z(N1529) );
  GTECH_AND2 C2157 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[34]), .Z(
        N1527) );
  GTECH_AND2 C2158 ( .A(div_frac_out_add), .B(div_frac_add[34]), .Z(N1528) );
  GTECH_AND2 C2159 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[33]), .Z(
        N1530) );
  GTECH_AND2 C2160 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[33]), .Z(
        N1532) );
  GTECH_AND2 C2161 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1534) );
  GTECH_OR2 C2162 ( .A(N1541), .B(N1542), .Z(div_frac_out_in[33]) );
  GTECH_OR2 C2163 ( .A(N1539), .B(N1540), .Z(N1541) );
  GTECH_OR2 C2164 ( .A(N1537), .B(N1538), .Z(N1539) );
  GTECH_OR2 C2165 ( .A(N1535), .B(N1536), .Z(N1537) );
  GTECH_AND2 C2166 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[33]), .Z(
        N1535) );
  GTECH_AND2 C2167 ( .A(div_frac_out_add), .B(div_frac_add[33]), .Z(N1536) );
  GTECH_AND2 C2168 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[32]), .Z(
        N1538) );
  GTECH_AND2 C2169 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[32]), .Z(
        N1540) );
  GTECH_AND2 C2170 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1542) );
  GTECH_OR2 C2171 ( .A(N1549), .B(N1550), .Z(div_frac_out_in[32]) );
  GTECH_OR2 C2172 ( .A(N1547), .B(N1548), .Z(N1549) );
  GTECH_OR2 C2173 ( .A(N1545), .B(N1546), .Z(N1547) );
  GTECH_OR2 C2174 ( .A(N1543), .B(N1544), .Z(N1545) );
  GTECH_AND2 C2175 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[32]), .Z(
        N1543) );
  GTECH_AND2 C2176 ( .A(div_frac_out_add), .B(div_frac_add[32]), .Z(N1544) );
  GTECH_AND2 C2177 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[31]), .Z(
        N1546) );
  GTECH_AND2 C2178 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[31]), .Z(
        N1548) );
  GTECH_AND2 C2179 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1550) );
  GTECH_OR2 C2180 ( .A(N1557), .B(N1558), .Z(div_frac_out_in[31]) );
  GTECH_OR2 C2181 ( .A(N1555), .B(N1556), .Z(N1557) );
  GTECH_OR2 C2182 ( .A(N1553), .B(N1554), .Z(N1555) );
  GTECH_OR2 C2183 ( .A(N1551), .B(N1552), .Z(N1553) );
  GTECH_AND2 C2184 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[31]), .Z(
        N1551) );
  GTECH_AND2 C2185 ( .A(div_frac_out_add), .B(div_frac_add[31]), .Z(N1552) );
  GTECH_AND2 C2186 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[30]), .Z(
        N1554) );
  GTECH_AND2 C2187 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[30]), .Z(
        N1556) );
  GTECH_AND2 C2188 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1558) );
  GTECH_OR2 C2189 ( .A(N1565), .B(N1566), .Z(div_frac_out_in[30]) );
  GTECH_OR2 C2190 ( .A(N1563), .B(N1564), .Z(N1565) );
  GTECH_OR2 C2191 ( .A(N1561), .B(N1562), .Z(N1563) );
  GTECH_OR2 C2192 ( .A(N1559), .B(N1560), .Z(N1561) );
  GTECH_AND2 C2193 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[30]), .Z(
        N1559) );
  GTECH_AND2 C2194 ( .A(div_frac_out_add), .B(div_frac_add[30]), .Z(N1560) );
  GTECH_AND2 C2195 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[29]), .Z(
        N1562) );
  GTECH_AND2 C2196 ( .A(div_frac_out_shl1_sng), .B(div_frac_outa[29]), .Z(
        N1564) );
  GTECH_AND2 C2197 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1566) );
  GTECH_OR2 C2198 ( .A(N1573), .B(N1574), .Z(div_frac_out_in[29]) );
  GTECH_OR2 C2199 ( .A(N1571), .B(N1572), .Z(N1573) );
  GTECH_OR2 C2200 ( .A(N1569), .B(N1570), .Z(N1571) );
  GTECH_OR2 C2201 ( .A(N1567), .B(N1568), .Z(N1569) );
  GTECH_AND2 C2202 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[29]), .Z(
        N1567) );
  GTECH_AND2 C2203 ( .A(div_frac_out_add), .B(div_frac_add[29]), .Z(N1568) );
  GTECH_AND2 C2204 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[28]), .Z(
        N1570) );
  GTECH_AND2 C2205 ( .A(div_frac_out_shl1_sng), .B(N857), .Z(N1572) );
  GTECH_AND2 C2206 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1574) );
  GTECH_OR2 C2207 ( .A(N1579), .B(N1580), .Z(div_frac_out_in[28]) );
  GTECH_OR2 C2208 ( .A(N1577), .B(N1578), .Z(N1579) );
  GTECH_OR2 C2209 ( .A(N1575), .B(N1576), .Z(N1577) );
  GTECH_AND2 C2210 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[28]), .Z(
        N1575) );
  GTECH_AND2 C2211 ( .A(div_frac_out_add), .B(div_frac_add[28]), .Z(N1576) );
  GTECH_AND2 C2212 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[27]), .Z(
        N1578) );
  GTECH_AND2 C2213 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1580) );
  GTECH_OR2 C2214 ( .A(N1585), .B(N1586), .Z(div_frac_out_in[27]) );
  GTECH_OR2 C2215 ( .A(N1583), .B(N1584), .Z(N1585) );
  GTECH_OR2 C2216 ( .A(N1581), .B(N1582), .Z(N1583) );
  GTECH_AND2 C2217 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[27]), .Z(
        N1581) );
  GTECH_AND2 C2218 ( .A(div_frac_out_add), .B(div_frac_add[27]), .Z(N1582) );
  GTECH_AND2 C2219 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[26]), .Z(
        N1584) );
  GTECH_AND2 C2220 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1586) );
  GTECH_OR2 C2221 ( .A(N1591), .B(N1592), .Z(div_frac_out_in[26]) );
  GTECH_OR2 C2222 ( .A(N1589), .B(N1590), .Z(N1591) );
  GTECH_OR2 C2223 ( .A(N1587), .B(N1588), .Z(N1589) );
  GTECH_AND2 C2224 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[26]), .Z(
        N1587) );
  GTECH_AND2 C2225 ( .A(div_frac_out_add), .B(div_frac_add[26]), .Z(N1588) );
  GTECH_AND2 C2226 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[25]), .Z(
        N1590) );
  GTECH_AND2 C2227 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1592) );
  GTECH_OR2 C2228 ( .A(N1597), .B(N1598), .Z(div_frac_out_in[25]) );
  GTECH_OR2 C2229 ( .A(N1595), .B(N1596), .Z(N1597) );
  GTECH_OR2 C2230 ( .A(N1593), .B(N1594), .Z(N1595) );
  GTECH_AND2 C2231 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[25]), .Z(
        N1593) );
  GTECH_AND2 C2232 ( .A(div_frac_out_add), .B(div_frac_add[25]), .Z(N1594) );
  GTECH_AND2 C2233 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[24]), .Z(
        N1596) );
  GTECH_AND2 C2234 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1598) );
  GTECH_OR2 C2235 ( .A(N1603), .B(N1604), .Z(div_frac_out_in[24]) );
  GTECH_OR2 C2236 ( .A(N1601), .B(N1602), .Z(N1603) );
  GTECH_OR2 C2237 ( .A(N1599), .B(N1600), .Z(N1601) );
  GTECH_AND2 C2238 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[24]), .Z(
        N1599) );
  GTECH_AND2 C2239 ( .A(div_frac_out_add), .B(div_frac_add[24]), .Z(N1600) );
  GTECH_AND2 C2240 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[23]), .Z(
        N1602) );
  GTECH_AND2 C2241 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1604) );
  GTECH_OR2 C2242 ( .A(N1609), .B(N1610), .Z(div_frac_out_in[23]) );
  GTECH_OR2 C2243 ( .A(N1607), .B(N1608), .Z(N1609) );
  GTECH_OR2 C2244 ( .A(N1605), .B(N1606), .Z(N1607) );
  GTECH_AND2 C2245 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[23]), .Z(
        N1605) );
  GTECH_AND2 C2246 ( .A(div_frac_out_add), .B(div_frac_add[23]), .Z(N1606) );
  GTECH_AND2 C2247 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[22]), .Z(
        N1608) );
  GTECH_AND2 C2248 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1610) );
  GTECH_OR2 C2249 ( .A(N1615), .B(N1616), .Z(div_frac_out_in[22]) );
  GTECH_OR2 C2250 ( .A(N1613), .B(N1614), .Z(N1615) );
  GTECH_OR2 C2251 ( .A(N1611), .B(N1612), .Z(N1613) );
  GTECH_AND2 C2252 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[22]), .Z(
        N1611) );
  GTECH_AND2 C2253 ( .A(div_frac_out_add), .B(div_frac_add[22]), .Z(N1612) );
  GTECH_AND2 C2254 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[21]), .Z(
        N1614) );
  GTECH_AND2 C2255 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1616) );
  GTECH_OR2 C2256 ( .A(N1621), .B(N1622), .Z(div_frac_out_in[21]) );
  GTECH_OR2 C2257 ( .A(N1619), .B(N1620), .Z(N1621) );
  GTECH_OR2 C2258 ( .A(N1617), .B(N1618), .Z(N1619) );
  GTECH_AND2 C2259 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[21]), .Z(
        N1617) );
  GTECH_AND2 C2260 ( .A(div_frac_out_add), .B(div_frac_add[21]), .Z(N1618) );
  GTECH_AND2 C2261 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[20]), .Z(
        N1620) );
  GTECH_AND2 C2262 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1622) );
  GTECH_OR2 C2263 ( .A(N1627), .B(N1628), .Z(div_frac_out_in[20]) );
  GTECH_OR2 C2264 ( .A(N1625), .B(N1626), .Z(N1627) );
  GTECH_OR2 C2265 ( .A(N1623), .B(N1624), .Z(N1625) );
  GTECH_AND2 C2266 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[20]), .Z(
        N1623) );
  GTECH_AND2 C2267 ( .A(div_frac_out_add), .B(div_frac_add[20]), .Z(N1624) );
  GTECH_AND2 C2268 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[19]), .Z(
        N1626) );
  GTECH_AND2 C2269 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1628) );
  GTECH_OR2 C2270 ( .A(N1633), .B(N1634), .Z(div_frac_out_in[19]) );
  GTECH_OR2 C2271 ( .A(N1631), .B(N1632), .Z(N1633) );
  GTECH_OR2 C2272 ( .A(N1629), .B(N1630), .Z(N1631) );
  GTECH_AND2 C2273 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[19]), .Z(
        N1629) );
  GTECH_AND2 C2274 ( .A(div_frac_out_add), .B(div_frac_add[19]), .Z(N1630) );
  GTECH_AND2 C2275 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[18]), .Z(
        N1632) );
  GTECH_AND2 C2276 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1634) );
  GTECH_OR2 C2277 ( .A(N1639), .B(N1640), .Z(div_frac_out_in[18]) );
  GTECH_OR2 C2278 ( .A(N1637), .B(N1638), .Z(N1639) );
  GTECH_OR2 C2279 ( .A(N1635), .B(N1636), .Z(N1637) );
  GTECH_AND2 C2280 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[18]), .Z(
        N1635) );
  GTECH_AND2 C2281 ( .A(div_frac_out_add), .B(div_frac_add[18]), .Z(N1636) );
  GTECH_AND2 C2282 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[17]), .Z(
        N1638) );
  GTECH_AND2 C2283 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1640) );
  GTECH_OR2 C2284 ( .A(N1645), .B(N1646), .Z(div_frac_out_in[17]) );
  GTECH_OR2 C2285 ( .A(N1643), .B(N1644), .Z(N1645) );
  GTECH_OR2 C2286 ( .A(N1641), .B(N1642), .Z(N1643) );
  GTECH_AND2 C2287 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[17]), .Z(
        N1641) );
  GTECH_AND2 C2288 ( .A(div_frac_out_add), .B(div_frac_add[17]), .Z(N1642) );
  GTECH_AND2 C2289 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[16]), .Z(
        N1644) );
  GTECH_AND2 C2290 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1646) );
  GTECH_OR2 C2291 ( .A(N1651), .B(N1652), .Z(div_frac_out_in[16]) );
  GTECH_OR2 C2292 ( .A(N1649), .B(N1650), .Z(N1651) );
  GTECH_OR2 C2293 ( .A(N1647), .B(N1648), .Z(N1649) );
  GTECH_AND2 C2294 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[16]), .Z(
        N1647) );
  GTECH_AND2 C2295 ( .A(div_frac_out_add), .B(div_frac_add[16]), .Z(N1648) );
  GTECH_AND2 C2296 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[15]), .Z(
        N1650) );
  GTECH_AND2 C2297 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1652) );
  GTECH_OR2 C2298 ( .A(N1657), .B(N1658), .Z(div_frac_out_in[15]) );
  GTECH_OR2 C2299 ( .A(N1655), .B(N1656), .Z(N1657) );
  GTECH_OR2 C2300 ( .A(N1653), .B(N1654), .Z(N1655) );
  GTECH_AND2 C2301 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[15]), .Z(
        N1653) );
  GTECH_AND2 C2302 ( .A(div_frac_out_add), .B(div_frac_add[15]), .Z(N1654) );
  GTECH_AND2 C2303 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[14]), .Z(
        N1656) );
  GTECH_AND2 C2304 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1658) );
  GTECH_OR2 C2305 ( .A(N1663), .B(N1664), .Z(div_frac_out_in[14]) );
  GTECH_OR2 C2306 ( .A(N1661), .B(N1662), .Z(N1663) );
  GTECH_OR2 C2307 ( .A(N1659), .B(N1660), .Z(N1661) );
  GTECH_AND2 C2308 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[14]), .Z(
        N1659) );
  GTECH_AND2 C2309 ( .A(div_frac_out_add), .B(div_frac_add[14]), .Z(N1660) );
  GTECH_AND2 C2310 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[13]), .Z(
        N1662) );
  GTECH_AND2 C2311 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1664) );
  GTECH_OR2 C2312 ( .A(N1669), .B(N1670), .Z(div_frac_out_in[13]) );
  GTECH_OR2 C2313 ( .A(N1667), .B(N1668), .Z(N1669) );
  GTECH_OR2 C2314 ( .A(N1665), .B(N1666), .Z(N1667) );
  GTECH_AND2 C2315 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[13]), .Z(
        N1665) );
  GTECH_AND2 C2316 ( .A(div_frac_out_add), .B(div_frac_add[13]), .Z(N1666) );
  GTECH_AND2 C2317 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[12]), .Z(
        N1668) );
  GTECH_AND2 C2318 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1670) );
  GTECH_OR2 C2319 ( .A(N1675), .B(N1676), .Z(div_frac_out_in[12]) );
  GTECH_OR2 C2320 ( .A(N1673), .B(N1674), .Z(N1675) );
  GTECH_OR2 C2321 ( .A(N1671), .B(N1672), .Z(N1673) );
  GTECH_AND2 C2322 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[12]), .Z(
        N1671) );
  GTECH_AND2 C2323 ( .A(div_frac_out_add), .B(div_frac_add[12]), .Z(N1672) );
  GTECH_AND2 C2324 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[11]), .Z(
        N1674) );
  GTECH_AND2 C2325 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1676) );
  GTECH_OR2 C2326 ( .A(N1681), .B(N1682), .Z(div_frac_out_in[11]) );
  GTECH_OR2 C2327 ( .A(N1679), .B(N1680), .Z(N1681) );
  GTECH_OR2 C2328 ( .A(N1677), .B(N1678), .Z(N1679) );
  GTECH_AND2 C2329 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[11]), .Z(
        N1677) );
  GTECH_AND2 C2330 ( .A(div_frac_out_add), .B(div_frac_add[11]), .Z(N1678) );
  GTECH_AND2 C2331 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[10]), .Z(
        N1680) );
  GTECH_AND2 C2332 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1682) );
  GTECH_OR2 C2333 ( .A(N1687), .B(N1688), .Z(div_frac_out_in[10]) );
  GTECH_OR2 C2334 ( .A(N1685), .B(N1686), .Z(N1687) );
  GTECH_OR2 C2335 ( .A(N1683), .B(N1684), .Z(N1685) );
  GTECH_AND2 C2336 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[10]), .Z(
        N1683) );
  GTECH_AND2 C2337 ( .A(div_frac_out_add), .B(div_frac_add[10]), .Z(N1684) );
  GTECH_AND2 C2338 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[9]), .Z(N1686) );
  GTECH_AND2 C2339 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1688) );
  GTECH_OR2 C2340 ( .A(N1693), .B(N1694), .Z(div_frac_out_in[9]) );
  GTECH_OR2 C2341 ( .A(N1691), .B(N1692), .Z(N1693) );
  GTECH_OR2 C2342 ( .A(N1689), .B(N1690), .Z(N1691) );
  GTECH_AND2 C2343 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[9]), .Z(
        N1689) );
  GTECH_AND2 C2344 ( .A(div_frac_out_add), .B(div_frac_add[9]), .Z(N1690) );
  GTECH_AND2 C2345 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[8]), .Z(N1692) );
  GTECH_AND2 C2346 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1694) );
  GTECH_OR2 C2347 ( .A(N1699), .B(N1700), .Z(div_frac_out_in[8]) );
  GTECH_OR2 C2348 ( .A(N1697), .B(N1698), .Z(N1699) );
  GTECH_OR2 C2349 ( .A(N1695), .B(N1696), .Z(N1697) );
  GTECH_AND2 C2350 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[8]), .Z(
        N1695) );
  GTECH_AND2 C2351 ( .A(div_frac_out_add), .B(div_frac_add[8]), .Z(N1696) );
  GTECH_AND2 C2352 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[7]), .Z(N1698) );
  GTECH_AND2 C2353 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1700) );
  GTECH_OR2 C2354 ( .A(N1705), .B(N1706), .Z(div_frac_out_in[7]) );
  GTECH_OR2 C2355 ( .A(N1703), .B(N1704), .Z(N1705) );
  GTECH_OR2 C2356 ( .A(N1701), .B(N1702), .Z(N1703) );
  GTECH_AND2 C2357 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[7]), .Z(
        N1701) );
  GTECH_AND2 C2358 ( .A(div_frac_out_add), .B(div_frac_add[7]), .Z(N1702) );
  GTECH_AND2 C2359 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[6]), .Z(N1704) );
  GTECH_AND2 C2360 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1706) );
  GTECH_OR2 C2361 ( .A(N1711), .B(N1712), .Z(div_frac_out_in[6]) );
  GTECH_OR2 C2362 ( .A(N1709), .B(N1710), .Z(N1711) );
  GTECH_OR2 C2363 ( .A(N1707), .B(N1708), .Z(N1709) );
  GTECH_AND2 C2364 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[6]), .Z(
        N1707) );
  GTECH_AND2 C2365 ( .A(div_frac_out_add), .B(div_frac_add[6]), .Z(N1708) );
  GTECH_AND2 C2366 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[5]), .Z(N1710) );
  GTECH_AND2 C2367 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1712) );
  GTECH_OR2 C2368 ( .A(N1717), .B(N1718), .Z(div_frac_out_in[5]) );
  GTECH_OR2 C2369 ( .A(N1715), .B(N1716), .Z(N1717) );
  GTECH_OR2 C2370 ( .A(N1713), .B(N1714), .Z(N1715) );
  GTECH_AND2 C2371 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[5]), .Z(
        N1713) );
  GTECH_AND2 C2372 ( .A(div_frac_out_add), .B(div_frac_add[5]), .Z(N1714) );
  GTECH_AND2 C2373 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[4]), .Z(N1716) );
  GTECH_AND2 C2374 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1718) );
  GTECH_OR2 C2375 ( .A(N1723), .B(N1724), .Z(div_frac_out_in[4]) );
  GTECH_OR2 C2376 ( .A(N1721), .B(N1722), .Z(N1723) );
  GTECH_OR2 C2377 ( .A(N1719), .B(N1720), .Z(N1721) );
  GTECH_AND2 C2378 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[4]), .Z(
        N1719) );
  GTECH_AND2 C2379 ( .A(div_frac_out_add), .B(div_frac_add[4]), .Z(N1720) );
  GTECH_AND2 C2380 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[3]), .Z(N1722) );
  GTECH_AND2 C2381 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1724) );
  GTECH_OR2 C2382 ( .A(N1729), .B(N1730), .Z(div_frac_out_in[3]) );
  GTECH_OR2 C2383 ( .A(N1727), .B(N1728), .Z(N1729) );
  GTECH_OR2 C2384 ( .A(N1725), .B(N1726), .Z(N1727) );
  GTECH_AND2 C2385 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[3]), .Z(
        N1725) );
  GTECH_AND2 C2386 ( .A(div_frac_out_add), .B(div_frac_add[3]), .Z(N1726) );
  GTECH_AND2 C2387 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[2]), .Z(N1728) );
  GTECH_AND2 C2388 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1730) );
  GTECH_OR2 C2389 ( .A(N1735), .B(N1736), .Z(div_frac_out_in[2]) );
  GTECH_OR2 C2390 ( .A(N1733), .B(N1734), .Z(N1735) );
  GTECH_OR2 C2391 ( .A(N1731), .B(N1732), .Z(N1733) );
  GTECH_AND2 C2392 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[2]), .Z(
        N1731) );
  GTECH_AND2 C2393 ( .A(div_frac_out_add), .B(div_frac_add[2]), .Z(N1732) );
  GTECH_AND2 C2394 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[1]), .Z(N1734) );
  GTECH_AND2 C2395 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1736) );
  GTECH_OR2 C2396 ( .A(N1741), .B(N1742), .Z(div_frac_out_in[1]) );
  GTECH_OR2 C2397 ( .A(N1739), .B(N1740), .Z(N1741) );
  GTECH_OR2 C2398 ( .A(N1737), .B(N1738), .Z(N1739) );
  GTECH_AND2 C2399 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[1]), .Z(
        N1737) );
  GTECH_AND2 C2400 ( .A(div_frac_out_add), .B(div_frac_add[1]), .Z(N1738) );
  GTECH_AND2 C2401 ( .A(div_frac_out_shl1_dbl), .B(div_frac_outa[0]), .Z(N1740) );
  GTECH_AND2 C2402 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1742) );
  GTECH_OR2 C2403 ( .A(N1747), .B(N1748), .Z(div_frac_out_in[0]) );
  GTECH_OR2 C2404 ( .A(N1745), .B(N1746), .Z(N1747) );
  GTECH_OR2 C2405 ( .A(N1743), .B(N1744), .Z(N1745) );
  GTECH_AND2 C2406 ( .A(div_frac_out_add_in1), .B(div_frac_add_in1[0]), .Z(
        N1743) );
  GTECH_AND2 C2407 ( .A(div_frac_out_add), .B(div_frac_add[0]), .Z(N1744) );
  GTECH_AND2 C2408 ( .A(div_frac_out_shl1_dbl), .B(N857), .Z(N1746) );
  GTECH_AND2 C2409 ( .A(div_frac_out_of), .B(d7stg_to_0), .Z(N1748) );
endmodule


module fpu_div ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_div, 
        div_dest_rdy, fdiv_clken_l, fdiv_clken_l_div_exp_buf1, arst_l, grst_l, 
        rclk, div_pipe_active, d1stg_step, d8stg_fdiv_in, div_id_out_in, 
        div_exc_out, d8stg_fdivd, d8stg_fdivs, div_sign_out, div_exp_outa, 
        div_frac_outa, se, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] div_id_out_in;
  output [4:0] div_exc_out;
  output [10:0] div_exp_outa;
  output [51:0] div_frac_outa;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_div, div_dest_rdy, fdiv_clken_l,
         fdiv_clken_l_div_exp_buf1, arst_l, grst_l, rclk, se, si;
  output div_pipe_active, d1stg_step, d8stg_fdiv_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, so;
  wire   div_frac_add_52_inva, div_frac_add_in1_neq_0, d6stg_frac_0,
         d6stg_frac_1, d6stg_frac_2, d6stg_frac_29, d6stg_frac_30,
         d6stg_frac_31, d1stg_snan_sng_in1, d1stg_snan_dbl_in1,
         d1stg_snan_sng_in2, d1stg_snan_dbl_in2, d1stg_dblop, d234stg_fdiv,
         d3stg_fdiv, d4stg_fdiv, d5stg_fdiva, d5stg_fdivb, d5stg_fdivs,
         d5stg_fdivd, d6stg_fdiv, d6stg_fdivs, d6stg_fdivd, d7stg_fdiv,
         d7stg_fdivd, div_norm_frac_in1_dbl_norm, div_norm_frac_in1_dbl_dnrm,
         div_norm_frac_in1_sng_norm, div_norm_frac_in1_sng_dnrm,
         div_norm_frac_in2_dbl_norm, div_norm_frac_in2_dbl_dnrm,
         div_norm_frac_in2_sng_norm, div_norm_frac_in2_sng_dnrm, div_norm_inf,
         div_norm_qnan, div_norm_zero, div_frac_add_in2_load,
         d6stg_frac_out_shl1, d6stg_frac_out_nosh, div_frac_add_in1_add,
         div_frac_add_in1_load, d7stg_rndup_inv, d7stg_to_0, d7stg_to_0_inv,
         div_frac_out_add_in1, div_frac_out_add, div_frac_out_shl1_dbl,
         div_frac_out_shl1_sng, div_frac_out_of, div_frac_out_load,
         div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl,
         div_expadd1_in2_exp_in2_sng, div_exp1_expadd1, div_exp1_0835,
         div_exp1_0118, div_exp1_zero, div_exp1_load, div_expadd2_in1_exp_out,
         div_expadd2_no_decr_inv, div_expadd2_cin, div_exp_out_expadd22_inv,
         div_exp_out_expadd2, div_exp_out_of, div_exp_out_exp_out,
         div_exp_out_load, scan_out_fpu_div_ctl, div_frac_add_52_inv,
         scan_out_fpu_div_exp_dp;
  wire   [12:0] div_exp1;
  wire   [12:0] div_exp_out;
  wire   [54:53] div_frac_out;
  wire   [12:12] div_expadd2;
  wire   [5:0] div_shl_cnt;

  fpu_div_ctl fpu_div_ctl ( .inq_in1_51(inq_in1[51]), .inq_in1_54(inq_in1[54]), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_51(inq_in2[51]), .inq_in2_54(
        inq_in2[54]), .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .inq_op(inq_op), .div_exp1(
        div_exp1), .div_dest_rdy(div_dest_rdy), .inq_rnd_mode(inq_rnd_mode), 
        .inq_id(inq_id), .inq_in1_63(inq_in1[63]), .inq_in2_63(inq_in2[63]), 
        .inq_div(inq_div), .div_exp_out(div_exp_out), .div_frac_add_52_inva(
        div_frac_add_52_inva), .div_frac_add_in1_neq_0(div_frac_add_in1_neq_0), 
        .div_frac_out_54(div_frac_out[54]), .d6stg_frac_0(d6stg_frac_0), 
        .d6stg_frac_1(d6stg_frac_1), .d6stg_frac_2(d6stg_frac_2), 
        .d6stg_frac_29(d6stg_frac_29), .d6stg_frac_30(d6stg_frac_30), 
        .d6stg_frac_31(d6stg_frac_31), .div_frac_out_53(div_frac_out[53]), 
        .div_expadd2_12(div_expadd2[12]), .arst_l(arst_l), .grst_l(grst_l), 
        .rclk(rclk), .div_pipe_active(div_pipe_active), .d1stg_snan_sng_in1(
        d1stg_snan_sng_in1), .d1stg_snan_dbl_in1(d1stg_snan_dbl_in1), 
        .d1stg_snan_sng_in2(d1stg_snan_sng_in2), .d1stg_snan_dbl_in2(
        d1stg_snan_dbl_in2), .d1stg_step(d1stg_step), .d1stg_dblop(d1stg_dblop), .d234stg_fdiv(d234stg_fdiv), .d3stg_fdiv(d3stg_fdiv), .d4stg_fdiv(d4stg_fdiv), .d5stg_fdiva(d5stg_fdiva), .d5stg_fdivb(d5stg_fdivb), .d5stg_fdivs(
        d5stg_fdivs), .d5stg_fdivd(d5stg_fdivd), .d6stg_fdiv(d6stg_fdiv), 
        .d6stg_fdivs(d6stg_fdivs), .d6stg_fdivd(d6stg_fdivd), .d7stg_fdiv(
        d7stg_fdiv), .d7stg_fdivd(d7stg_fdivd), .d8stg_fdiv_in(d8stg_fdiv_in), 
        .d8stg_fdivs(d8stg_fdivs), .d8stg_fdivd(d8stg_fdivd), .div_id_out_in(
        div_id_out_in), .div_sign_out(div_sign_out), .div_exc_out(div_exc_out), 
        .div_norm_frac_in1_dbl_norm(div_norm_frac_in1_dbl_norm), 
        .div_norm_frac_in1_dbl_dnrm(div_norm_frac_in1_dbl_dnrm), 
        .div_norm_frac_in1_sng_norm(div_norm_frac_in1_sng_norm), 
        .div_norm_frac_in1_sng_dnrm(div_norm_frac_in1_sng_dnrm), 
        .div_norm_frac_in2_dbl_norm(div_norm_frac_in2_dbl_norm), 
        .div_norm_frac_in2_dbl_dnrm(div_norm_frac_in2_dbl_dnrm), 
        .div_norm_frac_in2_sng_norm(div_norm_frac_in2_sng_norm), 
        .div_norm_frac_in2_sng_dnrm(div_norm_frac_in2_sng_dnrm), 
        .div_norm_inf(div_norm_inf), .div_norm_qnan(div_norm_qnan), 
        .div_norm_zero(div_norm_zero), .div_frac_add_in2_load(
        div_frac_add_in2_load), .d6stg_frac_out_shl1(d6stg_frac_out_shl1), 
        .d6stg_frac_out_nosh(d6stg_frac_out_nosh), .div_frac_add_in1_add(
        div_frac_add_in1_add), .div_frac_add_in1_load(div_frac_add_in1_load), 
        .d7stg_rndup_inv(d7stg_rndup_inv), .d7stg_to_0(d7stg_to_0), 
        .d7stg_to_0_inv(d7stg_to_0_inv), .div_frac_out_add_in1(
        div_frac_out_add_in1), .div_frac_out_add(div_frac_out_add), 
        .div_frac_out_shl1_dbl(div_frac_out_shl1_dbl), .div_frac_out_shl1_sng(
        div_frac_out_shl1_sng), .div_frac_out_of(div_frac_out_of), 
        .div_frac_out_load(div_frac_out_load), .div_expadd1_in1_dbl(
        div_expadd1_in1_dbl), .div_expadd1_in1_sng(div_expadd1_in1_sng), 
        .div_expadd1_in2_exp_in2_dbl(div_expadd1_in2_exp_in2_dbl), 
        .div_expadd1_in2_exp_in2_sng(div_expadd1_in2_exp_in2_sng), 
        .div_exp1_expadd1(div_exp1_expadd1), .div_exp1_0835(div_exp1_0835), 
        .div_exp1_0118(div_exp1_0118), .div_exp1_zero(div_exp1_zero), 
        .div_exp1_load(div_exp1_load), .div_expadd2_in1_exp_out(
        div_expadd2_in1_exp_out), .div_expadd2_no_decr_inv(
        div_expadd2_no_decr_inv), .div_expadd2_cin(div_expadd2_cin), 
        .div_exp_out_expadd22_inv(div_exp_out_expadd22_inv), 
        .div_exp_out_expadd2(div_exp_out_expadd2), .div_exp_out_of(
        div_exp_out_of), .div_exp_out_exp_out(div_exp_out_exp_out), 
        .div_exp_out_load(div_exp_out_load), .se(se), .si(si), .so(
        scan_out_fpu_div_ctl) );
  fpu_div_exp_dp fpu_div_exp_dp ( .inq_in1(inq_in1[62:52]), .inq_in2(
        inq_in2[62:52]), .d1stg_step(d1stg_step), .d234stg_fdiv(d234stg_fdiv), 
        .div_expadd1_in1_dbl(div_expadd1_in1_dbl), .div_expadd1_in1_sng(
        div_expadd1_in1_sng), .div_expadd1_in2_exp_in2_dbl(
        div_expadd1_in2_exp_in2_dbl), .div_expadd1_in2_exp_in2_sng(
        div_expadd1_in2_exp_in2_sng), .d3stg_fdiv(d3stg_fdiv), .d4stg_fdiv(
        d4stg_fdiv), .div_shl_cnt(div_shl_cnt), .div_exp1_expadd1(
        div_exp1_expadd1), .div_exp1_0835(div_exp1_0835), .div_exp1_0118(
        div_exp1_0118), .div_exp1_zero(div_exp1_zero), .div_exp1_load(
        div_exp1_load), .div_expadd2_in1_exp_out(div_expadd2_in1_exp_out), 
        .d5stg_fdiva(d5stg_fdiva), .d5stg_fdivd(d5stg_fdivd), .d5stg_fdivs(
        d5stg_fdivs), .d6stg_fdiv(d6stg_fdiv), .d7stg_fdiv(d7stg_fdiv), 
        .div_expadd2_no_decr_inv(div_expadd2_no_decr_inv), .div_expadd2_cin(
        div_expadd2_cin), .div_exp_out_expadd2(div_exp_out_expadd2), 
        .div_exp_out_expadd22_inv(div_exp_out_expadd22_inv), .div_exp_out_of(
        div_exp_out_of), .d7stg_to_0_inv(d7stg_to_0_inv), .d7stg_fdivd(
        d7stg_fdivd), .div_exp_out_exp_out(div_exp_out_exp_out), 
        .d7stg_rndup_inv(d7stg_rndup_inv), .div_frac_add_52_inv(
        div_frac_add_52_inv), .div_exp_out_load(div_exp_out_load), 
        .fdiv_clken_l(fdiv_clken_l_div_exp_buf1), .rclk(rclk), .div_exp1(
        div_exp1), .div_expadd2_12(div_expadd2[12]), .div_exp_out(div_exp_out), 
        .div_exp_outa(div_exp_outa), .se(se), .si(scan_out_fpu_div_ctl), .so(
        scan_out_fpu_div_exp_dp) );
  fpu_div_frac_dp fpu_div_frac_dp ( .inq_in1(inq_in1[54:0]), .inq_in2(
        inq_in2[54:0]), .d1stg_step(d1stg_step), .div_norm_frac_in1_dbl_norm(
        div_norm_frac_in1_dbl_norm), .div_norm_frac_in1_dbl_dnrm(
        div_norm_frac_in1_dbl_dnrm), .div_norm_frac_in1_sng_norm(
        div_norm_frac_in1_sng_norm), .div_norm_frac_in1_sng_dnrm(
        div_norm_frac_in1_sng_dnrm), .div_norm_frac_in2_dbl_norm(
        div_norm_frac_in2_dbl_norm), .div_norm_frac_in2_dbl_dnrm(
        div_norm_frac_in2_dbl_dnrm), .div_norm_frac_in2_sng_norm(
        div_norm_frac_in2_sng_norm), .div_norm_frac_in2_sng_dnrm(
        div_norm_frac_in2_sng_dnrm), .div_norm_inf(div_norm_inf), 
        .div_norm_qnan(div_norm_qnan), .d1stg_dblop(d1stg_dblop), 
        .div_norm_zero(div_norm_zero), .d1stg_snan_dbl_in1(d1stg_snan_dbl_in1), 
        .d1stg_snan_sng_in1(d1stg_snan_sng_in1), .d1stg_snan_dbl_in2(
        d1stg_snan_dbl_in2), .d1stg_snan_sng_in2(d1stg_snan_sng_in2), 
        .d3stg_fdiv(d3stg_fdiv), .d6stg_fdiv(d6stg_fdiv), .d6stg_fdivd(
        d6stg_fdivd), .d6stg_fdivs(d6stg_fdivs), .div_frac_add_in2_load(
        div_frac_add_in2_load), .d6stg_frac_out_shl1(d6stg_frac_out_shl1), 
        .d6stg_frac_out_nosh(d6stg_frac_out_nosh), .d4stg_fdiv(d4stg_fdiv), 
        .div_frac_add_in1_add(div_frac_add_in1_add), .div_frac_add_in1_load(
        div_frac_add_in1_load), .d5stg_fdivb(d5stg_fdivb), 
        .div_frac_out_add_in1(div_frac_out_add_in1), .div_frac_out_add(
        div_frac_out_add), .div_frac_out_shl1_dbl(div_frac_out_shl1_dbl), 
        .div_frac_out_shl1_sng(div_frac_out_shl1_sng), .div_frac_out_of(
        div_frac_out_of), .d7stg_to_0(d7stg_to_0), .div_frac_out_load(
        div_frac_out_load), .fdiv_clken_l(fdiv_clken_l), .rclk(rclk), 
        .div_shl_cnt(div_shl_cnt), .d6stg_frac_0(d6stg_frac_0), .d6stg_frac_1(
        d6stg_frac_1), .d6stg_frac_2(d6stg_frac_2), .d6stg_frac_29(
        d6stg_frac_29), .d6stg_frac_30(d6stg_frac_30), .d6stg_frac_31(
        d6stg_frac_31), .div_frac_add_in1_neq_0(div_frac_add_in1_neq_0), 
        .div_frac_add_52_inv(div_frac_add_52_inv), .div_frac_add_52_inva(
        div_frac_add_52_inva), .div_frac_out_54_53(div_frac_out), 
        .div_frac_outa(div_frac_outa), .se(se), .si(scan_out_fpu_div_exp_dp), 
        .so(so) );
endmodule


module fpu_out_ctl ( d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, 
        div_id_out_in, m6stg_id_in, add_id_out_in, arst_l, grst_l, rclk, 
        fp_cpx_req_cq, req_thread, dest_rdy, add_dest_rdy, mul_dest_rdy, 
        div_dest_rdy, se, si, so );
  input [9:0] div_id_out_in;
  input [9:0] m6stg_id_in;
  input [9:0] add_id_out_in;
  output [7:0] fp_cpx_req_cq;
  output [1:0] req_thread;
  output [2:0] dest_rdy;
  input d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, arst_l, grst_l, rclk, se,
         si;
  output add_dest_rdy, mul_dest_rdy, div_dest_rdy, so;
  wire   out_ctl_rst_l, reset, add_req, add_req_in, add_req_step, N0, N1, N2,
         N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, net12294, net12295, net12296, net12297, net12298,
         net12299, net12300, net12301, net12302, net12303, net12304, net12305,
         net12306, net12307, net12308, net12309, net12310, net12311, net12312;
  wire   [9:0] out_id;
  wire   [1:0] dest_rdy_in;

  dffrl_async_SIZE1 dffrl_out_ctl ( .din(grst_l), .clk(rclk), .rst_l(arst_l), 
        .q(out_ctl_rst_l), .se(se), .si(net12312) );
  dffre_SIZE1 i_add_req ( .din(add_req_in), .rst(reset), .en(add_req_step), 
        .clk(rclk), .q(add_req), .se(se), .si(net12311) );
  dff_SIZE8 i_fp_cpx_req_cq ( .din(out_id[9:2]), .clk(rclk), .q(fp_cpx_req_cq), 
        .se(se), .si({net12303, net12304, net12305, net12306, net12307, 
        net12308, net12309, net12310}) );
  dff_SIZE2 i_req_thread ( .din(out_id[1:0]), .clk(rclk), .q(req_thread), .se(
        se), .si({net12301, net12302}) );
  dff_SIZE3 i_dest_rdy ( .din({d8stg_fdiv_in, dest_rdy_in}), .clk(rclk), .q(
        dest_rdy), .se(se), .si({net12298, net12299, net12300}) );
  dff_SIZE1 i_add_dest_rdy ( .din(dest_rdy_in[0]), .clk(rclk), .q(add_dest_rdy), .se(se), .si(net12297) );
  dff_SIZE1 i_mul_dest_rdy ( .din(dest_rdy_in[1]), .clk(rclk), .q(mul_dest_rdy), .se(se), .si(net12296) );
  dff_SIZE1 i_div_dest_rdy ( .din(d8stg_fdiv_in), .clk(rclk), .q(div_dest_rdy), 
        .se(se), .si(net12295) );
  GTECH_NOT I_0 ( .A(out_ctl_rst_l), .Z(reset) );
  GTECH_NOT I_1 ( .A(add_req), .Z(add_req_in) );
  GTECH_OR2 C23 ( .A(dest_rdy_in[0]), .B(dest_rdy_in[1]), .Z(add_req_step) );
  GTECH_AND2 C24 ( .A(N3), .B(N4), .Z(dest_rdy_in[1]) );
  GTECH_AND2 C25 ( .A(m6stg_fmul_in), .B(N2), .Z(N3) );
  GTECH_OR2 C26 ( .A(N0), .B(N1), .Z(N2) );
  GTECH_NOT I_2 ( .A(add_req), .Z(N0) );
  GTECH_NOT I_3 ( .A(a6stg_fadd_in), .Z(N1) );
  GTECH_NOT I_4 ( .A(d8stg_fdiv_in), .Z(N4) );
  GTECH_AND2 C30 ( .A(N7), .B(N8), .Z(dest_rdy_in[0]) );
  GTECH_AND2 C31 ( .A(a6stg_fadd_in), .B(N6), .Z(N7) );
  GTECH_OR2 C32 ( .A(add_req), .B(N5), .Z(N6) );
  GTECH_NOT I_5 ( .A(m6stg_fmul_in), .Z(N5) );
  GTECH_NOT I_6 ( .A(d8stg_fdiv_in), .Z(N8) );
  GTECH_OR2 C35 ( .A(N11), .B(N12), .Z(out_id[9]) );
  GTECH_OR2 C36 ( .A(N9), .B(N10), .Z(N11) );
  GTECH_AND2 C37 ( .A(d8stg_fdiv_in), .B(div_id_out_in[9]), .Z(N9) );
  GTECH_AND2 C38 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[9]), .Z(N10) );
  GTECH_AND2 C39 ( .A(dest_rdy_in[0]), .B(add_id_out_in[9]), .Z(N12) );
  GTECH_OR2 C40 ( .A(N15), .B(N16), .Z(out_id[8]) );
  GTECH_OR2 C41 ( .A(N13), .B(N14), .Z(N15) );
  GTECH_AND2 C42 ( .A(d8stg_fdiv_in), .B(div_id_out_in[8]), .Z(N13) );
  GTECH_AND2 C43 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[8]), .Z(N14) );
  GTECH_AND2 C44 ( .A(dest_rdy_in[0]), .B(add_id_out_in[8]), .Z(N16) );
  GTECH_OR2 C45 ( .A(N19), .B(N20), .Z(out_id[7]) );
  GTECH_OR2 C46 ( .A(N17), .B(N18), .Z(N19) );
  GTECH_AND2 C47 ( .A(d8stg_fdiv_in), .B(div_id_out_in[7]), .Z(N17) );
  GTECH_AND2 C48 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[7]), .Z(N18) );
  GTECH_AND2 C49 ( .A(dest_rdy_in[0]), .B(add_id_out_in[7]), .Z(N20) );
  GTECH_OR2 C50 ( .A(N23), .B(N24), .Z(out_id[6]) );
  GTECH_OR2 C51 ( .A(N21), .B(N22), .Z(N23) );
  GTECH_AND2 C52 ( .A(d8stg_fdiv_in), .B(div_id_out_in[6]), .Z(N21) );
  GTECH_AND2 C53 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[6]), .Z(N22) );
  GTECH_AND2 C54 ( .A(dest_rdy_in[0]), .B(add_id_out_in[6]), .Z(N24) );
  GTECH_OR2 C55 ( .A(N27), .B(N28), .Z(out_id[5]) );
  GTECH_OR2 C56 ( .A(N25), .B(N26), .Z(N27) );
  GTECH_AND2 C57 ( .A(d8stg_fdiv_in), .B(div_id_out_in[5]), .Z(N25) );
  GTECH_AND2 C58 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[5]), .Z(N26) );
  GTECH_AND2 C59 ( .A(dest_rdy_in[0]), .B(add_id_out_in[5]), .Z(N28) );
  GTECH_OR2 C60 ( .A(N31), .B(N32), .Z(out_id[4]) );
  GTECH_OR2 C61 ( .A(N29), .B(N30), .Z(N31) );
  GTECH_AND2 C62 ( .A(d8stg_fdiv_in), .B(div_id_out_in[4]), .Z(N29) );
  GTECH_AND2 C63 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[4]), .Z(N30) );
  GTECH_AND2 C64 ( .A(dest_rdy_in[0]), .B(add_id_out_in[4]), .Z(N32) );
  GTECH_OR2 C65 ( .A(N35), .B(N36), .Z(out_id[3]) );
  GTECH_OR2 C66 ( .A(N33), .B(N34), .Z(N35) );
  GTECH_AND2 C67 ( .A(d8stg_fdiv_in), .B(div_id_out_in[3]), .Z(N33) );
  GTECH_AND2 C68 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[3]), .Z(N34) );
  GTECH_AND2 C69 ( .A(dest_rdy_in[0]), .B(add_id_out_in[3]), .Z(N36) );
  GTECH_OR2 C70 ( .A(N39), .B(N40), .Z(out_id[2]) );
  GTECH_OR2 C71 ( .A(N37), .B(N38), .Z(N39) );
  GTECH_AND2 C72 ( .A(d8stg_fdiv_in), .B(div_id_out_in[2]), .Z(N37) );
  GTECH_AND2 C73 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[2]), .Z(N38) );
  GTECH_AND2 C74 ( .A(dest_rdy_in[0]), .B(add_id_out_in[2]), .Z(N40) );
  GTECH_OR2 C75 ( .A(N43), .B(N44), .Z(out_id[1]) );
  GTECH_OR2 C76 ( .A(N41), .B(N42), .Z(N43) );
  GTECH_AND2 C77 ( .A(d8stg_fdiv_in), .B(div_id_out_in[1]), .Z(N41) );
  GTECH_AND2 C78 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[1]), .Z(N42) );
  GTECH_AND2 C79 ( .A(dest_rdy_in[0]), .B(add_id_out_in[1]), .Z(N44) );
  GTECH_OR2 C80 ( .A(N47), .B(N48), .Z(out_id[0]) );
  GTECH_OR2 C81 ( .A(N45), .B(N46), .Z(N47) );
  GTECH_AND2 C82 ( .A(d8stg_fdiv_in), .B(div_id_out_in[0]), .Z(N45) );
  GTECH_AND2 C83 ( .A(dest_rdy_in[1]), .B(m6stg_id_in[0]), .Z(N46) );
  GTECH_AND2 C84 ( .A(dest_rdy_in[0]), .B(add_id_out_in[0]), .Z(N48) );
endmodule


module dff_SIZE77 ( din, clk, q, se, si, so );
  input [76:0] din;
  output [76:0] q;
  input [76:0] si;
  output [76:0] so;
  input clk, se;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79;
  assign so[76] = q[76];
  assign so[75] = q[75];
  assign so[74] = q[74];
  assign so[73] = q[73];
  assign so[72] = q[72];
  assign so[71] = q[71];
  assign so[70] = q[70];
  assign so[69] = q[69];
  assign so[68] = q[68];
  assign so[67] = q[67];
  assign so[66] = q[66];
  assign so[65] = q[65];
  assign so[64] = q[64];
  assign so[63] = q[63];
  assign so[62] = q[62];
  assign so[61] = q[61];
  assign so[60] = q[60];
  assign so[59] = q[59];
  assign so[58] = q[58];
  assign so[57] = q[57];
  assign so[56] = q[56];
  assign so[55] = q[55];
  assign so[54] = q[54];
  assign so[53] = q[53];
  assign so[52] = q[52];
  assign so[51] = q[51];
  assign so[50] = q[50];
  assign so[49] = q[49];
  assign so[48] = q[48];
  assign so[47] = q[47];
  assign so[46] = q[46];
  assign so[45] = q[45];
  assign so[44] = q[44];
  assign so[43] = q[43];
  assign so[42] = q[42];
  assign so[41] = q[41];
  assign so[40] = q[40];
  assign so[39] = q[39];
  assign so[38] = q[38];
  assign so[37] = q[37];
  assign so[36] = q[36];
  assign so[35] = q[35];
  assign so[34] = q[34];
  assign so[33] = q[33];
  assign so[32] = q[32];
  assign so[31] = q[31];
  assign so[30] = q[30];
  assign so[29] = q[29];
  assign so[28] = q[28];
  assign so[27] = q[27];
  assign so[26] = q[26];
  assign so[25] = q[25];
  assign so[24] = q[24];
  assign so[23] = q[23];
  assign so[22] = q[22];
  assign so[21] = q[21];
  assign so[20] = q[20];
  assign so[19] = q[19];
  assign so[18] = q[18];
  assign so[17] = q[17];
  assign so[16] = q[16];
  assign so[15] = q[15];
  assign so[14] = q[14];
  assign so[13] = q[13];
  assign so[12] = q[12];
  assign so[11] = q[11];
  assign so[10] = q[10];
  assign so[9] = q[9];
  assign so[8] = q[8];
  assign so[7] = q[7];
  assign so[6] = q[6];
  assign so[5] = q[5];
  assign so[4] = q[4];
  assign so[3] = q[3];
  assign so[2] = q[2];
  assign so[1] = q[1];
  assign so[0] = q[0];

  \**SEQGEN**  \q_reg[76]  ( .clear(1'b0), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[75]  ( .clear(1'b0), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[74]  ( .clear(1'b0), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[73]  ( .clear(1'b0), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[72]  ( .clear(1'b0), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[71]  ( .clear(1'b0), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[70]  ( .clear(1'b0), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[69]  ( .clear(1'b0), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[68]  ( .clear(1'b0), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[67]  ( .clear(1'b0), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[66]  ( .clear(1'b0), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[65]  ( .clear(1'b0), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[64]  ( .clear(1'b0), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[63]  ( .clear(1'b0), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[62]  ( .clear(1'b0), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[61]  ( .clear(1'b0), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[60]  ( .clear(1'b0), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[59]  ( .clear(1'b0), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[58]  ( .clear(1'b0), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[57]  ( .clear(1'b0), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[56]  ( .clear(1'b0), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[55]  ( .clear(1'b0), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[54]  ( .clear(1'b0), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[53]  ( .clear(1'b0), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[52]  ( .clear(1'b0), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[51]  ( .clear(1'b0), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[50]  ( .clear(1'b0), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[49]  ( .clear(1'b0), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[48]  ( .clear(1'b0), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[47]  ( .clear(1'b0), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[46]  ( .clear(1'b0), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[45]  ( .clear(1'b0), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[44]  ( .clear(1'b0), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[43]  ( .clear(1'b0), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[42]  ( .clear(1'b0), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[41]  ( .clear(1'b0), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[40]  ( .clear(1'b0), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[39]  ( .clear(1'b0), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[38]  ( .clear(1'b0), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[37]  ( .clear(1'b0), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[36]  ( .clear(1'b0), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[35]  ( .clear(1'b0), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[34]  ( .clear(1'b0), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[33]  ( .clear(1'b0), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[32]  ( .clear(1'b0), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(N14), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(N13), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(N12), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(N11), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(N10), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(N9), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(N8), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(N6), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(N5), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(N4), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \q_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(q[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C87 ( .DATA1(si), .DATA2(din), .CONTROL1(N0), .CONTROL2(N1), .Z({
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, 
        N9, N8, N7, N6, N5, N4, N3}) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module fpu_out_dp ( dest_rdy, req_thread, div_exc_out, d8stg_fdivd, 
        d8stg_fdivs, div_sign_out, div_exp_out, div_frac_out, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, add_exc_out, a6stg_fcmpop, add_cc_out, add_fcc_out, 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        add_sign_out, add_exp_out, add_frac_out, rclk, fp_cpx_data_ca, se, si, 
        so );
  input [2:0] dest_rdy;
  input [1:0] req_thread;
  input [4:0] div_exc_out;
  input [10:0] div_exp_out;
  input [51:0] div_frac_out;
  input [4:0] mul_exc_out;
  input [10:0] mul_exp_out;
  input [51:0] mul_frac_out;
  input [4:0] add_exc_out;
  input [1:0] add_cc_out;
  input [1:0] add_fcc_out;
  input [10:0] add_exp_out;
  input [63:0] add_frac_out;
  output [144:0] fp_cpx_data_ca;
  input d8stg_fdivd, d8stg_fdivs, div_sign_out, m6stg_fmul_dbl_dst,
         m6stg_fmuls, mul_sign_out, a6stg_fcmpop, a6stg_dbl_dst, a6stg_sng_dst,
         a6stg_long_dst, a6stg_int_dst, add_sign_out, rclk, se, si;
  output so;
  wire   fp_cpx_data_ca_144, fp_cpx_data_ca_143, fp_cpx_data_ca_142,
         fp_cpx_data_ca_141, fp_cpx_data_ca_140, fp_cpx_data_ca_136,
         fp_cpx_data_ca_135, fp_cpx_data_ca_134, se_l, clk,
         fp_cpx_data_ca_84_77_in_1, fp_cpx_data_ca_84_77_in_0,
         fp_cpx_data_ca_76_0_in_76, fp_cpx_data_ca_76_0_in_75,
         fp_cpx_data_ca_76_0_in_74, fp_cpx_data_ca_76_0_in_73,
         fp_cpx_data_ca_76_0_in_72, fp_cpx_data_ca_76_0_in_69,
         fp_cpx_data_ca_76_0_in_68, fp_cpx_data_ca_76_0_in_67,
         fp_cpx_data_ca_76_0_in_66, fp_cpx_data_ca_76_0_in_65, N0, N1, N2, N3,
         N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, net12208, net12209, net12210, net12211, net12212,
         net12213, net12214, net12215, net12216, net12217, net12218, net12219,
         net12220, net12221, net12222, net12223, net12224, net12225, net12226,
         net12227, net12228, net12229, net12230, net12231, net12232, net12233,
         net12234, net12235, net12236, net12237, net12238, net12239, net12240,
         net12241, net12242, net12243, net12244, net12245, net12246, net12247,
         net12248, net12249, net12250, net12251, net12252, net12253, net12254,
         net12255, net12256, net12257, net12258, net12259, net12260, net12261,
         net12262, net12263, net12264, net12265, net12266, net12267, net12268,
         net12269, net12270, net12271, net12272, net12273, net12274, net12275,
         net12276, net12277, net12278, net12279, net12280, net12281, net12282,
         net12283, net12284, net12285, net12286, net12287, net12288, net12289,
         net12290, net12291, net12292, net12293;
  wire   [63:0] add_out;
  wire   [63:0] mul_out;
  wire   [63:0] div_out;
  wire   [7:6] fp_cpx_data_ca_84_77_in;
  wire   [63:0] fp_cpx_data_ca_76_0_in;
  assign fp_cpx_data_ca[77] = 1'b0;
  assign fp_cpx_data_ca[78] = 1'b0;
  assign fp_cpx_data_ca[79] = 1'b0;
  assign fp_cpx_data_ca[80] = 1'b0;
  assign fp_cpx_data_ca[81] = 1'b0;
  assign fp_cpx_data_ca[82] = 1'b0;
  assign fp_cpx_data_ca[83] = 1'b0;
  assign fp_cpx_data_ca[84] = 1'b0;
  assign fp_cpx_data_ca[85] = 1'b0;
  assign fp_cpx_data_ca[86] = 1'b0;
  assign fp_cpx_data_ca[87] = 1'b0;
  assign fp_cpx_data_ca[88] = 1'b0;
  assign fp_cpx_data_ca[89] = 1'b0;
  assign fp_cpx_data_ca[90] = 1'b0;
  assign fp_cpx_data_ca[91] = 1'b0;
  assign fp_cpx_data_ca[92] = 1'b0;
  assign fp_cpx_data_ca[93] = 1'b0;
  assign fp_cpx_data_ca[94] = 1'b0;
  assign fp_cpx_data_ca[95] = 1'b0;
  assign fp_cpx_data_ca[96] = 1'b0;
  assign fp_cpx_data_ca[97] = 1'b0;
  assign fp_cpx_data_ca[98] = 1'b0;
  assign fp_cpx_data_ca[99] = 1'b0;
  assign fp_cpx_data_ca[100] = 1'b0;
  assign fp_cpx_data_ca[101] = 1'b0;
  assign fp_cpx_data_ca[102] = 1'b0;
  assign fp_cpx_data_ca[103] = 1'b0;
  assign fp_cpx_data_ca[104] = 1'b0;
  assign fp_cpx_data_ca[105] = 1'b0;
  assign fp_cpx_data_ca[106] = 1'b0;
  assign fp_cpx_data_ca[107] = 1'b0;
  assign fp_cpx_data_ca[108] = 1'b0;
  assign fp_cpx_data_ca[109] = 1'b0;
  assign fp_cpx_data_ca[110] = 1'b0;
  assign fp_cpx_data_ca[111] = 1'b0;
  assign fp_cpx_data_ca[112] = 1'b0;
  assign fp_cpx_data_ca[113] = 1'b0;
  assign fp_cpx_data_ca[114] = 1'b0;
  assign fp_cpx_data_ca[115] = 1'b0;
  assign fp_cpx_data_ca[116] = 1'b0;
  assign fp_cpx_data_ca[117] = 1'b0;
  assign fp_cpx_data_ca[118] = 1'b0;
  assign fp_cpx_data_ca[119] = 1'b0;
  assign fp_cpx_data_ca[120] = 1'b0;
  assign fp_cpx_data_ca[121] = 1'b0;
  assign fp_cpx_data_ca[122] = 1'b0;
  assign fp_cpx_data_ca[123] = 1'b0;
  assign fp_cpx_data_ca[124] = 1'b0;
  assign fp_cpx_data_ca[125] = 1'b0;
  assign fp_cpx_data_ca[126] = 1'b0;
  assign fp_cpx_data_ca[127] = 1'b0;
  assign fp_cpx_data_ca[128] = 1'b0;
  assign fp_cpx_data_ca[129] = 1'b0;
  assign fp_cpx_data_ca[130] = 1'b0;
  assign fp_cpx_data_ca[131] = 1'b0;
  assign fp_cpx_data_ca[132] = 1'b0;
  assign fp_cpx_data_ca[133] = 1'b0;
  assign fp_cpx_data_ca[137] = 1'b0;
  assign fp_cpx_data_ca[138] = 1'b0;
  assign fp_cpx_data_ca[139] = 1'b0;
  assign fp_cpx_data_ca[144] = fp_cpx_data_ca_144;
  assign fp_cpx_data_ca[143] = fp_cpx_data_ca_143;
  assign fp_cpx_data_ca[142] = fp_cpx_data_ca_142;
  assign fp_cpx_data_ca[141] = fp_cpx_data_ca_141;
  assign fp_cpx_data_ca[140] = fp_cpx_data_ca_140;
  assign fp_cpx_data_ca[136] = fp_cpx_data_ca_136;
  assign fp_cpx_data_ca[135] = fp_cpx_data_ca_135;
  assign fp_cpx_data_ca[134] = fp_cpx_data_ca_134;

  clken_buf ckbuf_out_dp ( .clk(clk), .rclk(rclk), .enb_l(1'b0), .tmb_l(se_l)
         );
  dff_SIZE8 i_fp_cpx_data_ca_84_77 ( .din({fp_cpx_data_ca_84_77_in, 1'b0, 1'b0, 
        1'b0, 1'b0, fp_cpx_data_ca_84_77_in_1, fp_cpx_data_ca_84_77_in_0}), 
        .clk(clk), .q({fp_cpx_data_ca_144, fp_cpx_data_ca_143, 
        fp_cpx_data_ca_142, fp_cpx_data_ca_141, fp_cpx_data_ca_140, 
        fp_cpx_data_ca_136, fp_cpx_data_ca_135, fp_cpx_data_ca_134}), .se(se), 
        .si({net12286, net12287, net12288, net12289, net12290, net12291, 
        net12292, net12293}) );
  dff_SIZE77 i_fp_cpx_data_ca_76_0 ( .din({fp_cpx_data_ca_76_0_in_76, 
        fp_cpx_data_ca_76_0_in_75, fp_cpx_data_ca_76_0_in_74, 
        fp_cpx_data_ca_76_0_in_73, fp_cpx_data_ca_76_0_in_72, 1'b0, 1'b0, 
        fp_cpx_data_ca_76_0_in_69, fp_cpx_data_ca_76_0_in_68, 
        fp_cpx_data_ca_76_0_in_67, fp_cpx_data_ca_76_0_in_66, 
        fp_cpx_data_ca_76_0_in_65, 1'b0, fp_cpx_data_ca_76_0_in}), .clk(clk), 
        .q(fp_cpx_data_ca[76:0]), .se(se), .si({net12209, net12210, net12211, 
        net12212, net12213, net12214, net12215, net12216, net12217, net12218, 
        net12219, net12220, net12221, net12222, net12223, net12224, net12225, 
        net12226, net12227, net12228, net12229, net12230, net12231, net12232, 
        net12233, net12234, net12235, net12236, net12237, net12238, net12239, 
        net12240, net12241, net12242, net12243, net12244, net12245, net12246, 
        net12247, net12248, net12249, net12250, net12251, net12252, net12253, 
        net12254, net12255, net12256, net12257, net12258, net12259, net12260, 
        net12261, net12262, net12263, net12264, net12265, net12266, net12267, 
        net12268, net12269, net12270, net12271, net12272, net12273, net12274, 
        net12275, net12276, net12277, net12278, net12279, net12280, net12281, 
        net12282, net12283, net12284, net12285}) );
  GTECH_NOT I_0 ( .A(se), .Z(se_l) );
  GTECH_OR2 C279 ( .A(N4), .B(N5), .Z(add_out[63]) );
  GTECH_OR2 C280 ( .A(N2), .B(N3), .Z(N4) );
  GTECH_OR2 C281 ( .A(N0), .B(N1), .Z(N2) );
  GTECH_AND2 C282 ( .A(a6stg_dbl_dst), .B(add_sign_out), .Z(N0) );
  GTECH_AND2 C283 ( .A(a6stg_sng_dst), .B(add_sign_out), .Z(N1) );
  GTECH_AND2 C284 ( .A(a6stg_long_dst), .B(add_frac_out[63]), .Z(N3) );
  GTECH_AND2 C285 ( .A(a6stg_int_dst), .B(add_frac_out[63]), .Z(N5) );
  GTECH_OR2 C286 ( .A(N10), .B(N11), .Z(add_out[62]) );
  GTECH_OR2 C287 ( .A(N8), .B(N9), .Z(N10) );
  GTECH_OR2 C288 ( .A(N6), .B(N7), .Z(N8) );
  GTECH_AND2 C289 ( .A(a6stg_dbl_dst), .B(add_exp_out[10]), .Z(N6) );
  GTECH_AND2 C290 ( .A(a6stg_sng_dst), .B(add_exp_out[7]), .Z(N7) );
  GTECH_AND2 C291 ( .A(a6stg_long_dst), .B(add_frac_out[62]), .Z(N9) );
  GTECH_AND2 C292 ( .A(a6stg_int_dst), .B(add_frac_out[62]), .Z(N11) );
  GTECH_OR2 C293 ( .A(N16), .B(N17), .Z(add_out[61]) );
  GTECH_OR2 C294 ( .A(N14), .B(N15), .Z(N16) );
  GTECH_OR2 C295 ( .A(N12), .B(N13), .Z(N14) );
  GTECH_AND2 C296 ( .A(a6stg_dbl_dst), .B(add_exp_out[9]), .Z(N12) );
  GTECH_AND2 C297 ( .A(a6stg_sng_dst), .B(add_exp_out[6]), .Z(N13) );
  GTECH_AND2 C298 ( .A(a6stg_long_dst), .B(add_frac_out[61]), .Z(N15) );
  GTECH_AND2 C299 ( .A(a6stg_int_dst), .B(add_frac_out[61]), .Z(N17) );
  GTECH_OR2 C300 ( .A(N22), .B(N23), .Z(add_out[60]) );
  GTECH_OR2 C301 ( .A(N20), .B(N21), .Z(N22) );
  GTECH_OR2 C302 ( .A(N18), .B(N19), .Z(N20) );
  GTECH_AND2 C303 ( .A(a6stg_dbl_dst), .B(add_exp_out[8]), .Z(N18) );
  GTECH_AND2 C304 ( .A(a6stg_sng_dst), .B(add_exp_out[5]), .Z(N19) );
  GTECH_AND2 C305 ( .A(a6stg_long_dst), .B(add_frac_out[60]), .Z(N21) );
  GTECH_AND2 C306 ( .A(a6stg_int_dst), .B(add_frac_out[60]), .Z(N23) );
  GTECH_OR2 C307 ( .A(N28), .B(N29), .Z(add_out[59]) );
  GTECH_OR2 C308 ( .A(N26), .B(N27), .Z(N28) );
  GTECH_OR2 C309 ( .A(N24), .B(N25), .Z(N26) );
  GTECH_AND2 C310 ( .A(a6stg_dbl_dst), .B(add_exp_out[7]), .Z(N24) );
  GTECH_AND2 C311 ( .A(a6stg_sng_dst), .B(add_exp_out[4]), .Z(N25) );
  GTECH_AND2 C312 ( .A(a6stg_long_dst), .B(add_frac_out[59]), .Z(N27) );
  GTECH_AND2 C313 ( .A(a6stg_int_dst), .B(add_frac_out[59]), .Z(N29) );
  GTECH_OR2 C314 ( .A(N34), .B(N35), .Z(add_out[58]) );
  GTECH_OR2 C315 ( .A(N32), .B(N33), .Z(N34) );
  GTECH_OR2 C316 ( .A(N30), .B(N31), .Z(N32) );
  GTECH_AND2 C317 ( .A(a6stg_dbl_dst), .B(add_exp_out[6]), .Z(N30) );
  GTECH_AND2 C318 ( .A(a6stg_sng_dst), .B(add_exp_out[3]), .Z(N31) );
  GTECH_AND2 C319 ( .A(a6stg_long_dst), .B(add_frac_out[58]), .Z(N33) );
  GTECH_AND2 C320 ( .A(a6stg_int_dst), .B(add_frac_out[58]), .Z(N35) );
  GTECH_OR2 C321 ( .A(N40), .B(N41), .Z(add_out[57]) );
  GTECH_OR2 C322 ( .A(N38), .B(N39), .Z(N40) );
  GTECH_OR2 C323 ( .A(N36), .B(N37), .Z(N38) );
  GTECH_AND2 C324 ( .A(a6stg_dbl_dst), .B(add_exp_out[5]), .Z(N36) );
  GTECH_AND2 C325 ( .A(a6stg_sng_dst), .B(add_exp_out[2]), .Z(N37) );
  GTECH_AND2 C326 ( .A(a6stg_long_dst), .B(add_frac_out[57]), .Z(N39) );
  GTECH_AND2 C327 ( .A(a6stg_int_dst), .B(add_frac_out[57]), .Z(N41) );
  GTECH_OR2 C328 ( .A(N46), .B(N47), .Z(add_out[56]) );
  GTECH_OR2 C329 ( .A(N44), .B(N45), .Z(N46) );
  GTECH_OR2 C330 ( .A(N42), .B(N43), .Z(N44) );
  GTECH_AND2 C331 ( .A(a6stg_dbl_dst), .B(add_exp_out[4]), .Z(N42) );
  GTECH_AND2 C332 ( .A(a6stg_sng_dst), .B(add_exp_out[1]), .Z(N43) );
  GTECH_AND2 C333 ( .A(a6stg_long_dst), .B(add_frac_out[56]), .Z(N45) );
  GTECH_AND2 C334 ( .A(a6stg_int_dst), .B(add_frac_out[56]), .Z(N47) );
  GTECH_OR2 C335 ( .A(N52), .B(N53), .Z(add_out[55]) );
  GTECH_OR2 C336 ( .A(N50), .B(N51), .Z(N52) );
  GTECH_OR2 C337 ( .A(N48), .B(N49), .Z(N50) );
  GTECH_AND2 C338 ( .A(a6stg_dbl_dst), .B(add_exp_out[3]), .Z(N48) );
  GTECH_AND2 C339 ( .A(a6stg_sng_dst), .B(add_exp_out[0]), .Z(N49) );
  GTECH_AND2 C340 ( .A(a6stg_long_dst), .B(add_frac_out[55]), .Z(N51) );
  GTECH_AND2 C341 ( .A(a6stg_int_dst), .B(add_frac_out[55]), .Z(N53) );
  GTECH_OR2 C342 ( .A(N58), .B(N59), .Z(add_out[54]) );
  GTECH_OR2 C343 ( .A(N56), .B(N57), .Z(N58) );
  GTECH_OR2 C344 ( .A(N54), .B(N55), .Z(N56) );
  GTECH_AND2 C345 ( .A(a6stg_dbl_dst), .B(add_exp_out[2]), .Z(N54) );
  GTECH_AND2 C346 ( .A(a6stg_sng_dst), .B(add_frac_out[62]), .Z(N55) );
  GTECH_AND2 C347 ( .A(a6stg_long_dst), .B(add_frac_out[54]), .Z(N57) );
  GTECH_AND2 C348 ( .A(a6stg_int_dst), .B(add_frac_out[54]), .Z(N59) );
  GTECH_OR2 C349 ( .A(N64), .B(N65), .Z(add_out[53]) );
  GTECH_OR2 C350 ( .A(N62), .B(N63), .Z(N64) );
  GTECH_OR2 C351 ( .A(N60), .B(N61), .Z(N62) );
  GTECH_AND2 C352 ( .A(a6stg_dbl_dst), .B(add_exp_out[1]), .Z(N60) );
  GTECH_AND2 C353 ( .A(a6stg_sng_dst), .B(add_frac_out[61]), .Z(N61) );
  GTECH_AND2 C354 ( .A(a6stg_long_dst), .B(add_frac_out[53]), .Z(N63) );
  GTECH_AND2 C355 ( .A(a6stg_int_dst), .B(add_frac_out[53]), .Z(N65) );
  GTECH_OR2 C356 ( .A(N70), .B(N71), .Z(add_out[52]) );
  GTECH_OR2 C357 ( .A(N68), .B(N69), .Z(N70) );
  GTECH_OR2 C358 ( .A(N66), .B(N67), .Z(N68) );
  GTECH_AND2 C359 ( .A(a6stg_dbl_dst), .B(add_exp_out[0]), .Z(N66) );
  GTECH_AND2 C360 ( .A(a6stg_sng_dst), .B(add_frac_out[60]), .Z(N67) );
  GTECH_AND2 C361 ( .A(a6stg_long_dst), .B(add_frac_out[52]), .Z(N69) );
  GTECH_AND2 C362 ( .A(a6stg_int_dst), .B(add_frac_out[52]), .Z(N71) );
  GTECH_OR2 C363 ( .A(N76), .B(N77), .Z(add_out[51]) );
  GTECH_OR2 C364 ( .A(N74), .B(N75), .Z(N76) );
  GTECH_OR2 C365 ( .A(N72), .B(N73), .Z(N74) );
  GTECH_AND2 C366 ( .A(a6stg_dbl_dst), .B(add_frac_out[62]), .Z(N72) );
  GTECH_AND2 C367 ( .A(a6stg_sng_dst), .B(add_frac_out[59]), .Z(N73) );
  GTECH_AND2 C368 ( .A(a6stg_long_dst), .B(add_frac_out[51]), .Z(N75) );
  GTECH_AND2 C369 ( .A(a6stg_int_dst), .B(add_frac_out[51]), .Z(N77) );
  GTECH_OR2 C370 ( .A(N82), .B(N83), .Z(add_out[50]) );
  GTECH_OR2 C371 ( .A(N80), .B(N81), .Z(N82) );
  GTECH_OR2 C372 ( .A(N78), .B(N79), .Z(N80) );
  GTECH_AND2 C373 ( .A(a6stg_dbl_dst), .B(add_frac_out[61]), .Z(N78) );
  GTECH_AND2 C374 ( .A(a6stg_sng_dst), .B(add_frac_out[58]), .Z(N79) );
  GTECH_AND2 C375 ( .A(a6stg_long_dst), .B(add_frac_out[50]), .Z(N81) );
  GTECH_AND2 C376 ( .A(a6stg_int_dst), .B(add_frac_out[50]), .Z(N83) );
  GTECH_OR2 C377 ( .A(N88), .B(N89), .Z(add_out[49]) );
  GTECH_OR2 C378 ( .A(N86), .B(N87), .Z(N88) );
  GTECH_OR2 C379 ( .A(N84), .B(N85), .Z(N86) );
  GTECH_AND2 C380 ( .A(a6stg_dbl_dst), .B(add_frac_out[60]), .Z(N84) );
  GTECH_AND2 C381 ( .A(a6stg_sng_dst), .B(add_frac_out[57]), .Z(N85) );
  GTECH_AND2 C382 ( .A(a6stg_long_dst), .B(add_frac_out[49]), .Z(N87) );
  GTECH_AND2 C383 ( .A(a6stg_int_dst), .B(add_frac_out[49]), .Z(N89) );
  GTECH_OR2 C384 ( .A(N94), .B(N95), .Z(add_out[48]) );
  GTECH_OR2 C385 ( .A(N92), .B(N93), .Z(N94) );
  GTECH_OR2 C386 ( .A(N90), .B(N91), .Z(N92) );
  GTECH_AND2 C387 ( .A(a6stg_dbl_dst), .B(add_frac_out[59]), .Z(N90) );
  GTECH_AND2 C388 ( .A(a6stg_sng_dst), .B(add_frac_out[56]), .Z(N91) );
  GTECH_AND2 C389 ( .A(a6stg_long_dst), .B(add_frac_out[48]), .Z(N93) );
  GTECH_AND2 C390 ( .A(a6stg_int_dst), .B(add_frac_out[48]), .Z(N95) );
  GTECH_OR2 C391 ( .A(N100), .B(N101), .Z(add_out[47]) );
  GTECH_OR2 C392 ( .A(N98), .B(N99), .Z(N100) );
  GTECH_OR2 C393 ( .A(N96), .B(N97), .Z(N98) );
  GTECH_AND2 C394 ( .A(a6stg_dbl_dst), .B(add_frac_out[58]), .Z(N96) );
  GTECH_AND2 C395 ( .A(a6stg_sng_dst), .B(add_frac_out[55]), .Z(N97) );
  GTECH_AND2 C396 ( .A(a6stg_long_dst), .B(add_frac_out[47]), .Z(N99) );
  GTECH_AND2 C397 ( .A(a6stg_int_dst), .B(add_frac_out[47]), .Z(N101) );
  GTECH_OR2 C398 ( .A(N106), .B(N107), .Z(add_out[46]) );
  GTECH_OR2 C399 ( .A(N104), .B(N105), .Z(N106) );
  GTECH_OR2 C400 ( .A(N102), .B(N103), .Z(N104) );
  GTECH_AND2 C401 ( .A(a6stg_dbl_dst), .B(add_frac_out[57]), .Z(N102) );
  GTECH_AND2 C402 ( .A(a6stg_sng_dst), .B(add_frac_out[54]), .Z(N103) );
  GTECH_AND2 C403 ( .A(a6stg_long_dst), .B(add_frac_out[46]), .Z(N105) );
  GTECH_AND2 C404 ( .A(a6stg_int_dst), .B(add_frac_out[46]), .Z(N107) );
  GTECH_OR2 C405 ( .A(N112), .B(N113), .Z(add_out[45]) );
  GTECH_OR2 C406 ( .A(N110), .B(N111), .Z(N112) );
  GTECH_OR2 C407 ( .A(N108), .B(N109), .Z(N110) );
  GTECH_AND2 C408 ( .A(a6stg_dbl_dst), .B(add_frac_out[56]), .Z(N108) );
  GTECH_AND2 C409 ( .A(a6stg_sng_dst), .B(add_frac_out[53]), .Z(N109) );
  GTECH_AND2 C410 ( .A(a6stg_long_dst), .B(add_frac_out[45]), .Z(N111) );
  GTECH_AND2 C411 ( .A(a6stg_int_dst), .B(add_frac_out[45]), .Z(N113) );
  GTECH_OR2 C412 ( .A(N118), .B(N119), .Z(add_out[44]) );
  GTECH_OR2 C413 ( .A(N116), .B(N117), .Z(N118) );
  GTECH_OR2 C414 ( .A(N114), .B(N115), .Z(N116) );
  GTECH_AND2 C415 ( .A(a6stg_dbl_dst), .B(add_frac_out[55]), .Z(N114) );
  GTECH_AND2 C416 ( .A(a6stg_sng_dst), .B(add_frac_out[52]), .Z(N115) );
  GTECH_AND2 C417 ( .A(a6stg_long_dst), .B(add_frac_out[44]), .Z(N117) );
  GTECH_AND2 C418 ( .A(a6stg_int_dst), .B(add_frac_out[44]), .Z(N119) );
  GTECH_OR2 C419 ( .A(N124), .B(N125), .Z(add_out[43]) );
  GTECH_OR2 C420 ( .A(N122), .B(N123), .Z(N124) );
  GTECH_OR2 C421 ( .A(N120), .B(N121), .Z(N122) );
  GTECH_AND2 C422 ( .A(a6stg_dbl_dst), .B(add_frac_out[54]), .Z(N120) );
  GTECH_AND2 C423 ( .A(a6stg_sng_dst), .B(add_frac_out[51]), .Z(N121) );
  GTECH_AND2 C424 ( .A(a6stg_long_dst), .B(add_frac_out[43]), .Z(N123) );
  GTECH_AND2 C425 ( .A(a6stg_int_dst), .B(add_frac_out[43]), .Z(N125) );
  GTECH_OR2 C426 ( .A(N130), .B(N131), .Z(add_out[42]) );
  GTECH_OR2 C427 ( .A(N128), .B(N129), .Z(N130) );
  GTECH_OR2 C428 ( .A(N126), .B(N127), .Z(N128) );
  GTECH_AND2 C429 ( .A(a6stg_dbl_dst), .B(add_frac_out[53]), .Z(N126) );
  GTECH_AND2 C430 ( .A(a6stg_sng_dst), .B(add_frac_out[50]), .Z(N127) );
  GTECH_AND2 C431 ( .A(a6stg_long_dst), .B(add_frac_out[42]), .Z(N129) );
  GTECH_AND2 C432 ( .A(a6stg_int_dst), .B(add_frac_out[42]), .Z(N131) );
  GTECH_OR2 C433 ( .A(N136), .B(N137), .Z(add_out[41]) );
  GTECH_OR2 C434 ( .A(N134), .B(N135), .Z(N136) );
  GTECH_OR2 C435 ( .A(N132), .B(N133), .Z(N134) );
  GTECH_AND2 C436 ( .A(a6stg_dbl_dst), .B(add_frac_out[52]), .Z(N132) );
  GTECH_AND2 C437 ( .A(a6stg_sng_dst), .B(add_frac_out[49]), .Z(N133) );
  GTECH_AND2 C438 ( .A(a6stg_long_dst), .B(add_frac_out[41]), .Z(N135) );
  GTECH_AND2 C439 ( .A(a6stg_int_dst), .B(add_frac_out[41]), .Z(N137) );
  GTECH_OR2 C440 ( .A(N142), .B(N143), .Z(add_out[40]) );
  GTECH_OR2 C441 ( .A(N140), .B(N141), .Z(N142) );
  GTECH_OR2 C442 ( .A(N138), .B(N139), .Z(N140) );
  GTECH_AND2 C443 ( .A(a6stg_dbl_dst), .B(add_frac_out[51]), .Z(N138) );
  GTECH_AND2 C444 ( .A(a6stg_sng_dst), .B(add_frac_out[48]), .Z(N139) );
  GTECH_AND2 C445 ( .A(a6stg_long_dst), .B(add_frac_out[40]), .Z(N141) );
  GTECH_AND2 C446 ( .A(a6stg_int_dst), .B(add_frac_out[40]), .Z(N143) );
  GTECH_OR2 C447 ( .A(N148), .B(N149), .Z(add_out[39]) );
  GTECH_OR2 C448 ( .A(N146), .B(N147), .Z(N148) );
  GTECH_OR2 C449 ( .A(N144), .B(N145), .Z(N146) );
  GTECH_AND2 C450 ( .A(a6stg_dbl_dst), .B(add_frac_out[50]), .Z(N144) );
  GTECH_AND2 C451 ( .A(a6stg_sng_dst), .B(add_frac_out[47]), .Z(N145) );
  GTECH_AND2 C452 ( .A(a6stg_long_dst), .B(add_frac_out[39]), .Z(N147) );
  GTECH_AND2 C453 ( .A(a6stg_int_dst), .B(add_frac_out[39]), .Z(N149) );
  GTECH_OR2 C454 ( .A(N154), .B(N155), .Z(add_out[38]) );
  GTECH_OR2 C455 ( .A(N152), .B(N153), .Z(N154) );
  GTECH_OR2 C456 ( .A(N150), .B(N151), .Z(N152) );
  GTECH_AND2 C457 ( .A(a6stg_dbl_dst), .B(add_frac_out[49]), .Z(N150) );
  GTECH_AND2 C458 ( .A(a6stg_sng_dst), .B(add_frac_out[46]), .Z(N151) );
  GTECH_AND2 C459 ( .A(a6stg_long_dst), .B(add_frac_out[38]), .Z(N153) );
  GTECH_AND2 C460 ( .A(a6stg_int_dst), .B(add_frac_out[38]), .Z(N155) );
  GTECH_OR2 C461 ( .A(N160), .B(N161), .Z(add_out[37]) );
  GTECH_OR2 C462 ( .A(N158), .B(N159), .Z(N160) );
  GTECH_OR2 C463 ( .A(N156), .B(N157), .Z(N158) );
  GTECH_AND2 C464 ( .A(a6stg_dbl_dst), .B(add_frac_out[48]), .Z(N156) );
  GTECH_AND2 C465 ( .A(a6stg_sng_dst), .B(add_frac_out[45]), .Z(N157) );
  GTECH_AND2 C466 ( .A(a6stg_long_dst), .B(add_frac_out[37]), .Z(N159) );
  GTECH_AND2 C467 ( .A(a6stg_int_dst), .B(add_frac_out[37]), .Z(N161) );
  GTECH_OR2 C468 ( .A(N166), .B(N167), .Z(add_out[36]) );
  GTECH_OR2 C469 ( .A(N164), .B(N165), .Z(N166) );
  GTECH_OR2 C470 ( .A(N162), .B(N163), .Z(N164) );
  GTECH_AND2 C471 ( .A(a6stg_dbl_dst), .B(add_frac_out[47]), .Z(N162) );
  GTECH_AND2 C472 ( .A(a6stg_sng_dst), .B(add_frac_out[44]), .Z(N163) );
  GTECH_AND2 C473 ( .A(a6stg_long_dst), .B(add_frac_out[36]), .Z(N165) );
  GTECH_AND2 C474 ( .A(a6stg_int_dst), .B(add_frac_out[36]), .Z(N167) );
  GTECH_OR2 C475 ( .A(N172), .B(N173), .Z(add_out[35]) );
  GTECH_OR2 C476 ( .A(N170), .B(N171), .Z(N172) );
  GTECH_OR2 C477 ( .A(N168), .B(N169), .Z(N170) );
  GTECH_AND2 C478 ( .A(a6stg_dbl_dst), .B(add_frac_out[46]), .Z(N168) );
  GTECH_AND2 C479 ( .A(a6stg_sng_dst), .B(add_frac_out[43]), .Z(N169) );
  GTECH_AND2 C480 ( .A(a6stg_long_dst), .B(add_frac_out[35]), .Z(N171) );
  GTECH_AND2 C481 ( .A(a6stg_int_dst), .B(add_frac_out[35]), .Z(N173) );
  GTECH_OR2 C482 ( .A(N178), .B(N179), .Z(add_out[34]) );
  GTECH_OR2 C483 ( .A(N176), .B(N177), .Z(N178) );
  GTECH_OR2 C484 ( .A(N174), .B(N175), .Z(N176) );
  GTECH_AND2 C485 ( .A(a6stg_dbl_dst), .B(add_frac_out[45]), .Z(N174) );
  GTECH_AND2 C486 ( .A(a6stg_sng_dst), .B(add_frac_out[42]), .Z(N175) );
  GTECH_AND2 C487 ( .A(a6stg_long_dst), .B(add_frac_out[34]), .Z(N177) );
  GTECH_AND2 C488 ( .A(a6stg_int_dst), .B(add_frac_out[34]), .Z(N179) );
  GTECH_OR2 C489 ( .A(N184), .B(N185), .Z(add_out[33]) );
  GTECH_OR2 C490 ( .A(N182), .B(N183), .Z(N184) );
  GTECH_OR2 C491 ( .A(N180), .B(N181), .Z(N182) );
  GTECH_AND2 C492 ( .A(a6stg_dbl_dst), .B(add_frac_out[44]), .Z(N180) );
  GTECH_AND2 C493 ( .A(a6stg_sng_dst), .B(add_frac_out[41]), .Z(N181) );
  GTECH_AND2 C494 ( .A(a6stg_long_dst), .B(add_frac_out[33]), .Z(N183) );
  GTECH_AND2 C495 ( .A(a6stg_int_dst), .B(add_frac_out[33]), .Z(N185) );
  GTECH_OR2 C496 ( .A(N190), .B(N191), .Z(add_out[32]) );
  GTECH_OR2 C497 ( .A(N188), .B(N189), .Z(N190) );
  GTECH_OR2 C498 ( .A(N186), .B(N187), .Z(N188) );
  GTECH_AND2 C499 ( .A(a6stg_dbl_dst), .B(add_frac_out[43]), .Z(N186) );
  GTECH_AND2 C500 ( .A(a6stg_sng_dst), .B(add_frac_out[40]), .Z(N187) );
  GTECH_AND2 C501 ( .A(a6stg_long_dst), .B(add_frac_out[32]), .Z(N189) );
  GTECH_AND2 C502 ( .A(a6stg_int_dst), .B(add_frac_out[32]), .Z(N191) );
  GTECH_OR2 C503 ( .A(N192), .B(N193), .Z(add_out[31]) );
  GTECH_AND2 C504 ( .A(a6stg_dbl_dst), .B(add_frac_out[42]), .Z(N192) );
  GTECH_AND2 C505 ( .A(a6stg_long_dst), .B(add_frac_out[31]), .Z(N193) );
  GTECH_OR2 C506 ( .A(N194), .B(N195), .Z(add_out[30]) );
  GTECH_AND2 C507 ( .A(a6stg_dbl_dst), .B(add_frac_out[41]), .Z(N194) );
  GTECH_AND2 C508 ( .A(a6stg_long_dst), .B(add_frac_out[30]), .Z(N195) );
  GTECH_OR2 C509 ( .A(N196), .B(N197), .Z(add_out[29]) );
  GTECH_AND2 C510 ( .A(a6stg_dbl_dst), .B(add_frac_out[40]), .Z(N196) );
  GTECH_AND2 C511 ( .A(a6stg_long_dst), .B(add_frac_out[29]), .Z(N197) );
  GTECH_OR2 C512 ( .A(N198), .B(N199), .Z(add_out[28]) );
  GTECH_AND2 C513 ( .A(a6stg_dbl_dst), .B(add_frac_out[39]), .Z(N198) );
  GTECH_AND2 C514 ( .A(a6stg_long_dst), .B(add_frac_out[28]), .Z(N199) );
  GTECH_OR2 C515 ( .A(N200), .B(N201), .Z(add_out[27]) );
  GTECH_AND2 C516 ( .A(a6stg_dbl_dst), .B(add_frac_out[38]), .Z(N200) );
  GTECH_AND2 C517 ( .A(a6stg_long_dst), .B(add_frac_out[27]), .Z(N201) );
  GTECH_OR2 C518 ( .A(N202), .B(N203), .Z(add_out[26]) );
  GTECH_AND2 C519 ( .A(a6stg_dbl_dst), .B(add_frac_out[37]), .Z(N202) );
  GTECH_AND2 C520 ( .A(a6stg_long_dst), .B(add_frac_out[26]), .Z(N203) );
  GTECH_OR2 C521 ( .A(N204), .B(N205), .Z(add_out[25]) );
  GTECH_AND2 C522 ( .A(a6stg_dbl_dst), .B(add_frac_out[36]), .Z(N204) );
  GTECH_AND2 C523 ( .A(a6stg_long_dst), .B(add_frac_out[25]), .Z(N205) );
  GTECH_OR2 C524 ( .A(N206), .B(N207), .Z(add_out[24]) );
  GTECH_AND2 C525 ( .A(a6stg_dbl_dst), .B(add_frac_out[35]), .Z(N206) );
  GTECH_AND2 C526 ( .A(a6stg_long_dst), .B(add_frac_out[24]), .Z(N207) );
  GTECH_OR2 C527 ( .A(N208), .B(N209), .Z(add_out[23]) );
  GTECH_AND2 C528 ( .A(a6stg_dbl_dst), .B(add_frac_out[34]), .Z(N208) );
  GTECH_AND2 C529 ( .A(a6stg_long_dst), .B(add_frac_out[23]), .Z(N209) );
  GTECH_OR2 C530 ( .A(N210), .B(N211), .Z(add_out[22]) );
  GTECH_AND2 C531 ( .A(a6stg_dbl_dst), .B(add_frac_out[33]), .Z(N210) );
  GTECH_AND2 C532 ( .A(a6stg_long_dst), .B(add_frac_out[22]), .Z(N211) );
  GTECH_OR2 C533 ( .A(N212), .B(N213), .Z(add_out[21]) );
  GTECH_AND2 C534 ( .A(a6stg_dbl_dst), .B(add_frac_out[32]), .Z(N212) );
  GTECH_AND2 C535 ( .A(a6stg_long_dst), .B(add_frac_out[21]), .Z(N213) );
  GTECH_OR2 C536 ( .A(N214), .B(N215), .Z(add_out[20]) );
  GTECH_AND2 C537 ( .A(a6stg_dbl_dst), .B(add_frac_out[31]), .Z(N214) );
  GTECH_AND2 C538 ( .A(a6stg_long_dst), .B(add_frac_out[20]), .Z(N215) );
  GTECH_OR2 C539 ( .A(N216), .B(N217), .Z(add_out[19]) );
  GTECH_AND2 C540 ( .A(a6stg_dbl_dst), .B(add_frac_out[30]), .Z(N216) );
  GTECH_AND2 C541 ( .A(a6stg_long_dst), .B(add_frac_out[19]), .Z(N217) );
  GTECH_OR2 C542 ( .A(N218), .B(N219), .Z(add_out[18]) );
  GTECH_AND2 C543 ( .A(a6stg_dbl_dst), .B(add_frac_out[29]), .Z(N218) );
  GTECH_AND2 C544 ( .A(a6stg_long_dst), .B(add_frac_out[18]), .Z(N219) );
  GTECH_OR2 C545 ( .A(N220), .B(N221), .Z(add_out[17]) );
  GTECH_AND2 C546 ( .A(a6stg_dbl_dst), .B(add_frac_out[28]), .Z(N220) );
  GTECH_AND2 C547 ( .A(a6stg_long_dst), .B(add_frac_out[17]), .Z(N221) );
  GTECH_OR2 C548 ( .A(N222), .B(N223), .Z(add_out[16]) );
  GTECH_AND2 C549 ( .A(a6stg_dbl_dst), .B(add_frac_out[27]), .Z(N222) );
  GTECH_AND2 C550 ( .A(a6stg_long_dst), .B(add_frac_out[16]), .Z(N223) );
  GTECH_OR2 C551 ( .A(N224), .B(N225), .Z(add_out[15]) );
  GTECH_AND2 C552 ( .A(a6stg_dbl_dst), .B(add_frac_out[26]), .Z(N224) );
  GTECH_AND2 C553 ( .A(a6stg_long_dst), .B(add_frac_out[15]), .Z(N225) );
  GTECH_OR2 C554 ( .A(N226), .B(N227), .Z(add_out[14]) );
  GTECH_AND2 C555 ( .A(a6stg_dbl_dst), .B(add_frac_out[25]), .Z(N226) );
  GTECH_AND2 C556 ( .A(a6stg_long_dst), .B(add_frac_out[14]), .Z(N227) );
  GTECH_OR2 C557 ( .A(N228), .B(N229), .Z(add_out[13]) );
  GTECH_AND2 C558 ( .A(a6stg_dbl_dst), .B(add_frac_out[24]), .Z(N228) );
  GTECH_AND2 C559 ( .A(a6stg_long_dst), .B(add_frac_out[13]), .Z(N229) );
  GTECH_OR2 C560 ( .A(N230), .B(N231), .Z(add_out[12]) );
  GTECH_AND2 C561 ( .A(a6stg_dbl_dst), .B(add_frac_out[23]), .Z(N230) );
  GTECH_AND2 C562 ( .A(a6stg_long_dst), .B(add_frac_out[12]), .Z(N231) );
  GTECH_OR2 C563 ( .A(N232), .B(N233), .Z(add_out[11]) );
  GTECH_AND2 C564 ( .A(a6stg_dbl_dst), .B(add_frac_out[22]), .Z(N232) );
  GTECH_AND2 C565 ( .A(a6stg_long_dst), .B(add_frac_out[11]), .Z(N233) );
  GTECH_OR2 C566 ( .A(N234), .B(N235), .Z(add_out[10]) );
  GTECH_AND2 C567 ( .A(a6stg_dbl_dst), .B(add_frac_out[21]), .Z(N234) );
  GTECH_AND2 C568 ( .A(a6stg_long_dst), .B(add_frac_out[10]), .Z(N235) );
  GTECH_OR2 C569 ( .A(N236), .B(N237), .Z(add_out[9]) );
  GTECH_AND2 C570 ( .A(a6stg_dbl_dst), .B(add_frac_out[20]), .Z(N236) );
  GTECH_AND2 C571 ( .A(a6stg_long_dst), .B(add_frac_out[9]), .Z(N237) );
  GTECH_OR2 C572 ( .A(N238), .B(N239), .Z(add_out[8]) );
  GTECH_AND2 C573 ( .A(a6stg_dbl_dst), .B(add_frac_out[19]), .Z(N238) );
  GTECH_AND2 C574 ( .A(a6stg_long_dst), .B(add_frac_out[8]), .Z(N239) );
  GTECH_OR2 C575 ( .A(N240), .B(N241), .Z(add_out[7]) );
  GTECH_AND2 C576 ( .A(a6stg_dbl_dst), .B(add_frac_out[18]), .Z(N240) );
  GTECH_AND2 C577 ( .A(a6stg_long_dst), .B(add_frac_out[7]), .Z(N241) );
  GTECH_OR2 C578 ( .A(N242), .B(N243), .Z(add_out[6]) );
  GTECH_AND2 C579 ( .A(a6stg_dbl_dst), .B(add_frac_out[17]), .Z(N242) );
  GTECH_AND2 C580 ( .A(a6stg_long_dst), .B(add_frac_out[6]), .Z(N243) );
  GTECH_OR2 C581 ( .A(N244), .B(N245), .Z(add_out[5]) );
  GTECH_AND2 C582 ( .A(a6stg_dbl_dst), .B(add_frac_out[16]), .Z(N244) );
  GTECH_AND2 C583 ( .A(a6stg_long_dst), .B(add_frac_out[5]), .Z(N245) );
  GTECH_OR2 C584 ( .A(N246), .B(N247), .Z(add_out[4]) );
  GTECH_AND2 C585 ( .A(a6stg_dbl_dst), .B(add_frac_out[15]), .Z(N246) );
  GTECH_AND2 C586 ( .A(a6stg_long_dst), .B(add_frac_out[4]), .Z(N247) );
  GTECH_OR2 C587 ( .A(N248), .B(N249), .Z(add_out[3]) );
  GTECH_AND2 C588 ( .A(a6stg_dbl_dst), .B(add_frac_out[14]), .Z(N248) );
  GTECH_AND2 C589 ( .A(a6stg_long_dst), .B(add_frac_out[3]), .Z(N249) );
  GTECH_OR2 C590 ( .A(N250), .B(N251), .Z(add_out[2]) );
  GTECH_AND2 C591 ( .A(a6stg_dbl_dst), .B(add_frac_out[13]), .Z(N250) );
  GTECH_AND2 C592 ( .A(a6stg_long_dst), .B(add_frac_out[2]), .Z(N251) );
  GTECH_OR2 C593 ( .A(N252), .B(N253), .Z(add_out[1]) );
  GTECH_AND2 C594 ( .A(a6stg_dbl_dst), .B(add_frac_out[12]), .Z(N252) );
  GTECH_AND2 C595 ( .A(a6stg_long_dst), .B(add_frac_out[1]), .Z(N253) );
  GTECH_OR2 C596 ( .A(N254), .B(N255), .Z(add_out[0]) );
  GTECH_AND2 C597 ( .A(a6stg_dbl_dst), .B(add_frac_out[11]), .Z(N254) );
  GTECH_AND2 C598 ( .A(a6stg_long_dst), .B(add_frac_out[0]), .Z(N255) );
  GTECH_OR2 C599 ( .A(N256), .B(N257), .Z(mul_out[63]) );
  GTECH_AND2 C600 ( .A(m6stg_fmul_dbl_dst), .B(mul_sign_out), .Z(N256) );
  GTECH_AND2 C601 ( .A(m6stg_fmuls), .B(mul_sign_out), .Z(N257) );
  GTECH_OR2 C602 ( .A(N258), .B(N259), .Z(mul_out[62]) );
  GTECH_AND2 C603 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[10]), .Z(N258) );
  GTECH_AND2 C604 ( .A(m6stg_fmuls), .B(mul_exp_out[7]), .Z(N259) );
  GTECH_OR2 C605 ( .A(N260), .B(N261), .Z(mul_out[61]) );
  GTECH_AND2 C606 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[9]), .Z(N260) );
  GTECH_AND2 C607 ( .A(m6stg_fmuls), .B(mul_exp_out[6]), .Z(N261) );
  GTECH_OR2 C608 ( .A(N262), .B(N263), .Z(mul_out[60]) );
  GTECH_AND2 C609 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[8]), .Z(N262) );
  GTECH_AND2 C610 ( .A(m6stg_fmuls), .B(mul_exp_out[5]), .Z(N263) );
  GTECH_OR2 C611 ( .A(N264), .B(N265), .Z(mul_out[59]) );
  GTECH_AND2 C612 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[7]), .Z(N264) );
  GTECH_AND2 C613 ( .A(m6stg_fmuls), .B(mul_exp_out[4]), .Z(N265) );
  GTECH_OR2 C614 ( .A(N266), .B(N267), .Z(mul_out[58]) );
  GTECH_AND2 C615 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[6]), .Z(N266) );
  GTECH_AND2 C616 ( .A(m6stg_fmuls), .B(mul_exp_out[3]), .Z(N267) );
  GTECH_OR2 C617 ( .A(N268), .B(N269), .Z(mul_out[57]) );
  GTECH_AND2 C618 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[5]), .Z(N268) );
  GTECH_AND2 C619 ( .A(m6stg_fmuls), .B(mul_exp_out[2]), .Z(N269) );
  GTECH_OR2 C620 ( .A(N270), .B(N271), .Z(mul_out[56]) );
  GTECH_AND2 C621 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[4]), .Z(N270) );
  GTECH_AND2 C622 ( .A(m6stg_fmuls), .B(mul_exp_out[1]), .Z(N271) );
  GTECH_OR2 C623 ( .A(N272), .B(N273), .Z(mul_out[55]) );
  GTECH_AND2 C624 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[3]), .Z(N272) );
  GTECH_AND2 C625 ( .A(m6stg_fmuls), .B(mul_exp_out[0]), .Z(N273) );
  GTECH_OR2 C626 ( .A(N274), .B(N275), .Z(mul_out[54]) );
  GTECH_AND2 C627 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[2]), .Z(N274) );
  GTECH_AND2 C628 ( .A(m6stg_fmuls), .B(mul_frac_out[51]), .Z(N275) );
  GTECH_OR2 C629 ( .A(N276), .B(N277), .Z(mul_out[53]) );
  GTECH_AND2 C630 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[1]), .Z(N276) );
  GTECH_AND2 C631 ( .A(m6stg_fmuls), .B(mul_frac_out[50]), .Z(N277) );
  GTECH_OR2 C632 ( .A(N278), .B(N279), .Z(mul_out[52]) );
  GTECH_AND2 C633 ( .A(m6stg_fmul_dbl_dst), .B(mul_exp_out[0]), .Z(N278) );
  GTECH_AND2 C634 ( .A(m6stg_fmuls), .B(mul_frac_out[49]), .Z(N279) );
  GTECH_OR2 C635 ( .A(N280), .B(N281), .Z(mul_out[51]) );
  GTECH_AND2 C636 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[51]), .Z(N280) );
  GTECH_AND2 C637 ( .A(m6stg_fmuls), .B(mul_frac_out[48]), .Z(N281) );
  GTECH_OR2 C638 ( .A(N282), .B(N283), .Z(mul_out[50]) );
  GTECH_AND2 C639 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[50]), .Z(N282) );
  GTECH_AND2 C640 ( .A(m6stg_fmuls), .B(mul_frac_out[47]), .Z(N283) );
  GTECH_OR2 C641 ( .A(N284), .B(N285), .Z(mul_out[49]) );
  GTECH_AND2 C642 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[49]), .Z(N284) );
  GTECH_AND2 C643 ( .A(m6stg_fmuls), .B(mul_frac_out[46]), .Z(N285) );
  GTECH_OR2 C644 ( .A(N286), .B(N287), .Z(mul_out[48]) );
  GTECH_AND2 C645 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[48]), .Z(N286) );
  GTECH_AND2 C646 ( .A(m6stg_fmuls), .B(mul_frac_out[45]), .Z(N287) );
  GTECH_OR2 C647 ( .A(N288), .B(N289), .Z(mul_out[47]) );
  GTECH_AND2 C648 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[47]), .Z(N288) );
  GTECH_AND2 C649 ( .A(m6stg_fmuls), .B(mul_frac_out[44]), .Z(N289) );
  GTECH_OR2 C650 ( .A(N290), .B(N291), .Z(mul_out[46]) );
  GTECH_AND2 C651 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[46]), .Z(N290) );
  GTECH_AND2 C652 ( .A(m6stg_fmuls), .B(mul_frac_out[43]), .Z(N291) );
  GTECH_OR2 C653 ( .A(N292), .B(N293), .Z(mul_out[45]) );
  GTECH_AND2 C654 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[45]), .Z(N292) );
  GTECH_AND2 C655 ( .A(m6stg_fmuls), .B(mul_frac_out[42]), .Z(N293) );
  GTECH_OR2 C656 ( .A(N294), .B(N295), .Z(mul_out[44]) );
  GTECH_AND2 C657 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[44]), .Z(N294) );
  GTECH_AND2 C658 ( .A(m6stg_fmuls), .B(mul_frac_out[41]), .Z(N295) );
  GTECH_OR2 C659 ( .A(N296), .B(N297), .Z(mul_out[43]) );
  GTECH_AND2 C660 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[43]), .Z(N296) );
  GTECH_AND2 C661 ( .A(m6stg_fmuls), .B(mul_frac_out[40]), .Z(N297) );
  GTECH_OR2 C662 ( .A(N298), .B(N299), .Z(mul_out[42]) );
  GTECH_AND2 C663 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[42]), .Z(N298) );
  GTECH_AND2 C664 ( .A(m6stg_fmuls), .B(mul_frac_out[39]), .Z(N299) );
  GTECH_OR2 C665 ( .A(N300), .B(N301), .Z(mul_out[41]) );
  GTECH_AND2 C666 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[41]), .Z(N300) );
  GTECH_AND2 C667 ( .A(m6stg_fmuls), .B(mul_frac_out[38]), .Z(N301) );
  GTECH_OR2 C668 ( .A(N302), .B(N303), .Z(mul_out[40]) );
  GTECH_AND2 C669 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[40]), .Z(N302) );
  GTECH_AND2 C670 ( .A(m6stg_fmuls), .B(mul_frac_out[37]), .Z(N303) );
  GTECH_OR2 C671 ( .A(N304), .B(N305), .Z(mul_out[39]) );
  GTECH_AND2 C672 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[39]), .Z(N304) );
  GTECH_AND2 C673 ( .A(m6stg_fmuls), .B(mul_frac_out[36]), .Z(N305) );
  GTECH_OR2 C674 ( .A(N306), .B(N307), .Z(mul_out[38]) );
  GTECH_AND2 C675 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[38]), .Z(N306) );
  GTECH_AND2 C676 ( .A(m6stg_fmuls), .B(mul_frac_out[35]), .Z(N307) );
  GTECH_OR2 C677 ( .A(N308), .B(N309), .Z(mul_out[37]) );
  GTECH_AND2 C678 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[37]), .Z(N308) );
  GTECH_AND2 C679 ( .A(m6stg_fmuls), .B(mul_frac_out[34]), .Z(N309) );
  GTECH_OR2 C680 ( .A(N310), .B(N311), .Z(mul_out[36]) );
  GTECH_AND2 C681 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[36]), .Z(N310) );
  GTECH_AND2 C682 ( .A(m6stg_fmuls), .B(mul_frac_out[33]), .Z(N311) );
  GTECH_OR2 C683 ( .A(N312), .B(N313), .Z(mul_out[35]) );
  GTECH_AND2 C684 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[35]), .Z(N312) );
  GTECH_AND2 C685 ( .A(m6stg_fmuls), .B(mul_frac_out[32]), .Z(N313) );
  GTECH_OR2 C686 ( .A(N314), .B(N315), .Z(mul_out[34]) );
  GTECH_AND2 C687 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[34]), .Z(N314) );
  GTECH_AND2 C688 ( .A(m6stg_fmuls), .B(mul_frac_out[31]), .Z(N315) );
  GTECH_OR2 C689 ( .A(N316), .B(N317), .Z(mul_out[33]) );
  GTECH_AND2 C690 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[33]), .Z(N316) );
  GTECH_AND2 C691 ( .A(m6stg_fmuls), .B(mul_frac_out[30]), .Z(N317) );
  GTECH_OR2 C692 ( .A(N318), .B(N319), .Z(mul_out[32]) );
  GTECH_AND2 C693 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[32]), .Z(N318) );
  GTECH_AND2 C694 ( .A(m6stg_fmuls), .B(mul_frac_out[29]), .Z(N319) );
  GTECH_AND2 C695 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[31]), .Z(
        mul_out[31]) );
  GTECH_AND2 C696 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[30]), .Z(
        mul_out[30]) );
  GTECH_AND2 C697 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[29]), .Z(
        mul_out[29]) );
  GTECH_AND2 C698 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[28]), .Z(
        mul_out[28]) );
  GTECH_AND2 C699 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[27]), .Z(
        mul_out[27]) );
  GTECH_AND2 C700 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[26]), .Z(
        mul_out[26]) );
  GTECH_AND2 C701 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[25]), .Z(
        mul_out[25]) );
  GTECH_AND2 C702 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[24]), .Z(
        mul_out[24]) );
  GTECH_AND2 C703 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[23]), .Z(
        mul_out[23]) );
  GTECH_AND2 C704 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[22]), .Z(
        mul_out[22]) );
  GTECH_AND2 C705 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[21]), .Z(
        mul_out[21]) );
  GTECH_AND2 C706 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[20]), .Z(
        mul_out[20]) );
  GTECH_AND2 C707 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[19]), .Z(
        mul_out[19]) );
  GTECH_AND2 C708 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[18]), .Z(
        mul_out[18]) );
  GTECH_AND2 C709 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[17]), .Z(
        mul_out[17]) );
  GTECH_AND2 C710 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[16]), .Z(
        mul_out[16]) );
  GTECH_AND2 C711 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[15]), .Z(
        mul_out[15]) );
  GTECH_AND2 C712 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[14]), .Z(
        mul_out[14]) );
  GTECH_AND2 C713 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[13]), .Z(
        mul_out[13]) );
  GTECH_AND2 C714 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[12]), .Z(
        mul_out[12]) );
  GTECH_AND2 C715 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[11]), .Z(
        mul_out[11]) );
  GTECH_AND2 C716 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[10]), .Z(
        mul_out[10]) );
  GTECH_AND2 C717 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[9]), .Z(mul_out[9]) );
  GTECH_AND2 C718 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[8]), .Z(mul_out[8]) );
  GTECH_AND2 C719 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[7]), .Z(mul_out[7]) );
  GTECH_AND2 C720 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[6]), .Z(mul_out[6]) );
  GTECH_AND2 C721 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[5]), .Z(mul_out[5]) );
  GTECH_AND2 C722 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[4]), .Z(mul_out[4]) );
  GTECH_AND2 C723 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[3]), .Z(mul_out[3]) );
  GTECH_AND2 C724 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[2]), .Z(mul_out[2]) );
  GTECH_AND2 C725 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[1]), .Z(mul_out[1]) );
  GTECH_AND2 C726 ( .A(m6stg_fmul_dbl_dst), .B(mul_frac_out[0]), .Z(mul_out[0]) );
  GTECH_OR2 C727 ( .A(N320), .B(N321), .Z(div_out[63]) );
  GTECH_AND2 C728 ( .A(d8stg_fdivd), .B(div_sign_out), .Z(N320) );
  GTECH_AND2 C729 ( .A(d8stg_fdivs), .B(div_sign_out), .Z(N321) );
  GTECH_OR2 C730 ( .A(N322), .B(N323), .Z(div_out[62]) );
  GTECH_AND2 C731 ( .A(d8stg_fdivd), .B(div_exp_out[10]), .Z(N322) );
  GTECH_AND2 C732 ( .A(d8stg_fdivs), .B(div_exp_out[7]), .Z(N323) );
  GTECH_OR2 C733 ( .A(N324), .B(N325), .Z(div_out[61]) );
  GTECH_AND2 C734 ( .A(d8stg_fdivd), .B(div_exp_out[9]), .Z(N324) );
  GTECH_AND2 C735 ( .A(d8stg_fdivs), .B(div_exp_out[6]), .Z(N325) );
  GTECH_OR2 C736 ( .A(N326), .B(N327), .Z(div_out[60]) );
  GTECH_AND2 C737 ( .A(d8stg_fdivd), .B(div_exp_out[8]), .Z(N326) );
  GTECH_AND2 C738 ( .A(d8stg_fdivs), .B(div_exp_out[5]), .Z(N327) );
  GTECH_OR2 C739 ( .A(N328), .B(N329), .Z(div_out[59]) );
  GTECH_AND2 C740 ( .A(d8stg_fdivd), .B(div_exp_out[7]), .Z(N328) );
  GTECH_AND2 C741 ( .A(d8stg_fdivs), .B(div_exp_out[4]), .Z(N329) );
  GTECH_OR2 C742 ( .A(N330), .B(N331), .Z(div_out[58]) );
  GTECH_AND2 C743 ( .A(d8stg_fdivd), .B(div_exp_out[6]), .Z(N330) );
  GTECH_AND2 C744 ( .A(d8stg_fdivs), .B(div_exp_out[3]), .Z(N331) );
  GTECH_OR2 C745 ( .A(N332), .B(N333), .Z(div_out[57]) );
  GTECH_AND2 C746 ( .A(d8stg_fdivd), .B(div_exp_out[5]), .Z(N332) );
  GTECH_AND2 C747 ( .A(d8stg_fdivs), .B(div_exp_out[2]), .Z(N333) );
  GTECH_OR2 C748 ( .A(N334), .B(N335), .Z(div_out[56]) );
  GTECH_AND2 C749 ( .A(d8stg_fdivd), .B(div_exp_out[4]), .Z(N334) );
  GTECH_AND2 C750 ( .A(d8stg_fdivs), .B(div_exp_out[1]), .Z(N335) );
  GTECH_OR2 C751 ( .A(N336), .B(N337), .Z(div_out[55]) );
  GTECH_AND2 C752 ( .A(d8stg_fdivd), .B(div_exp_out[3]), .Z(N336) );
  GTECH_AND2 C753 ( .A(d8stg_fdivs), .B(div_exp_out[0]), .Z(N337) );
  GTECH_OR2 C754 ( .A(N338), .B(N339), .Z(div_out[54]) );
  GTECH_AND2 C755 ( .A(d8stg_fdivd), .B(div_exp_out[2]), .Z(N338) );
  GTECH_AND2 C756 ( .A(d8stg_fdivs), .B(div_frac_out[51]), .Z(N339) );
  GTECH_OR2 C757 ( .A(N340), .B(N341), .Z(div_out[53]) );
  GTECH_AND2 C758 ( .A(d8stg_fdivd), .B(div_exp_out[1]), .Z(N340) );
  GTECH_AND2 C759 ( .A(d8stg_fdivs), .B(div_frac_out[50]), .Z(N341) );
  GTECH_OR2 C760 ( .A(N342), .B(N343), .Z(div_out[52]) );
  GTECH_AND2 C761 ( .A(d8stg_fdivd), .B(div_exp_out[0]), .Z(N342) );
  GTECH_AND2 C762 ( .A(d8stg_fdivs), .B(div_frac_out[49]), .Z(N343) );
  GTECH_OR2 C763 ( .A(N344), .B(N345), .Z(div_out[51]) );
  GTECH_AND2 C764 ( .A(d8stg_fdivd), .B(div_frac_out[51]), .Z(N344) );
  GTECH_AND2 C765 ( .A(d8stg_fdivs), .B(div_frac_out[48]), .Z(N345) );
  GTECH_OR2 C766 ( .A(N346), .B(N347), .Z(div_out[50]) );
  GTECH_AND2 C767 ( .A(d8stg_fdivd), .B(div_frac_out[50]), .Z(N346) );
  GTECH_AND2 C768 ( .A(d8stg_fdivs), .B(div_frac_out[47]), .Z(N347) );
  GTECH_OR2 C769 ( .A(N348), .B(N349), .Z(div_out[49]) );
  GTECH_AND2 C770 ( .A(d8stg_fdivd), .B(div_frac_out[49]), .Z(N348) );
  GTECH_AND2 C771 ( .A(d8stg_fdivs), .B(div_frac_out[46]), .Z(N349) );
  GTECH_OR2 C772 ( .A(N350), .B(N351), .Z(div_out[48]) );
  GTECH_AND2 C773 ( .A(d8stg_fdivd), .B(div_frac_out[48]), .Z(N350) );
  GTECH_AND2 C774 ( .A(d8stg_fdivs), .B(div_frac_out[45]), .Z(N351) );
  GTECH_OR2 C775 ( .A(N352), .B(N353), .Z(div_out[47]) );
  GTECH_AND2 C776 ( .A(d8stg_fdivd), .B(div_frac_out[47]), .Z(N352) );
  GTECH_AND2 C777 ( .A(d8stg_fdivs), .B(div_frac_out[44]), .Z(N353) );
  GTECH_OR2 C778 ( .A(N354), .B(N355), .Z(div_out[46]) );
  GTECH_AND2 C779 ( .A(d8stg_fdivd), .B(div_frac_out[46]), .Z(N354) );
  GTECH_AND2 C780 ( .A(d8stg_fdivs), .B(div_frac_out[43]), .Z(N355) );
  GTECH_OR2 C781 ( .A(N356), .B(N357), .Z(div_out[45]) );
  GTECH_AND2 C782 ( .A(d8stg_fdivd), .B(div_frac_out[45]), .Z(N356) );
  GTECH_AND2 C783 ( .A(d8stg_fdivs), .B(div_frac_out[42]), .Z(N357) );
  GTECH_OR2 C784 ( .A(N358), .B(N359), .Z(div_out[44]) );
  GTECH_AND2 C785 ( .A(d8stg_fdivd), .B(div_frac_out[44]), .Z(N358) );
  GTECH_AND2 C786 ( .A(d8stg_fdivs), .B(div_frac_out[41]), .Z(N359) );
  GTECH_OR2 C787 ( .A(N360), .B(N361), .Z(div_out[43]) );
  GTECH_AND2 C788 ( .A(d8stg_fdivd), .B(div_frac_out[43]), .Z(N360) );
  GTECH_AND2 C789 ( .A(d8stg_fdivs), .B(div_frac_out[40]), .Z(N361) );
  GTECH_OR2 C790 ( .A(N362), .B(N363), .Z(div_out[42]) );
  GTECH_AND2 C791 ( .A(d8stg_fdivd), .B(div_frac_out[42]), .Z(N362) );
  GTECH_AND2 C792 ( .A(d8stg_fdivs), .B(div_frac_out[39]), .Z(N363) );
  GTECH_OR2 C793 ( .A(N364), .B(N365), .Z(div_out[41]) );
  GTECH_AND2 C794 ( .A(d8stg_fdivd), .B(div_frac_out[41]), .Z(N364) );
  GTECH_AND2 C795 ( .A(d8stg_fdivs), .B(div_frac_out[38]), .Z(N365) );
  GTECH_OR2 C796 ( .A(N366), .B(N367), .Z(div_out[40]) );
  GTECH_AND2 C797 ( .A(d8stg_fdivd), .B(div_frac_out[40]), .Z(N366) );
  GTECH_AND2 C798 ( .A(d8stg_fdivs), .B(div_frac_out[37]), .Z(N367) );
  GTECH_OR2 C799 ( .A(N368), .B(N369), .Z(div_out[39]) );
  GTECH_AND2 C800 ( .A(d8stg_fdivd), .B(div_frac_out[39]), .Z(N368) );
  GTECH_AND2 C801 ( .A(d8stg_fdivs), .B(div_frac_out[36]), .Z(N369) );
  GTECH_OR2 C802 ( .A(N370), .B(N371), .Z(div_out[38]) );
  GTECH_AND2 C803 ( .A(d8stg_fdivd), .B(div_frac_out[38]), .Z(N370) );
  GTECH_AND2 C804 ( .A(d8stg_fdivs), .B(div_frac_out[35]), .Z(N371) );
  GTECH_OR2 C805 ( .A(N372), .B(N373), .Z(div_out[37]) );
  GTECH_AND2 C806 ( .A(d8stg_fdivd), .B(div_frac_out[37]), .Z(N372) );
  GTECH_AND2 C807 ( .A(d8stg_fdivs), .B(div_frac_out[34]), .Z(N373) );
  GTECH_OR2 C808 ( .A(N374), .B(N375), .Z(div_out[36]) );
  GTECH_AND2 C809 ( .A(d8stg_fdivd), .B(div_frac_out[36]), .Z(N374) );
  GTECH_AND2 C810 ( .A(d8stg_fdivs), .B(div_frac_out[33]), .Z(N375) );
  GTECH_OR2 C811 ( .A(N376), .B(N377), .Z(div_out[35]) );
  GTECH_AND2 C812 ( .A(d8stg_fdivd), .B(div_frac_out[35]), .Z(N376) );
  GTECH_AND2 C813 ( .A(d8stg_fdivs), .B(div_frac_out[32]), .Z(N377) );
  GTECH_OR2 C814 ( .A(N378), .B(N379), .Z(div_out[34]) );
  GTECH_AND2 C815 ( .A(d8stg_fdivd), .B(div_frac_out[34]), .Z(N378) );
  GTECH_AND2 C816 ( .A(d8stg_fdivs), .B(div_frac_out[31]), .Z(N379) );
  GTECH_OR2 C817 ( .A(N380), .B(N381), .Z(div_out[33]) );
  GTECH_AND2 C818 ( .A(d8stg_fdivd), .B(div_frac_out[33]), .Z(N380) );
  GTECH_AND2 C819 ( .A(d8stg_fdivs), .B(div_frac_out[30]), .Z(N381) );
  GTECH_OR2 C820 ( .A(N382), .B(N383), .Z(div_out[32]) );
  GTECH_AND2 C821 ( .A(d8stg_fdivd), .B(div_frac_out[32]), .Z(N382) );
  GTECH_AND2 C822 ( .A(d8stg_fdivs), .B(div_frac_out[29]), .Z(N383) );
  GTECH_AND2 C823 ( .A(d8stg_fdivd), .B(div_frac_out[31]), .Z(div_out[31]) );
  GTECH_AND2 C824 ( .A(d8stg_fdivd), .B(div_frac_out[30]), .Z(div_out[30]) );
  GTECH_AND2 C825 ( .A(d8stg_fdivd), .B(div_frac_out[29]), .Z(div_out[29]) );
  GTECH_AND2 C826 ( .A(d8stg_fdivd), .B(div_frac_out[28]), .Z(div_out[28]) );
  GTECH_AND2 C827 ( .A(d8stg_fdivd), .B(div_frac_out[27]), .Z(div_out[27]) );
  GTECH_AND2 C828 ( .A(d8stg_fdivd), .B(div_frac_out[26]), .Z(div_out[26]) );
  GTECH_AND2 C829 ( .A(d8stg_fdivd), .B(div_frac_out[25]), .Z(div_out[25]) );
  GTECH_AND2 C830 ( .A(d8stg_fdivd), .B(div_frac_out[24]), .Z(div_out[24]) );
  GTECH_AND2 C831 ( .A(d8stg_fdivd), .B(div_frac_out[23]), .Z(div_out[23]) );
  GTECH_AND2 C832 ( .A(d8stg_fdivd), .B(div_frac_out[22]), .Z(div_out[22]) );
  GTECH_AND2 C833 ( .A(d8stg_fdivd), .B(div_frac_out[21]), .Z(div_out[21]) );
  GTECH_AND2 C834 ( .A(d8stg_fdivd), .B(div_frac_out[20]), .Z(div_out[20]) );
  GTECH_AND2 C835 ( .A(d8stg_fdivd), .B(div_frac_out[19]), .Z(div_out[19]) );
  GTECH_AND2 C836 ( .A(d8stg_fdivd), .B(div_frac_out[18]), .Z(div_out[18]) );
  GTECH_AND2 C837 ( .A(d8stg_fdivd), .B(div_frac_out[17]), .Z(div_out[17]) );
  GTECH_AND2 C838 ( .A(d8stg_fdivd), .B(div_frac_out[16]), .Z(div_out[16]) );
  GTECH_AND2 C839 ( .A(d8stg_fdivd), .B(div_frac_out[15]), .Z(div_out[15]) );
  GTECH_AND2 C840 ( .A(d8stg_fdivd), .B(div_frac_out[14]), .Z(div_out[14]) );
  GTECH_AND2 C841 ( .A(d8stg_fdivd), .B(div_frac_out[13]), .Z(div_out[13]) );
  GTECH_AND2 C842 ( .A(d8stg_fdivd), .B(div_frac_out[12]), .Z(div_out[12]) );
  GTECH_AND2 C843 ( .A(d8stg_fdivd), .B(div_frac_out[11]), .Z(div_out[11]) );
  GTECH_AND2 C844 ( .A(d8stg_fdivd), .B(div_frac_out[10]), .Z(div_out[10]) );
  GTECH_AND2 C845 ( .A(d8stg_fdivd), .B(div_frac_out[9]), .Z(div_out[9]) );
  GTECH_AND2 C846 ( .A(d8stg_fdivd), .B(div_frac_out[8]), .Z(div_out[8]) );
  GTECH_AND2 C847 ( .A(d8stg_fdivd), .B(div_frac_out[7]), .Z(div_out[7]) );
  GTECH_AND2 C848 ( .A(d8stg_fdivd), .B(div_frac_out[6]), .Z(div_out[6]) );
  GTECH_AND2 C849 ( .A(d8stg_fdivd), .B(div_frac_out[5]), .Z(div_out[5]) );
  GTECH_AND2 C850 ( .A(d8stg_fdivd), .B(div_frac_out[4]), .Z(div_out[4]) );
  GTECH_AND2 C851 ( .A(d8stg_fdivd), .B(div_frac_out[3]), .Z(div_out[3]) );
  GTECH_AND2 C852 ( .A(d8stg_fdivd), .B(div_frac_out[2]), .Z(div_out[2]) );
  GTECH_AND2 C853 ( .A(d8stg_fdivd), .B(div_frac_out[1]), .Z(div_out[1]) );
  GTECH_AND2 C854 ( .A(d8stg_fdivd), .B(div_frac_out[0]), .Z(div_out[0]) );
  GTECH_OR2 C855 ( .A(N384), .B(dest_rdy[0]), .Z(fp_cpx_data_ca_84_77_in[7])
         );
  GTECH_OR2 C856 ( .A(dest_rdy[2]), .B(dest_rdy[1]), .Z(N384) );
  GTECH_OR2 C857 ( .A(N385), .B(dest_rdy[0]), .Z(fp_cpx_data_ca_84_77_in[6])
         );
  GTECH_OR2 C858 ( .A(dest_rdy[2]), .B(dest_rdy[1]), .Z(N385) );
  GTECH_AND2 C859 ( .A(N387), .B(req_thread[1]), .Z(fp_cpx_data_ca_84_77_in_1)
         );
  GTECH_OR2 C860 ( .A(N386), .B(dest_rdy[0]), .Z(N387) );
  GTECH_OR2 C861 ( .A(dest_rdy[2]), .B(dest_rdy[1]), .Z(N386) );
  GTECH_AND2 C862 ( .A(N389), .B(req_thread[0]), .Z(fp_cpx_data_ca_84_77_in_0)
         );
  GTECH_OR2 C863 ( .A(N388), .B(dest_rdy[0]), .Z(N389) );
  GTECH_OR2 C864 ( .A(dest_rdy[2]), .B(dest_rdy[1]), .Z(N388) );
  GTECH_OR2 C865 ( .A(N392), .B(N393), .Z(fp_cpx_data_ca_76_0_in_76) );
  GTECH_OR2 C866 ( .A(N390), .B(N391), .Z(N392) );
  GTECH_AND2 C867 ( .A(dest_rdy[2]), .B(div_exc_out[4]), .Z(N390) );
  GTECH_AND2 C868 ( .A(dest_rdy[1]), .B(mul_exc_out[4]), .Z(N391) );
  GTECH_AND2 C869 ( .A(dest_rdy[0]), .B(add_exc_out[4]), .Z(N393) );
  GTECH_OR2 C870 ( .A(N396), .B(N397), .Z(fp_cpx_data_ca_76_0_in_75) );
  GTECH_OR2 C871 ( .A(N394), .B(N395), .Z(N396) );
  GTECH_AND2 C872 ( .A(dest_rdy[2]), .B(div_exc_out[3]), .Z(N394) );
  GTECH_AND2 C873 ( .A(dest_rdy[1]), .B(mul_exc_out[3]), .Z(N395) );
  GTECH_AND2 C874 ( .A(dest_rdy[0]), .B(add_exc_out[3]), .Z(N397) );
  GTECH_OR2 C875 ( .A(N400), .B(N401), .Z(fp_cpx_data_ca_76_0_in_74) );
  GTECH_OR2 C876 ( .A(N398), .B(N399), .Z(N400) );
  GTECH_AND2 C877 ( .A(dest_rdy[2]), .B(div_exc_out[2]), .Z(N398) );
  GTECH_AND2 C878 ( .A(dest_rdy[1]), .B(mul_exc_out[2]), .Z(N399) );
  GTECH_AND2 C879 ( .A(dest_rdy[0]), .B(add_exc_out[2]), .Z(N401) );
  GTECH_OR2 C880 ( .A(N404), .B(N405), .Z(fp_cpx_data_ca_76_0_in_73) );
  GTECH_OR2 C881 ( .A(N402), .B(N403), .Z(N404) );
  GTECH_AND2 C882 ( .A(dest_rdy[2]), .B(div_exc_out[1]), .Z(N402) );
  GTECH_AND2 C883 ( .A(dest_rdy[1]), .B(mul_exc_out[1]), .Z(N403) );
  GTECH_AND2 C884 ( .A(dest_rdy[0]), .B(add_exc_out[1]), .Z(N405) );
  GTECH_OR2 C885 ( .A(N408), .B(N409), .Z(fp_cpx_data_ca_76_0_in_72) );
  GTECH_OR2 C886 ( .A(N406), .B(N407), .Z(N408) );
  GTECH_AND2 C887 ( .A(dest_rdy[2]), .B(div_exc_out[0]), .Z(N406) );
  GTECH_AND2 C888 ( .A(dest_rdy[1]), .B(mul_exc_out[0]), .Z(N407) );
  GTECH_AND2 C889 ( .A(dest_rdy[0]), .B(add_exc_out[0]), .Z(N409) );
  GTECH_AND2 C890 ( .A(dest_rdy[0]), .B(a6stg_fcmpop), .Z(
        fp_cpx_data_ca_76_0_in_69) );
  GTECH_AND2 C891 ( .A(dest_rdy[0]), .B(add_cc_out[1]), .Z(
        fp_cpx_data_ca_76_0_in_68) );
  GTECH_AND2 C892 ( .A(dest_rdy[0]), .B(add_cc_out[0]), .Z(
        fp_cpx_data_ca_76_0_in_67) );
  GTECH_AND2 C893 ( .A(dest_rdy[0]), .B(add_fcc_out[1]), .Z(
        fp_cpx_data_ca_76_0_in_66) );
  GTECH_AND2 C894 ( .A(dest_rdy[0]), .B(add_fcc_out[0]), .Z(
        fp_cpx_data_ca_76_0_in_65) );
  GTECH_OR2 C895 ( .A(N412), .B(N413), .Z(fp_cpx_data_ca_76_0_in[63]) );
  GTECH_OR2 C896 ( .A(N410), .B(N411), .Z(N412) );
  GTECH_AND2 C897 ( .A(dest_rdy[2]), .B(div_out[63]), .Z(N410) );
  GTECH_AND2 C898 ( .A(dest_rdy[1]), .B(mul_out[63]), .Z(N411) );
  GTECH_AND2 C899 ( .A(dest_rdy[0]), .B(add_out[63]), .Z(N413) );
  GTECH_OR2 C900 ( .A(N416), .B(N417), .Z(fp_cpx_data_ca_76_0_in[62]) );
  GTECH_OR2 C901 ( .A(N414), .B(N415), .Z(N416) );
  GTECH_AND2 C902 ( .A(dest_rdy[2]), .B(div_out[62]), .Z(N414) );
  GTECH_AND2 C903 ( .A(dest_rdy[1]), .B(mul_out[62]), .Z(N415) );
  GTECH_AND2 C904 ( .A(dest_rdy[0]), .B(add_out[62]), .Z(N417) );
  GTECH_OR2 C905 ( .A(N420), .B(N421), .Z(fp_cpx_data_ca_76_0_in[61]) );
  GTECH_OR2 C906 ( .A(N418), .B(N419), .Z(N420) );
  GTECH_AND2 C907 ( .A(dest_rdy[2]), .B(div_out[61]), .Z(N418) );
  GTECH_AND2 C908 ( .A(dest_rdy[1]), .B(mul_out[61]), .Z(N419) );
  GTECH_AND2 C909 ( .A(dest_rdy[0]), .B(add_out[61]), .Z(N421) );
  GTECH_OR2 C910 ( .A(N424), .B(N425), .Z(fp_cpx_data_ca_76_0_in[60]) );
  GTECH_OR2 C911 ( .A(N422), .B(N423), .Z(N424) );
  GTECH_AND2 C912 ( .A(dest_rdy[2]), .B(div_out[60]), .Z(N422) );
  GTECH_AND2 C913 ( .A(dest_rdy[1]), .B(mul_out[60]), .Z(N423) );
  GTECH_AND2 C914 ( .A(dest_rdy[0]), .B(add_out[60]), .Z(N425) );
  GTECH_OR2 C915 ( .A(N428), .B(N429), .Z(fp_cpx_data_ca_76_0_in[59]) );
  GTECH_OR2 C916 ( .A(N426), .B(N427), .Z(N428) );
  GTECH_AND2 C917 ( .A(dest_rdy[2]), .B(div_out[59]), .Z(N426) );
  GTECH_AND2 C918 ( .A(dest_rdy[1]), .B(mul_out[59]), .Z(N427) );
  GTECH_AND2 C919 ( .A(dest_rdy[0]), .B(add_out[59]), .Z(N429) );
  GTECH_OR2 C920 ( .A(N432), .B(N433), .Z(fp_cpx_data_ca_76_0_in[58]) );
  GTECH_OR2 C921 ( .A(N430), .B(N431), .Z(N432) );
  GTECH_AND2 C922 ( .A(dest_rdy[2]), .B(div_out[58]), .Z(N430) );
  GTECH_AND2 C923 ( .A(dest_rdy[1]), .B(mul_out[58]), .Z(N431) );
  GTECH_AND2 C924 ( .A(dest_rdy[0]), .B(add_out[58]), .Z(N433) );
  GTECH_OR2 C925 ( .A(N436), .B(N437), .Z(fp_cpx_data_ca_76_0_in[57]) );
  GTECH_OR2 C926 ( .A(N434), .B(N435), .Z(N436) );
  GTECH_AND2 C927 ( .A(dest_rdy[2]), .B(div_out[57]), .Z(N434) );
  GTECH_AND2 C928 ( .A(dest_rdy[1]), .B(mul_out[57]), .Z(N435) );
  GTECH_AND2 C929 ( .A(dest_rdy[0]), .B(add_out[57]), .Z(N437) );
  GTECH_OR2 C930 ( .A(N440), .B(N441), .Z(fp_cpx_data_ca_76_0_in[56]) );
  GTECH_OR2 C931 ( .A(N438), .B(N439), .Z(N440) );
  GTECH_AND2 C932 ( .A(dest_rdy[2]), .B(div_out[56]), .Z(N438) );
  GTECH_AND2 C933 ( .A(dest_rdy[1]), .B(mul_out[56]), .Z(N439) );
  GTECH_AND2 C934 ( .A(dest_rdy[0]), .B(add_out[56]), .Z(N441) );
  GTECH_OR2 C935 ( .A(N444), .B(N445), .Z(fp_cpx_data_ca_76_0_in[55]) );
  GTECH_OR2 C936 ( .A(N442), .B(N443), .Z(N444) );
  GTECH_AND2 C937 ( .A(dest_rdy[2]), .B(div_out[55]), .Z(N442) );
  GTECH_AND2 C938 ( .A(dest_rdy[1]), .B(mul_out[55]), .Z(N443) );
  GTECH_AND2 C939 ( .A(dest_rdy[0]), .B(add_out[55]), .Z(N445) );
  GTECH_OR2 C940 ( .A(N448), .B(N449), .Z(fp_cpx_data_ca_76_0_in[54]) );
  GTECH_OR2 C941 ( .A(N446), .B(N447), .Z(N448) );
  GTECH_AND2 C942 ( .A(dest_rdy[2]), .B(div_out[54]), .Z(N446) );
  GTECH_AND2 C943 ( .A(dest_rdy[1]), .B(mul_out[54]), .Z(N447) );
  GTECH_AND2 C944 ( .A(dest_rdy[0]), .B(add_out[54]), .Z(N449) );
  GTECH_OR2 C945 ( .A(N452), .B(N453), .Z(fp_cpx_data_ca_76_0_in[53]) );
  GTECH_OR2 C946 ( .A(N450), .B(N451), .Z(N452) );
  GTECH_AND2 C947 ( .A(dest_rdy[2]), .B(div_out[53]), .Z(N450) );
  GTECH_AND2 C948 ( .A(dest_rdy[1]), .B(mul_out[53]), .Z(N451) );
  GTECH_AND2 C949 ( .A(dest_rdy[0]), .B(add_out[53]), .Z(N453) );
  GTECH_OR2 C950 ( .A(N456), .B(N457), .Z(fp_cpx_data_ca_76_0_in[52]) );
  GTECH_OR2 C951 ( .A(N454), .B(N455), .Z(N456) );
  GTECH_AND2 C952 ( .A(dest_rdy[2]), .B(div_out[52]), .Z(N454) );
  GTECH_AND2 C953 ( .A(dest_rdy[1]), .B(mul_out[52]), .Z(N455) );
  GTECH_AND2 C954 ( .A(dest_rdy[0]), .B(add_out[52]), .Z(N457) );
  GTECH_OR2 C955 ( .A(N460), .B(N461), .Z(fp_cpx_data_ca_76_0_in[51]) );
  GTECH_OR2 C956 ( .A(N458), .B(N459), .Z(N460) );
  GTECH_AND2 C957 ( .A(dest_rdy[2]), .B(div_out[51]), .Z(N458) );
  GTECH_AND2 C958 ( .A(dest_rdy[1]), .B(mul_out[51]), .Z(N459) );
  GTECH_AND2 C959 ( .A(dest_rdy[0]), .B(add_out[51]), .Z(N461) );
  GTECH_OR2 C960 ( .A(N464), .B(N465), .Z(fp_cpx_data_ca_76_0_in[50]) );
  GTECH_OR2 C961 ( .A(N462), .B(N463), .Z(N464) );
  GTECH_AND2 C962 ( .A(dest_rdy[2]), .B(div_out[50]), .Z(N462) );
  GTECH_AND2 C963 ( .A(dest_rdy[1]), .B(mul_out[50]), .Z(N463) );
  GTECH_AND2 C964 ( .A(dest_rdy[0]), .B(add_out[50]), .Z(N465) );
  GTECH_OR2 C965 ( .A(N468), .B(N469), .Z(fp_cpx_data_ca_76_0_in[49]) );
  GTECH_OR2 C966 ( .A(N466), .B(N467), .Z(N468) );
  GTECH_AND2 C967 ( .A(dest_rdy[2]), .B(div_out[49]), .Z(N466) );
  GTECH_AND2 C968 ( .A(dest_rdy[1]), .B(mul_out[49]), .Z(N467) );
  GTECH_AND2 C969 ( .A(dest_rdy[0]), .B(add_out[49]), .Z(N469) );
  GTECH_OR2 C970 ( .A(N472), .B(N473), .Z(fp_cpx_data_ca_76_0_in[48]) );
  GTECH_OR2 C971 ( .A(N470), .B(N471), .Z(N472) );
  GTECH_AND2 C972 ( .A(dest_rdy[2]), .B(div_out[48]), .Z(N470) );
  GTECH_AND2 C973 ( .A(dest_rdy[1]), .B(mul_out[48]), .Z(N471) );
  GTECH_AND2 C974 ( .A(dest_rdy[0]), .B(add_out[48]), .Z(N473) );
  GTECH_OR2 C975 ( .A(N476), .B(N477), .Z(fp_cpx_data_ca_76_0_in[47]) );
  GTECH_OR2 C976 ( .A(N474), .B(N475), .Z(N476) );
  GTECH_AND2 C977 ( .A(dest_rdy[2]), .B(div_out[47]), .Z(N474) );
  GTECH_AND2 C978 ( .A(dest_rdy[1]), .B(mul_out[47]), .Z(N475) );
  GTECH_AND2 C979 ( .A(dest_rdy[0]), .B(add_out[47]), .Z(N477) );
  GTECH_OR2 C980 ( .A(N480), .B(N481), .Z(fp_cpx_data_ca_76_0_in[46]) );
  GTECH_OR2 C981 ( .A(N478), .B(N479), .Z(N480) );
  GTECH_AND2 C982 ( .A(dest_rdy[2]), .B(div_out[46]), .Z(N478) );
  GTECH_AND2 C983 ( .A(dest_rdy[1]), .B(mul_out[46]), .Z(N479) );
  GTECH_AND2 C984 ( .A(dest_rdy[0]), .B(add_out[46]), .Z(N481) );
  GTECH_OR2 C985 ( .A(N484), .B(N485), .Z(fp_cpx_data_ca_76_0_in[45]) );
  GTECH_OR2 C986 ( .A(N482), .B(N483), .Z(N484) );
  GTECH_AND2 C987 ( .A(dest_rdy[2]), .B(div_out[45]), .Z(N482) );
  GTECH_AND2 C988 ( .A(dest_rdy[1]), .B(mul_out[45]), .Z(N483) );
  GTECH_AND2 C989 ( .A(dest_rdy[0]), .B(add_out[45]), .Z(N485) );
  GTECH_OR2 C990 ( .A(N488), .B(N489), .Z(fp_cpx_data_ca_76_0_in[44]) );
  GTECH_OR2 C991 ( .A(N486), .B(N487), .Z(N488) );
  GTECH_AND2 C992 ( .A(dest_rdy[2]), .B(div_out[44]), .Z(N486) );
  GTECH_AND2 C993 ( .A(dest_rdy[1]), .B(mul_out[44]), .Z(N487) );
  GTECH_AND2 C994 ( .A(dest_rdy[0]), .B(add_out[44]), .Z(N489) );
  GTECH_OR2 C995 ( .A(N492), .B(N493), .Z(fp_cpx_data_ca_76_0_in[43]) );
  GTECH_OR2 C996 ( .A(N490), .B(N491), .Z(N492) );
  GTECH_AND2 C997 ( .A(dest_rdy[2]), .B(div_out[43]), .Z(N490) );
  GTECH_AND2 C998 ( .A(dest_rdy[1]), .B(mul_out[43]), .Z(N491) );
  GTECH_AND2 C999 ( .A(dest_rdy[0]), .B(add_out[43]), .Z(N493) );
  GTECH_OR2 C1000 ( .A(N496), .B(N497), .Z(fp_cpx_data_ca_76_0_in[42]) );
  GTECH_OR2 C1001 ( .A(N494), .B(N495), .Z(N496) );
  GTECH_AND2 C1002 ( .A(dest_rdy[2]), .B(div_out[42]), .Z(N494) );
  GTECH_AND2 C1003 ( .A(dest_rdy[1]), .B(mul_out[42]), .Z(N495) );
  GTECH_AND2 C1004 ( .A(dest_rdy[0]), .B(add_out[42]), .Z(N497) );
  GTECH_OR2 C1005 ( .A(N500), .B(N501), .Z(fp_cpx_data_ca_76_0_in[41]) );
  GTECH_OR2 C1006 ( .A(N498), .B(N499), .Z(N500) );
  GTECH_AND2 C1007 ( .A(dest_rdy[2]), .B(div_out[41]), .Z(N498) );
  GTECH_AND2 C1008 ( .A(dest_rdy[1]), .B(mul_out[41]), .Z(N499) );
  GTECH_AND2 C1009 ( .A(dest_rdy[0]), .B(add_out[41]), .Z(N501) );
  GTECH_OR2 C1010 ( .A(N504), .B(N505), .Z(fp_cpx_data_ca_76_0_in[40]) );
  GTECH_OR2 C1011 ( .A(N502), .B(N503), .Z(N504) );
  GTECH_AND2 C1012 ( .A(dest_rdy[2]), .B(div_out[40]), .Z(N502) );
  GTECH_AND2 C1013 ( .A(dest_rdy[1]), .B(mul_out[40]), .Z(N503) );
  GTECH_AND2 C1014 ( .A(dest_rdy[0]), .B(add_out[40]), .Z(N505) );
  GTECH_OR2 C1015 ( .A(N508), .B(N509), .Z(fp_cpx_data_ca_76_0_in[39]) );
  GTECH_OR2 C1016 ( .A(N506), .B(N507), .Z(N508) );
  GTECH_AND2 C1017 ( .A(dest_rdy[2]), .B(div_out[39]), .Z(N506) );
  GTECH_AND2 C1018 ( .A(dest_rdy[1]), .B(mul_out[39]), .Z(N507) );
  GTECH_AND2 C1019 ( .A(dest_rdy[0]), .B(add_out[39]), .Z(N509) );
  GTECH_OR2 C1020 ( .A(N512), .B(N513), .Z(fp_cpx_data_ca_76_0_in[38]) );
  GTECH_OR2 C1021 ( .A(N510), .B(N511), .Z(N512) );
  GTECH_AND2 C1022 ( .A(dest_rdy[2]), .B(div_out[38]), .Z(N510) );
  GTECH_AND2 C1023 ( .A(dest_rdy[1]), .B(mul_out[38]), .Z(N511) );
  GTECH_AND2 C1024 ( .A(dest_rdy[0]), .B(add_out[38]), .Z(N513) );
  GTECH_OR2 C1025 ( .A(N516), .B(N517), .Z(fp_cpx_data_ca_76_0_in[37]) );
  GTECH_OR2 C1026 ( .A(N514), .B(N515), .Z(N516) );
  GTECH_AND2 C1027 ( .A(dest_rdy[2]), .B(div_out[37]), .Z(N514) );
  GTECH_AND2 C1028 ( .A(dest_rdy[1]), .B(mul_out[37]), .Z(N515) );
  GTECH_AND2 C1029 ( .A(dest_rdy[0]), .B(add_out[37]), .Z(N517) );
  GTECH_OR2 C1030 ( .A(N520), .B(N521), .Z(fp_cpx_data_ca_76_0_in[36]) );
  GTECH_OR2 C1031 ( .A(N518), .B(N519), .Z(N520) );
  GTECH_AND2 C1032 ( .A(dest_rdy[2]), .B(div_out[36]), .Z(N518) );
  GTECH_AND2 C1033 ( .A(dest_rdy[1]), .B(mul_out[36]), .Z(N519) );
  GTECH_AND2 C1034 ( .A(dest_rdy[0]), .B(add_out[36]), .Z(N521) );
  GTECH_OR2 C1035 ( .A(N524), .B(N525), .Z(fp_cpx_data_ca_76_0_in[35]) );
  GTECH_OR2 C1036 ( .A(N522), .B(N523), .Z(N524) );
  GTECH_AND2 C1037 ( .A(dest_rdy[2]), .B(div_out[35]), .Z(N522) );
  GTECH_AND2 C1038 ( .A(dest_rdy[1]), .B(mul_out[35]), .Z(N523) );
  GTECH_AND2 C1039 ( .A(dest_rdy[0]), .B(add_out[35]), .Z(N525) );
  GTECH_OR2 C1040 ( .A(N528), .B(N529), .Z(fp_cpx_data_ca_76_0_in[34]) );
  GTECH_OR2 C1041 ( .A(N526), .B(N527), .Z(N528) );
  GTECH_AND2 C1042 ( .A(dest_rdy[2]), .B(div_out[34]), .Z(N526) );
  GTECH_AND2 C1043 ( .A(dest_rdy[1]), .B(mul_out[34]), .Z(N527) );
  GTECH_AND2 C1044 ( .A(dest_rdy[0]), .B(add_out[34]), .Z(N529) );
  GTECH_OR2 C1045 ( .A(N532), .B(N533), .Z(fp_cpx_data_ca_76_0_in[33]) );
  GTECH_OR2 C1046 ( .A(N530), .B(N531), .Z(N532) );
  GTECH_AND2 C1047 ( .A(dest_rdy[2]), .B(div_out[33]), .Z(N530) );
  GTECH_AND2 C1048 ( .A(dest_rdy[1]), .B(mul_out[33]), .Z(N531) );
  GTECH_AND2 C1049 ( .A(dest_rdy[0]), .B(add_out[33]), .Z(N533) );
  GTECH_OR2 C1050 ( .A(N536), .B(N537), .Z(fp_cpx_data_ca_76_0_in[32]) );
  GTECH_OR2 C1051 ( .A(N534), .B(N535), .Z(N536) );
  GTECH_AND2 C1052 ( .A(dest_rdy[2]), .B(div_out[32]), .Z(N534) );
  GTECH_AND2 C1053 ( .A(dest_rdy[1]), .B(mul_out[32]), .Z(N535) );
  GTECH_AND2 C1054 ( .A(dest_rdy[0]), .B(add_out[32]), .Z(N537) );
  GTECH_OR2 C1055 ( .A(N540), .B(N541), .Z(fp_cpx_data_ca_76_0_in[31]) );
  GTECH_OR2 C1056 ( .A(N538), .B(N539), .Z(N540) );
  GTECH_AND2 C1057 ( .A(dest_rdy[2]), .B(div_out[31]), .Z(N538) );
  GTECH_AND2 C1058 ( .A(dest_rdy[1]), .B(mul_out[31]), .Z(N539) );
  GTECH_AND2 C1059 ( .A(dest_rdy[0]), .B(add_out[31]), .Z(N541) );
  GTECH_OR2 C1060 ( .A(N544), .B(N545), .Z(fp_cpx_data_ca_76_0_in[30]) );
  GTECH_OR2 C1061 ( .A(N542), .B(N543), .Z(N544) );
  GTECH_AND2 C1062 ( .A(dest_rdy[2]), .B(div_out[30]), .Z(N542) );
  GTECH_AND2 C1063 ( .A(dest_rdy[1]), .B(mul_out[30]), .Z(N543) );
  GTECH_AND2 C1064 ( .A(dest_rdy[0]), .B(add_out[30]), .Z(N545) );
  GTECH_OR2 C1065 ( .A(N548), .B(N549), .Z(fp_cpx_data_ca_76_0_in[29]) );
  GTECH_OR2 C1066 ( .A(N546), .B(N547), .Z(N548) );
  GTECH_AND2 C1067 ( .A(dest_rdy[2]), .B(div_out[29]), .Z(N546) );
  GTECH_AND2 C1068 ( .A(dest_rdy[1]), .B(mul_out[29]), .Z(N547) );
  GTECH_AND2 C1069 ( .A(dest_rdy[0]), .B(add_out[29]), .Z(N549) );
  GTECH_OR2 C1070 ( .A(N552), .B(N553), .Z(fp_cpx_data_ca_76_0_in[28]) );
  GTECH_OR2 C1071 ( .A(N550), .B(N551), .Z(N552) );
  GTECH_AND2 C1072 ( .A(dest_rdy[2]), .B(div_out[28]), .Z(N550) );
  GTECH_AND2 C1073 ( .A(dest_rdy[1]), .B(mul_out[28]), .Z(N551) );
  GTECH_AND2 C1074 ( .A(dest_rdy[0]), .B(add_out[28]), .Z(N553) );
  GTECH_OR2 C1075 ( .A(N556), .B(N557), .Z(fp_cpx_data_ca_76_0_in[27]) );
  GTECH_OR2 C1076 ( .A(N554), .B(N555), .Z(N556) );
  GTECH_AND2 C1077 ( .A(dest_rdy[2]), .B(div_out[27]), .Z(N554) );
  GTECH_AND2 C1078 ( .A(dest_rdy[1]), .B(mul_out[27]), .Z(N555) );
  GTECH_AND2 C1079 ( .A(dest_rdy[0]), .B(add_out[27]), .Z(N557) );
  GTECH_OR2 C1080 ( .A(N560), .B(N561), .Z(fp_cpx_data_ca_76_0_in[26]) );
  GTECH_OR2 C1081 ( .A(N558), .B(N559), .Z(N560) );
  GTECH_AND2 C1082 ( .A(dest_rdy[2]), .B(div_out[26]), .Z(N558) );
  GTECH_AND2 C1083 ( .A(dest_rdy[1]), .B(mul_out[26]), .Z(N559) );
  GTECH_AND2 C1084 ( .A(dest_rdy[0]), .B(add_out[26]), .Z(N561) );
  GTECH_OR2 C1085 ( .A(N564), .B(N565), .Z(fp_cpx_data_ca_76_0_in[25]) );
  GTECH_OR2 C1086 ( .A(N562), .B(N563), .Z(N564) );
  GTECH_AND2 C1087 ( .A(dest_rdy[2]), .B(div_out[25]), .Z(N562) );
  GTECH_AND2 C1088 ( .A(dest_rdy[1]), .B(mul_out[25]), .Z(N563) );
  GTECH_AND2 C1089 ( .A(dest_rdy[0]), .B(add_out[25]), .Z(N565) );
  GTECH_OR2 C1090 ( .A(N568), .B(N569), .Z(fp_cpx_data_ca_76_0_in[24]) );
  GTECH_OR2 C1091 ( .A(N566), .B(N567), .Z(N568) );
  GTECH_AND2 C1092 ( .A(dest_rdy[2]), .B(div_out[24]), .Z(N566) );
  GTECH_AND2 C1093 ( .A(dest_rdy[1]), .B(mul_out[24]), .Z(N567) );
  GTECH_AND2 C1094 ( .A(dest_rdy[0]), .B(add_out[24]), .Z(N569) );
  GTECH_OR2 C1095 ( .A(N572), .B(N573), .Z(fp_cpx_data_ca_76_0_in[23]) );
  GTECH_OR2 C1096 ( .A(N570), .B(N571), .Z(N572) );
  GTECH_AND2 C1097 ( .A(dest_rdy[2]), .B(div_out[23]), .Z(N570) );
  GTECH_AND2 C1098 ( .A(dest_rdy[1]), .B(mul_out[23]), .Z(N571) );
  GTECH_AND2 C1099 ( .A(dest_rdy[0]), .B(add_out[23]), .Z(N573) );
  GTECH_OR2 C1100 ( .A(N576), .B(N577), .Z(fp_cpx_data_ca_76_0_in[22]) );
  GTECH_OR2 C1101 ( .A(N574), .B(N575), .Z(N576) );
  GTECH_AND2 C1102 ( .A(dest_rdy[2]), .B(div_out[22]), .Z(N574) );
  GTECH_AND2 C1103 ( .A(dest_rdy[1]), .B(mul_out[22]), .Z(N575) );
  GTECH_AND2 C1104 ( .A(dest_rdy[0]), .B(add_out[22]), .Z(N577) );
  GTECH_OR2 C1105 ( .A(N580), .B(N581), .Z(fp_cpx_data_ca_76_0_in[21]) );
  GTECH_OR2 C1106 ( .A(N578), .B(N579), .Z(N580) );
  GTECH_AND2 C1107 ( .A(dest_rdy[2]), .B(div_out[21]), .Z(N578) );
  GTECH_AND2 C1108 ( .A(dest_rdy[1]), .B(mul_out[21]), .Z(N579) );
  GTECH_AND2 C1109 ( .A(dest_rdy[0]), .B(add_out[21]), .Z(N581) );
  GTECH_OR2 C1110 ( .A(N584), .B(N585), .Z(fp_cpx_data_ca_76_0_in[20]) );
  GTECH_OR2 C1111 ( .A(N582), .B(N583), .Z(N584) );
  GTECH_AND2 C1112 ( .A(dest_rdy[2]), .B(div_out[20]), .Z(N582) );
  GTECH_AND2 C1113 ( .A(dest_rdy[1]), .B(mul_out[20]), .Z(N583) );
  GTECH_AND2 C1114 ( .A(dest_rdy[0]), .B(add_out[20]), .Z(N585) );
  GTECH_OR2 C1115 ( .A(N588), .B(N589), .Z(fp_cpx_data_ca_76_0_in[19]) );
  GTECH_OR2 C1116 ( .A(N586), .B(N587), .Z(N588) );
  GTECH_AND2 C1117 ( .A(dest_rdy[2]), .B(div_out[19]), .Z(N586) );
  GTECH_AND2 C1118 ( .A(dest_rdy[1]), .B(mul_out[19]), .Z(N587) );
  GTECH_AND2 C1119 ( .A(dest_rdy[0]), .B(add_out[19]), .Z(N589) );
  GTECH_OR2 C1120 ( .A(N592), .B(N593), .Z(fp_cpx_data_ca_76_0_in[18]) );
  GTECH_OR2 C1121 ( .A(N590), .B(N591), .Z(N592) );
  GTECH_AND2 C1122 ( .A(dest_rdy[2]), .B(div_out[18]), .Z(N590) );
  GTECH_AND2 C1123 ( .A(dest_rdy[1]), .B(mul_out[18]), .Z(N591) );
  GTECH_AND2 C1124 ( .A(dest_rdy[0]), .B(add_out[18]), .Z(N593) );
  GTECH_OR2 C1125 ( .A(N596), .B(N597), .Z(fp_cpx_data_ca_76_0_in[17]) );
  GTECH_OR2 C1126 ( .A(N594), .B(N595), .Z(N596) );
  GTECH_AND2 C1127 ( .A(dest_rdy[2]), .B(div_out[17]), .Z(N594) );
  GTECH_AND2 C1128 ( .A(dest_rdy[1]), .B(mul_out[17]), .Z(N595) );
  GTECH_AND2 C1129 ( .A(dest_rdy[0]), .B(add_out[17]), .Z(N597) );
  GTECH_OR2 C1130 ( .A(N600), .B(N601), .Z(fp_cpx_data_ca_76_0_in[16]) );
  GTECH_OR2 C1131 ( .A(N598), .B(N599), .Z(N600) );
  GTECH_AND2 C1132 ( .A(dest_rdy[2]), .B(div_out[16]), .Z(N598) );
  GTECH_AND2 C1133 ( .A(dest_rdy[1]), .B(mul_out[16]), .Z(N599) );
  GTECH_AND2 C1134 ( .A(dest_rdy[0]), .B(add_out[16]), .Z(N601) );
  GTECH_OR2 C1135 ( .A(N604), .B(N605), .Z(fp_cpx_data_ca_76_0_in[15]) );
  GTECH_OR2 C1136 ( .A(N602), .B(N603), .Z(N604) );
  GTECH_AND2 C1137 ( .A(dest_rdy[2]), .B(div_out[15]), .Z(N602) );
  GTECH_AND2 C1138 ( .A(dest_rdy[1]), .B(mul_out[15]), .Z(N603) );
  GTECH_AND2 C1139 ( .A(dest_rdy[0]), .B(add_out[15]), .Z(N605) );
  GTECH_OR2 C1140 ( .A(N608), .B(N609), .Z(fp_cpx_data_ca_76_0_in[14]) );
  GTECH_OR2 C1141 ( .A(N606), .B(N607), .Z(N608) );
  GTECH_AND2 C1142 ( .A(dest_rdy[2]), .B(div_out[14]), .Z(N606) );
  GTECH_AND2 C1143 ( .A(dest_rdy[1]), .B(mul_out[14]), .Z(N607) );
  GTECH_AND2 C1144 ( .A(dest_rdy[0]), .B(add_out[14]), .Z(N609) );
  GTECH_OR2 C1145 ( .A(N612), .B(N613), .Z(fp_cpx_data_ca_76_0_in[13]) );
  GTECH_OR2 C1146 ( .A(N610), .B(N611), .Z(N612) );
  GTECH_AND2 C1147 ( .A(dest_rdy[2]), .B(div_out[13]), .Z(N610) );
  GTECH_AND2 C1148 ( .A(dest_rdy[1]), .B(mul_out[13]), .Z(N611) );
  GTECH_AND2 C1149 ( .A(dest_rdy[0]), .B(add_out[13]), .Z(N613) );
  GTECH_OR2 C1150 ( .A(N616), .B(N617), .Z(fp_cpx_data_ca_76_0_in[12]) );
  GTECH_OR2 C1151 ( .A(N614), .B(N615), .Z(N616) );
  GTECH_AND2 C1152 ( .A(dest_rdy[2]), .B(div_out[12]), .Z(N614) );
  GTECH_AND2 C1153 ( .A(dest_rdy[1]), .B(mul_out[12]), .Z(N615) );
  GTECH_AND2 C1154 ( .A(dest_rdy[0]), .B(add_out[12]), .Z(N617) );
  GTECH_OR2 C1155 ( .A(N620), .B(N621), .Z(fp_cpx_data_ca_76_0_in[11]) );
  GTECH_OR2 C1156 ( .A(N618), .B(N619), .Z(N620) );
  GTECH_AND2 C1157 ( .A(dest_rdy[2]), .B(div_out[11]), .Z(N618) );
  GTECH_AND2 C1158 ( .A(dest_rdy[1]), .B(mul_out[11]), .Z(N619) );
  GTECH_AND2 C1159 ( .A(dest_rdy[0]), .B(add_out[11]), .Z(N621) );
  GTECH_OR2 C1160 ( .A(N624), .B(N625), .Z(fp_cpx_data_ca_76_0_in[10]) );
  GTECH_OR2 C1161 ( .A(N622), .B(N623), .Z(N624) );
  GTECH_AND2 C1162 ( .A(dest_rdy[2]), .B(div_out[10]), .Z(N622) );
  GTECH_AND2 C1163 ( .A(dest_rdy[1]), .B(mul_out[10]), .Z(N623) );
  GTECH_AND2 C1164 ( .A(dest_rdy[0]), .B(add_out[10]), .Z(N625) );
  GTECH_OR2 C1165 ( .A(N628), .B(N629), .Z(fp_cpx_data_ca_76_0_in[9]) );
  GTECH_OR2 C1166 ( .A(N626), .B(N627), .Z(N628) );
  GTECH_AND2 C1167 ( .A(dest_rdy[2]), .B(div_out[9]), .Z(N626) );
  GTECH_AND2 C1168 ( .A(dest_rdy[1]), .B(mul_out[9]), .Z(N627) );
  GTECH_AND2 C1169 ( .A(dest_rdy[0]), .B(add_out[9]), .Z(N629) );
  GTECH_OR2 C1170 ( .A(N632), .B(N633), .Z(fp_cpx_data_ca_76_0_in[8]) );
  GTECH_OR2 C1171 ( .A(N630), .B(N631), .Z(N632) );
  GTECH_AND2 C1172 ( .A(dest_rdy[2]), .B(div_out[8]), .Z(N630) );
  GTECH_AND2 C1173 ( .A(dest_rdy[1]), .B(mul_out[8]), .Z(N631) );
  GTECH_AND2 C1174 ( .A(dest_rdy[0]), .B(add_out[8]), .Z(N633) );
  GTECH_OR2 C1175 ( .A(N636), .B(N637), .Z(fp_cpx_data_ca_76_0_in[7]) );
  GTECH_OR2 C1176 ( .A(N634), .B(N635), .Z(N636) );
  GTECH_AND2 C1177 ( .A(dest_rdy[2]), .B(div_out[7]), .Z(N634) );
  GTECH_AND2 C1178 ( .A(dest_rdy[1]), .B(mul_out[7]), .Z(N635) );
  GTECH_AND2 C1179 ( .A(dest_rdy[0]), .B(add_out[7]), .Z(N637) );
  GTECH_OR2 C1180 ( .A(N640), .B(N641), .Z(fp_cpx_data_ca_76_0_in[6]) );
  GTECH_OR2 C1181 ( .A(N638), .B(N639), .Z(N640) );
  GTECH_AND2 C1182 ( .A(dest_rdy[2]), .B(div_out[6]), .Z(N638) );
  GTECH_AND2 C1183 ( .A(dest_rdy[1]), .B(mul_out[6]), .Z(N639) );
  GTECH_AND2 C1184 ( .A(dest_rdy[0]), .B(add_out[6]), .Z(N641) );
  GTECH_OR2 C1185 ( .A(N644), .B(N645), .Z(fp_cpx_data_ca_76_0_in[5]) );
  GTECH_OR2 C1186 ( .A(N642), .B(N643), .Z(N644) );
  GTECH_AND2 C1187 ( .A(dest_rdy[2]), .B(div_out[5]), .Z(N642) );
  GTECH_AND2 C1188 ( .A(dest_rdy[1]), .B(mul_out[5]), .Z(N643) );
  GTECH_AND2 C1189 ( .A(dest_rdy[0]), .B(add_out[5]), .Z(N645) );
  GTECH_OR2 C1190 ( .A(N648), .B(N649), .Z(fp_cpx_data_ca_76_0_in[4]) );
  GTECH_OR2 C1191 ( .A(N646), .B(N647), .Z(N648) );
  GTECH_AND2 C1192 ( .A(dest_rdy[2]), .B(div_out[4]), .Z(N646) );
  GTECH_AND2 C1193 ( .A(dest_rdy[1]), .B(mul_out[4]), .Z(N647) );
  GTECH_AND2 C1194 ( .A(dest_rdy[0]), .B(add_out[4]), .Z(N649) );
  GTECH_OR2 C1195 ( .A(N652), .B(N653), .Z(fp_cpx_data_ca_76_0_in[3]) );
  GTECH_OR2 C1196 ( .A(N650), .B(N651), .Z(N652) );
  GTECH_AND2 C1197 ( .A(dest_rdy[2]), .B(div_out[3]), .Z(N650) );
  GTECH_AND2 C1198 ( .A(dest_rdy[1]), .B(mul_out[3]), .Z(N651) );
  GTECH_AND2 C1199 ( .A(dest_rdy[0]), .B(add_out[3]), .Z(N653) );
  GTECH_OR2 C1200 ( .A(N656), .B(N657), .Z(fp_cpx_data_ca_76_0_in[2]) );
  GTECH_OR2 C1201 ( .A(N654), .B(N655), .Z(N656) );
  GTECH_AND2 C1202 ( .A(dest_rdy[2]), .B(div_out[2]), .Z(N654) );
  GTECH_AND2 C1203 ( .A(dest_rdy[1]), .B(mul_out[2]), .Z(N655) );
  GTECH_AND2 C1204 ( .A(dest_rdy[0]), .B(add_out[2]), .Z(N657) );
  GTECH_OR2 C1205 ( .A(N660), .B(N661), .Z(fp_cpx_data_ca_76_0_in[1]) );
  GTECH_OR2 C1206 ( .A(N658), .B(N659), .Z(N660) );
  GTECH_AND2 C1207 ( .A(dest_rdy[2]), .B(div_out[1]), .Z(N658) );
  GTECH_AND2 C1208 ( .A(dest_rdy[1]), .B(mul_out[1]), .Z(N659) );
  GTECH_AND2 C1209 ( .A(dest_rdy[0]), .B(add_out[1]), .Z(N661) );
  GTECH_OR2 C1210 ( .A(N664), .B(N665), .Z(fp_cpx_data_ca_76_0_in[0]) );
  GTECH_OR2 C1211 ( .A(N662), .B(N663), .Z(N664) );
  GTECH_AND2 C1212 ( .A(dest_rdy[2]), .B(div_out[0]), .Z(N662) );
  GTECH_AND2 C1213 ( .A(dest_rdy[1]), .B(mul_out[0]), .Z(N663) );
  GTECH_AND2 C1214 ( .A(dest_rdy[0]), .B(add_out[0]), .Z(N665) );
endmodule


module fpu_out ( d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, div_id_out_in, 
        m6stg_id_in, add_id_out_in, div_exc_out, d8stg_fdivd, d8stg_fdivs, 
        div_sign_out, div_exp_out, div_frac_out, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, add_exc_out, a6stg_fcmpop, add_cc_out, add_fcc_out, 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        add_sign_out, add_exp_out, add_frac_out, arst_l, grst_l, rclk, 
        fp_cpx_req_cq, add_dest_rdy, mul_dest_rdy, div_dest_rdy, 
        fp_cpx_data_ca, se, si, so );
  input [9:0] div_id_out_in;
  input [9:0] m6stg_id_in;
  input [9:0] add_id_out_in;
  input [4:0] div_exc_out;
  input [10:0] div_exp_out;
  input [51:0] div_frac_out;
  input [4:0] mul_exc_out;
  input [10:0] mul_exp_out;
  input [51:0] mul_frac_out;
  input [4:0] add_exc_out;
  input [1:0] add_cc_out;
  input [1:0] add_fcc_out;
  input [10:0] add_exp_out;
  input [63:0] add_frac_out;
  output [7:0] fp_cpx_req_cq;
  output [144:0] fp_cpx_data_ca;
  input d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out,
         a6stg_fcmpop, a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst,
         a6stg_int_dst, add_sign_out, arst_l, grst_l, rclk, se, si;
  output add_dest_rdy, mul_dest_rdy, div_dest_rdy, so;
  wire   scan_out_fpu_out_ctl;
  wire   [1:0] req_thread;
  wire   [2:0] dest_rdy;

  fpu_out_ctl fpu_out_ctl ( .d8stg_fdiv_in(d8stg_fdiv_in), .m6stg_fmul_in(
        m6stg_fmul_in), .a6stg_fadd_in(a6stg_fadd_in), .div_id_out_in(
        div_id_out_in), .m6stg_id_in(m6stg_id_in), .add_id_out_in(
        add_id_out_in), .arst_l(arst_l), .grst_l(grst_l), .rclk(rclk), 
        .fp_cpx_req_cq(fp_cpx_req_cq), .req_thread(req_thread), .dest_rdy(
        dest_rdy), .add_dest_rdy(add_dest_rdy), .mul_dest_rdy(mul_dest_rdy), 
        .div_dest_rdy(div_dest_rdy), .se(se), .si(si), .so(
        scan_out_fpu_out_ctl) );
  fpu_out_dp fpu_out_dp ( .dest_rdy(dest_rdy), .req_thread(req_thread), 
        .div_exc_out(div_exc_out), .d8stg_fdivd(d8stg_fdivd), .d8stg_fdivs(
        d8stg_fdivs), .div_sign_out(div_sign_out), .div_exp_out(div_exp_out), 
        .div_frac_out(div_frac_out), .mul_exc_out(mul_exc_out), 
        .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), .m6stg_fmuls(m6stg_fmuls), 
        .mul_sign_out(mul_sign_out), .mul_exp_out(mul_exp_out), .mul_frac_out(
        mul_frac_out), .add_exc_out(add_exc_out), .a6stg_fcmpop(a6stg_fcmpop), 
        .add_cc_out(add_cc_out), .add_fcc_out(add_fcc_out), .a6stg_dbl_dst(
        a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), .a6stg_long_dst(
        a6stg_long_dst), .a6stg_int_dst(a6stg_int_dst), .add_sign_out(
        add_sign_out), .add_exp_out(add_exp_out), .add_frac_out(add_frac_out), 
        .rclk(rclk), .fp_cpx_data_ca(fp_cpx_data_ca), .se(se), .si(
        scan_out_fpu_out_ctl), .so(so) );
endmodule


module test_stub_scan ( mux_drive_disable, mem_write_disable, sehold, se, 
        testmode_l, mem_bypass, so_0, so_1, so_2, ctu_tst_pre_grst_l, arst_l, 
        global_shift_enable, ctu_tst_scan_disable, ctu_tst_scanmode, 
        ctu_tst_macrotest, ctu_tst_short_chain, long_chain_so_0, 
        short_chain_so_0, long_chain_so_1, short_chain_so_1, long_chain_so_2, 
        short_chain_so_2 );
  input ctu_tst_pre_grst_l, arst_l, global_shift_enable, ctu_tst_scan_disable,
         ctu_tst_scanmode, ctu_tst_macrotest, ctu_tst_short_chain,
         long_chain_so_0, short_chain_so_0, long_chain_so_1, short_chain_so_1,
         long_chain_so_2, short_chain_so_2;
  output mux_drive_disable, mem_write_disable, sehold, se, testmode_l,
         mem_bypass, so_0, so_1, so_2;
  wire   N0, N1, se, short_chain_select, short_chain_en, N2, N3, N4, N5, N6,
         N7, N8, N9;
  assign se = global_shift_enable;

  SELECT_OP C30 ( .DATA1(short_chain_so_0), .DATA2(long_chain_so_0), 
        .CONTROL1(N0), .CONTROL2(N1), .Z(so_0) );
  GTECH_BUF B_0 ( .A(short_chain_select), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  SELECT_OP C31 ( .DATA1(short_chain_so_1), .DATA2(long_chain_so_1), 
        .CONTROL1(N0), .CONTROL2(N1), .Z(so_1) );
  SELECT_OP C32 ( .DATA1(short_chain_so_2), .DATA2(long_chain_so_2), 
        .CONTROL1(N0), .CONTROL2(N1), .Z(so_2) );
  GTECH_OR2 C34 ( .A(N4), .B(se), .Z(mux_drive_disable) );
  GTECH_OR2 C35 ( .A(N3), .B(short_chain_select), .Z(N4) );
  GTECH_NOT I_0 ( .A(ctu_tst_pre_grst_l), .Z(N3) );
  GTECH_OR2 C37 ( .A(N3), .B(se), .Z(mem_write_disable) );
  GTECH_AND2 C39 ( .A(ctu_tst_macrotest), .B(N5), .Z(sehold) );
  GTECH_NOT I_1 ( .A(se), .Z(N5) );
  GTECH_NOT I_2 ( .A(ctu_tst_scanmode), .Z(testmode_l) );
  GTECH_AND2 C42 ( .A(N6), .B(N7), .Z(mem_bypass) );
  GTECH_NOT I_3 ( .A(ctu_tst_macrotest), .Z(N6) );
  GTECH_NOT I_4 ( .A(testmode_l), .Z(N7) );
  GTECH_NOT I_5 ( .A(N8), .Z(short_chain_en) );
  GTECH_AND2 C46 ( .A(ctu_tst_scan_disable), .B(se), .Z(N8) );
  GTECH_AND2 C47 ( .A(N9), .B(short_chain_en), .Z(short_chain_select) );
  GTECH_AND2 C48 ( .A(ctu_tst_short_chain), .B(N7), .Z(N9) );
  GTECH_NOT I_6 ( .A(short_chain_select), .Z(N2) );
endmodule


module bw_u1_syncff_4x ( q, so, ck, d, se, sd );
  input ck, d, se, sd;
  output q, so;
  wire   N0, N1, q, N2, N3;
  assign so = q;

  \**SEQGEN**  q_r_reg ( .clear(1'b0), .preset(1'b0), .next_state(N3), 
        .clocked_on(ck), .data_in(1'b0), .enable(1'b0), .Q(q), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1)
         );
  SELECT_OP C11 ( .DATA1(sd), .DATA2(d), .CONTROL1(N0), .CONTROL2(N1), .Z(N3)
         );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  GTECH_NOT I_0 ( .A(se), .Z(N2) );
endmodule


module bw_u1_scanl_2x ( so, sd, ck );
  input sd, ck;
  output so;
  wire   so_l, N0, N1;

  \**SEQGEN**  so_l_reg ( .clear(1'b0), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(1'b0), .data_in(N1), .enable(N0), .Q(so_l), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b0)
         );
  GTECH_NOT I_0 ( .A(so_l), .Z(so) );
  GTECH_NOT I_1 ( .A(ck), .Z(N0) );
  GTECH_NOT I_2 ( .A(sd), .Z(N1) );
endmodule


module zsoffasr_prim ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12;

  \**SEQGEN**  q_reg ( .clear(N5), .preset(1'b0), .next_state(N10), 
        .clocked_on(ck), .data_in(r_l), .enable(N11), .Q(q), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1) );
  GTECH_NOT I_0 ( .A(s_l), .Z(N6) );
  SELECT_OP C33 ( .DATA1(N8), .DATA2(N9), .CONTROL1(N0), .CONTROL2(N1), .Z(N10) );
  GTECH_BUF B_0 ( .A(se), .Z(N0) );
  GTECH_BUF B_1 ( .A(N7), .Z(N1) );
  SELECT_OP C34 ( .DATA1(1'b1), .DATA2(1'b0), .CONTROL1(N2), .CONTROL2(N3), 
        .Z(N11) );
  GTECH_BUF B_2 ( .A(N6), .Z(N2) );
  GTECH_BUF B_3 ( .A(s_l), .Z(N3) );
  GTECH_AND2 C37 ( .A(r_l), .B(s_l), .Z(N4) );
  GTECH_NOT I_1 ( .A(r_l), .Z(N5) );
  GTECH_NOT I_2 ( .A(se), .Z(N7) );
  GTECH_AND2 C42 ( .A(N4), .B(sd), .Z(N8) );
  GTECH_AND2 C43 ( .A(N12), .B(d), .Z(N9) );
  GTECH_AND2 C44 ( .A(N4), .B(N7), .Z(N12) );
  GTECH_OR2 C46 ( .A(q), .B(N7), .Z(so) );
endmodule


module bw_u1_soffasr_2x ( q, so, ck, d, r_l, s_l, se, sd );
  input ck, d, r_l, s_l, se, sd;
  output q, so;


  zsoffasr_prim i0 ( .q(q), .so(so), .ck(ck), .d(d), .r_l(r_l), .s_l(s_l), 
        .se(se), .sd(sd) );
endmodule


module synchronizer_asr ( sync_out, so, async_in, gclk, rclk, arst_l, si, se
 );
  input async_in, gclk, rclk, arst_l, si, se;
  output sync_out, so;
  wire   pre_sync_out, so_rptr, so_lockup;

  bw_u1_soffasr_2x repeater ( .q(pre_sync_out), .so(so_rptr), .ck(gclk), .d(
        async_in), .r_l(arst_l), .s_l(1'b1), .se(se), .sd(si) );
  bw_u1_scanl_2x lockup ( .so(so_lockup), .sd(so_rptr), .ck(gclk) );
  bw_u1_soffasr_2x syncff ( .q(sync_out), .so(so), .ck(rclk), .d(pre_sync_out), 
        .r_l(arst_l), .s_l(1'b1), .se(se), .sd(so_lockup) );
endmodule


module cluster_header ( dbginit_l, cluster_grst_l, rclk, so, gclk, 
        cluster_cken, arst_l, grst_l, adbginit_l, gdbginit_l, si, se );
  input gclk, cluster_cken, arst_l, grst_l, adbginit_l, gdbginit_l, si, se;
  output dbginit_l, cluster_grst_l, rclk, so;
  wire   pre_sync_enable, sync_enable, rst_sync_so;

  bw_u1_syncff_4x sync_cluster_master ( .q(pre_sync_enable), .ck(gclk), .d(
        cluster_cken), .se(1'b0), .sd(1'b0) );
  bw_u1_scanl_2x sync_cluster_slave ( .so(sync_enable), .sd(pre_sync_enable), 
        .ck(gclk) );
  synchronizer_asr rst_repeater ( .sync_out(cluster_grst_l), .so(rst_sync_so), 
        .async_in(grst_l), .gclk(gclk), .rclk(rclk), .arst_l(arst_l), .si(si), 
        .se(se) );
  synchronizer_asr dbginit_repeater ( .sync_out(dbginit_l), .so(so), 
        .async_in(gdbginit_l), .gclk(gclk), .rclk(rclk), .arst_l(adbginit_l), 
        .si(rst_sync_so), .se(se) );
  GTECH_AND2 C8 ( .A(gclk), .B(sync_enable), .Z(rclk) );
endmodule


module bw_clk_cl_fpu_cmp ( so, dbginit_l, cluster_grst_l, rclk, si, se, 
        adbginit_l, gdbginit_l, arst_l, grst_l, cluster_cken, gclk );
  input si, se, adbginit_l, gdbginit_l, arst_l, grst_l, cluster_cken, gclk;
  output so, dbginit_l, cluster_grst_l, rclk;


  cluster_header I0 ( .dbginit_l(dbginit_l), .cluster_grst_l(cluster_grst_l), 
        .rclk(rclk), .so(so), .gclk(gclk), .cluster_cken(cluster_cken), 
        .arst_l(arst_l), .grst_l(grst_l), .adbginit_l(adbginit_l), 
        .gdbginit_l(gdbginit_l), .si(si), .se(se) );
endmodule


module fpu_bufrpt_grp32 ( in, out );
  input [31:0] in;
  output [31:0] out;

  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp64 ( in, out );
  input [63:0] in;
  output [63:0] out;

  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[55];
  assign out[54] = in[54];
  assign out[53] = in[53];
  assign out[52] = in[52];
  assign out[51] = in[51];
  assign out[50] = in[50];
  assign out[49] = in[49];
  assign out[48] = in[48];
  assign out[47] = in[47];
  assign out[46] = in[46];
  assign out[45] = in[45];
  assign out[44] = in[44];
  assign out[43] = in[43];
  assign out[42] = in[42];
  assign out[41] = in[41];
  assign out[40] = in[40];
  assign out[39] = in[39];
  assign out[38] = in[38];
  assign out[37] = in[37];
  assign out[36] = in[36];
  assign out[35] = in[35];
  assign out[34] = in[34];
  assign out[33] = in[33];
  assign out[32] = in[32];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_bufrpt_grp4 ( in, out );
  input [3:0] in;
  output [3:0] out;

  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_pcx_fpio_grp16 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_fp_cpx_grp16 ( in, out );
  input [15:0] in;
  output [15:0] out;

  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_inq ( in, out );
  input [155:0] in;
  output [155:0] out;

  assign out[155] = in[155];
  assign out[154] = in[154];
  assign out[153] = in[153];
  assign out[152] = in[152];
  assign out[151] = in[151];
  assign out[150] = in[150];
  assign out[149] = in[149];
  assign out[148] = in[148];
  assign out[147] = in[147];
  assign out[146] = in[146];
  assign out[145] = in[145];
  assign out[144] = in[144];
  assign out[143] = in[143];
  assign out[142] = in[142];
  assign out[141] = in[141];
  assign out[140] = in[140];
  assign out[139] = in[139];
  assign out[138] = in[138];
  assign out[137] = in[137];
  assign out[136] = in[136];
  assign out[135] = in[135];
  assign out[134] = in[134];
  assign out[133] = in[133];
  assign out[132] = in[132];
  assign out[131] = in[131];
  assign out[130] = in[130];
  assign out[129] = in[129];
  assign out[128] = in[128];
  assign out[127] = in[127];
  assign out[126] = in[126];
  assign out[125] = in[125];
  assign out[124] = in[124];
  assign out[123] = in[123];
  assign out[122] = in[122];
  assign out[121] = in[121];
  assign out[120] = in[120];
  assign out[119] = in[119];
  assign out[118] = in[118];
  assign out[117] = in[117];
  assign out[116] = in[116];
  assign out[115] = in[115];
  assign out[114] = in[114];
  assign out[113] = in[113];
  assign out[112] = in[112];
  assign out[111] = in[111];
  assign out[110] = in[110];
  assign out[109] = in[109];
  assign out[108] = in[108];
  assign out[107] = in[107];
  assign out[106] = in[106];
  assign out[105] = in[105];
  assign out[104] = in[104];
  assign out[103] = in[103];
  assign out[102] = in[102];
  assign out[101] = in[101];
  assign out[100] = in[100];
  assign out[99] = in[99];
  assign out[98] = in[98];
  assign out[97] = in[97];
  assign out[96] = in[96];
  assign out[95] = in[95];
  assign out[94] = in[94];
  assign out[93] = in[93];
  assign out[92] = in[92];
  assign out[91] = in[91];
  assign out[90] = in[90];
  assign out[89] = in[89];
  assign out[88] = in[88];
  assign out[87] = in[87];
  assign out[86] = in[86];
  assign out[85] = in[85];
  assign out[84] = in[84];
  assign out[83] = in[83];
  assign out[82] = in[82];
  assign out[81] = in[81];
  assign out[80] = in[80];
  assign out[79] = in[79];
  assign out[78] = in[78];
  assign out[77] = in[77];
  assign out[76] = in[76];
  assign out[75] = in[75];
  assign out[74] = in[74];
  assign out[73] = in[73];
  assign out[72] = in[72];
  assign out[71] = in[71];
  assign out[70] = in[70];
  assign out[69] = in[69];
  assign out[68] = in[68];
  assign out[67] = in[67];
  assign out[66] = in[66];
  assign out[65] = in[65];
  assign out[64] = in[64];
  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[55];
  assign out[54] = in[54];
  assign out[53] = in[53];
  assign out[52] = in[52];
  assign out[51] = in[51];
  assign out[50] = in[50];
  assign out[49] = in[49];
  assign out[48] = in[48];
  assign out[47] = in[47];
  assign out[46] = in[46];
  assign out[45] = in[45];
  assign out[44] = in[44];
  assign out[43] = in[43];
  assign out[42] = in[42];
  assign out[41] = in[41];
  assign out[40] = in[40];
  assign out[39] = in[39];
  assign out[38] = in[38];
  assign out[37] = in[37];
  assign out[36] = in[36];
  assign out[35] = in[35];
  assign out[34] = in[34];
  assign out[33] = in[33];
  assign out[32] = in[32];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[23];
  assign out[22] = in[22];
  assign out[21] = in[21];
  assign out[20] = in[20];
  assign out[19] = in[19];
  assign out[18] = in[18];
  assign out[17] = in[17];
  assign out[16] = in[16];
  assign out[15] = in[15];
  assign out[14] = in[14];
  assign out[13] = in[13];
  assign out[12] = in[12];
  assign out[11] = in[11];
  assign out[10] = in[10];
  assign out[9] = in[9];
  assign out[8] = in[8];
  assign out[7] = in[7];
  assign out[6] = in[6];
  assign out[5] = in[5];
  assign out[4] = in[4];
  assign out[3] = in[3];
  assign out[2] = in[2];
  assign out[1] = in[1];
  assign out[0] = in[0];

endmodule


module fpu_rptr_groups ( inq_in1, inq_in2, inq_id, inq_op, inq_rnd_mode, 
        inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0, 
        inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, 
        inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l, 
        ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain, 
        global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l, 
        fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf, 
        pcx_fpio_data_px2, pcx_fpio_data_rdy_px2, fp_cpx_req_cq, 
        fp_cpx_data_ca, inq_sram_din_unbuf, inq_in1_add_buf1, inq_in1_mul_buf1, 
        inq_in1_div_buf1, inq_in2_add_buf1, inq_in2_mul_buf1, inq_in2_div_buf1, 
        inq_id_add_buf1, inq_id_mul_buf1, inq_id_div_buf1, inq_op_add_buf1, 
        inq_op_div_buf1, inq_op_mul_buf1, inq_rnd_mode_add_buf1, 
        inq_rnd_mode_div_buf1, inq_rnd_mode_mul_buf1, 
        inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1, 
        inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1, 
        inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1, 
        inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1, 
        inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1, 
        inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1, 
        inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1, 
        inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1, 
        inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1, 
        inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1, 
        inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1, 
        inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1, 
        inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1, 
        inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1, 
        inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1, 
        ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1, 
        ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1, 
        ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1, 
        cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2, 
        se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4, 
        se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2, 
        arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3, 
        arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2, 
        fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1, 
        fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so, 
        pcx_fpio_data_px2_buf1, pcx_fpio_data_rdy_px2_buf1, fp_cpx_req_cq_buf1, 
        fp_cpx_data_ca_buf1, inq_sram_din_buf1 );
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  input [4:0] inq_id;
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [123:0] pcx_fpio_data_px2;
  input [7:0] fp_cpx_req_cq;
  input [144:0] fp_cpx_data_ca;
  input [155:0] inq_sram_din_unbuf;
  output [63:0] inq_in1_add_buf1;
  output [63:0] inq_in1_mul_buf1;
  output [63:0] inq_in1_div_buf1;
  output [63:0] inq_in2_add_buf1;
  output [63:0] inq_in2_mul_buf1;
  output [63:0] inq_in2_div_buf1;
  output [4:0] inq_id_add_buf1;
  output [4:0] inq_id_mul_buf1;
  output [4:0] inq_id_div_buf1;
  output [7:0] inq_op_add_buf1;
  output [7:0] inq_op_div_buf1;
  output [7:0] inq_op_mul_buf1;
  output [1:0] inq_rnd_mode_add_buf1;
  output [1:0] inq_rnd_mode_div_buf1;
  output [1:0] inq_rnd_mode_mul_buf1;
  output [123:0] pcx_fpio_data_px2_buf1;
  output [7:0] fp_cpx_req_cq_buf1;
  output [144:0] fp_cpx_data_ca_buf1;
  output [155:0] inq_sram_din_buf1;
  input inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0,
         inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l,
         ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain,
         global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l,
         fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf,
         pcx_fpio_data_rdy_px2;
  output inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1,
         inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1,
         inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1,
         inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1,
         inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1,
         inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1,
         inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1,
         inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1,
         inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1,
         inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1,
         inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1,
         inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1,
         inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1,
         inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1,
         inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1,
         ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1,
         ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1,
         ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1,
         cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2,
         se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4,
         se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2,
         arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3,
         arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2,
         fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1,
         fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so,
         pcx_fpio_data_rdy_px2_buf1;
  wire   se_add_buf1, se_mul64_buf1, so_buf1, se_buf1_unused,
         se_add_buf2_unused, arst_l_buf1;
  wire   [3:0] inq_id_add_buf1_unused;
  wire   [2:0] inq_id_mul_buf1_unused;
  wire   [4:0] inq_id_div_buf1_unused;
  wire   [1:0] ctu_tst_buf1_lo_unused;
  wire   [1:0] cluster_cken_buf1_unused;
  wire   [1:0] se_mul64_buf2_unused;
  wire   [2:0] arst_l_buf1_unused;
  wire   [1:0] fdiv_clken_l_buf1_unused;
  wire   [2:0] so_cluster_header_buf1_unused;
  wire   [2:0] si_buf1_unused;
  wire   [2:0] pcx_fpio_data_px2_buf1_unused;
  wire   [5:0] fp_cpx_buf1_9_unused;

  fpu_bufrpt_grp32 i_inq_in1_add_buf1_hi ( .in(inq_in1[63:32]), .out(
        inq_in1_add_buf1[63:32]) );
  fpu_bufrpt_grp32 i_inq_in1_add_buf1_lo ( .in(inq_in1[31:0]), .out(
        inq_in1_add_buf1[31:0]) );
  fpu_bufrpt_grp32 i_inq_in1_mul_buf1_hi ( .in(inq_in1[63:32]), .out(
        inq_in1_mul_buf1[63:32]) );
  fpu_bufrpt_grp32 i_inq_in1_mul_buf1_lo ( .in(inq_in1[31:0]), .out(
        inq_in1_mul_buf1[31:0]) );
  fpu_bufrpt_grp64 i_inq_in1_div_buf1 ( .in(inq_in1), .out(inq_in1_div_buf1)
         );
  fpu_bufrpt_grp32 i_inq_in2_add_buf1_hi ( .in(inq_in2[63:32]), .out(
        inq_in2_add_buf1[63:32]) );
  fpu_bufrpt_grp32 i_inq_in2_add_buf1_lo ( .in(inq_in2[31:0]), .out(
        inq_in2_add_buf1[31:0]) );
  fpu_bufrpt_grp32 i_inq_in2_mul_buf1_hi ( .in(inq_in2[63:32]), .out(
        inq_in2_mul_buf1[63:32]) );
  fpu_bufrpt_grp32 i_inq_in2_mul_buf1_lo ( .in(inq_in2[31:0]), .out(
        inq_in2_mul_buf1[31:0]) );
  fpu_bufrpt_grp64 i_inq_in2_div_buf1 ( .in(inq_in2), .out(inq_in2_div_buf1)
         );
  fpu_bufrpt_grp32 i_inq_id_add_buf1 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 
        se_out_buf2, arst_l_out_buf3, fpu_grst_l_in_buf2, inq_id, inq_op, 
        inq_rnd_mode, inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, 
        inq_in2_50_0_neq_0, inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs}), .out({inq_id_add_buf1_unused, 
        se_in_buf3, arst_l_add_buf4, fpu_grst_l_add_buf3, inq_id_add_buf1, 
        inq_op_add_buf1, inq_rnd_mode_add_buf1, inq_in1_50_0_neq_0_add_buf1, 
        inq_in1_53_0_neq_0_add_buf1, inq_in1_53_32_neq_0_add_buf1, 
        inq_in1_exp_eq_0_add_buf1, inq_in1_exp_neq_ffs_add_buf1, 
        inq_in2_50_0_neq_0_add_buf1, inq_in2_53_0_neq_0_add_buf1, 
        inq_in2_53_32_neq_0_add_buf1, inq_in2_exp_eq_0_add_buf1, 
        inq_in2_exp_neq_ffs_add_buf1}) );
  fpu_bufrpt_grp32 i_inq_id_mul_buf1 ( .in({1'b0, 1'b0, 1'b0, se_in_buf3, 
        arst_l_mul_buf2, fpu_grst_l_mul_buf1, fmul_clken_l, inq_id, inq_op, 
        inq_rnd_mode, inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, 
        inq_in1_53_32_neq_0, inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, 
        inq_in2_50_0_neq_0, inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs}), .out({inq_id_mul_buf1_unused, 
        se_mul_buf4, arst_l_out_buf3, fpu_grst_l_in_buf2, fmul_clken_l_buf1, 
        inq_id_mul_buf1, inq_op_mul_buf1, inq_rnd_mode_mul_buf1, 
        inq_in1_50_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_mul_buf1, 
        inq_in1_53_32_neq_0_mul_buf1, inq_in1_exp_eq_0_mul_buf1, 
        inq_in1_exp_neq_ffs_mul_buf1, inq_in2_50_0_neq_0_mul_buf1, 
        inq_in2_53_0_neq_0_mul_buf1, inq_in2_53_32_neq_0_mul_buf1, 
        inq_in2_exp_eq_0_mul_buf1, inq_in2_exp_neq_ffs_mul_buf1}) );
  fpu_bufrpt_grp32 i_inq_id_div_buf1 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        se_mul_buf4, arst_l_mul_buf2, inq_id, inq_op, inq_rnd_mode, 
        inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0, 
        inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, 
        inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs}), .out({inq_id_div_buf1_unused, se_div_buf5, 
        arst_l_in_buf3, inq_id_div_buf1, inq_op_div_buf1, 
        inq_rnd_mode_div_buf1, inq_in1_50_0_neq_0_div_buf1, 
        inq_in1_53_0_neq_0_div_buf1, inq_in1_53_32_neq_0_div_buf1, 
        inq_in1_exp_eq_0_div_buf1, inq_in1_exp_neq_ffs_div_buf1, 
        inq_in2_50_0_neq_0_div_buf1, inq_in2_53_0_neq_0_div_buf1, 
        inq_in2_53_32_neq_0_div_buf1, inq_in2_exp_eq_0_div_buf1, 
        inq_in2_exp_neq_ffs_div_buf1}) );
  fpu_bufrpt_grp4 i_ctu_tst_buf1_hi ( .in({ctu_tst_short_chain, 
        ctu_tst_macrotest, ctu_tst_scan_disable, ctu_tst_pre_grst_l}), .out({
        ctu_tst_short_chain_buf1, ctu_tst_macrotest_buf1, 
        ctu_tst_scan_disable_buf1, ctu_tst_pre_grst_l_buf1}) );
  fpu_bufrpt_grp4 i_ctu_tst_buf1_lo ( .in({ctu_tst_scanmode, 
        global_shift_enable, 1'b0, 1'b0}), .out({ctu_tst_scanmode_buf1, 
        global_shift_enable_buf1, ctu_tst_buf1_lo_unused}) );
  fpu_bufrpt_grp4 i_cluster_cken_buf1 ( .in({cluster_cken, grst_l, 1'b0, 1'b0}), .out({cluster_cken_buf1, grst_l_buf1, cluster_cken_buf1_unused}) );
  fpu_bufrpt_grp4 i_se_buf1 ( .in({se, se, so_unbuf, 1'b0}), .out({se_add_buf1, 
        se_mul64_buf1, so_buf1, se_buf1_unused}) );
  fpu_bufrpt_grp4 i_se_add_buf2 ( .in({se_add_buf1, se_add_buf1, se_add_buf1, 
        1'b0}), .out({se_add_exp_buf2, se_add_frac_buf2, se_out_buf2, 
        se_add_buf2_unused}) );
  fpu_bufrpt_grp4 i_se_mul64_buf2 ( .in({se_mul64_buf1, se_mul64_buf1, 1'b0, 
        1'b0}), .out({se_mul64_buf2, se_cluster_header_buf2, 
        se_mul64_buf2_unused}) );
  fpu_bufrpt_grp4 i_arst_l_buf1 ( .in({arst_l, 1'b0, 1'b0, 1'b0}), .out({
        arst_l_buf1, arst_l_buf1_unused}) );
  fpu_bufrpt_grp4 i_arst_l_buf2 ( .in({arst_l_buf1, arst_l_buf1, arst_l_buf1, 
        fpu_grst_l}), .out({arst_l_mul_buf2, arst_l_cluster_header_buf2, 
        arst_l_div_buf2, fpu_grst_l_mul_buf1}) );
  fpu_bufrpt_grp4 i_fdiv_clken_l_buf1 ( .in({fdiv_clken_l, fdiv_clken_l, 1'b0, 
        1'b0}), .out({fdiv_clken_l_div_exp_buf1, fdiv_clken_l_div_frac_buf1, 
        fdiv_clken_l_buf1_unused}) );
  fpu_bufrpt_grp4 i_so_cluster_header_buf1 ( .in({scan_manual_6, 1'b0, 1'b0, 
        1'b0}), .out({scan_manual_6_buf1, so_cluster_header_buf1_unused}) );
  fpu_bufrpt_grp4 i_si_buf1 ( .in({si, 1'b0, 1'b0, 1'b0}), .out({si_buf1, 
        si_buf1_unused}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_0 ( .in({pcx_fpio_data_px2[108], 
        pcx_fpio_data_px2[109], pcx_fpio_data_px2[110], pcx_fpio_data_px2[111], 
        pcx_fpio_data_px2[112], pcx_fpio_data_px2[113], pcx_fpio_data_px2[114], 
        pcx_fpio_data_px2[115], pcx_fpio_data_px2[116], pcx_fpio_data_px2[117], 
        pcx_fpio_data_px2[118], pcx_fpio_data_px2[119], pcx_fpio_data_px2[120], 
        pcx_fpio_data_px2[121], pcx_fpio_data_px2[122], pcx_fpio_data_px2[123]}), .out({pcx_fpio_data_px2_buf1[108], pcx_fpio_data_px2_buf1[109], 
        pcx_fpio_data_px2_buf1[110], pcx_fpio_data_px2_buf1[111], 
        pcx_fpio_data_px2_buf1[112], pcx_fpio_data_px2_buf1[113], 
        pcx_fpio_data_px2_buf1[114], pcx_fpio_data_px2_buf1[115], 
        pcx_fpio_data_px2_buf1[116], pcx_fpio_data_px2_buf1[117], 
        pcx_fpio_data_px2_buf1[118], pcx_fpio_data_px2_buf1[119], 
        pcx_fpio_data_px2_buf1[120], pcx_fpio_data_px2_buf1[121], 
        pcx_fpio_data_px2_buf1[122], pcx_fpio_data_px2_buf1[123]}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_1 ( .in({pcx_fpio_data_px2[92], 
        pcx_fpio_data_px2[93], pcx_fpio_data_px2[94], pcx_fpio_data_px2[95], 
        pcx_fpio_data_px2[96], pcx_fpio_data_px2[97], pcx_fpio_data_px2[98], 
        pcx_fpio_data_px2[99], pcx_fpio_data_px2[100], pcx_fpio_data_px2[101], 
        pcx_fpio_data_px2[102], pcx_fpio_data_px2[103], pcx_fpio_data_px2[104], 
        pcx_fpio_data_px2[105], pcx_fpio_data_px2[106], pcx_fpio_data_px2[107]}), .out({pcx_fpio_data_px2_buf1[92], pcx_fpio_data_px2_buf1[93], 
        pcx_fpio_data_px2_buf1[94], pcx_fpio_data_px2_buf1[95], 
        pcx_fpio_data_px2_buf1[96], pcx_fpio_data_px2_buf1[97], 
        pcx_fpio_data_px2_buf1[98], pcx_fpio_data_px2_buf1[99], 
        pcx_fpio_data_px2_buf1[100], pcx_fpio_data_px2_buf1[101], 
        pcx_fpio_data_px2_buf1[102], pcx_fpio_data_px2_buf1[103], 
        pcx_fpio_data_px2_buf1[104], pcx_fpio_data_px2_buf1[105], 
        pcx_fpio_data_px2_buf1[106], pcx_fpio_data_px2_buf1[107]}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_2 ( .in({pcx_fpio_data_px2[76], 
        pcx_fpio_data_px2[77], pcx_fpio_data_px2[78], pcx_fpio_data_px2[79], 
        pcx_fpio_data_px2[80], pcx_fpio_data_px2[81], pcx_fpio_data_px2[82], 
        pcx_fpio_data_px2[83], pcx_fpio_data_px2[84], pcx_fpio_data_px2[85], 
        pcx_fpio_data_px2[86], pcx_fpio_data_px2[87], pcx_fpio_data_px2[88], 
        pcx_fpio_data_px2[89], pcx_fpio_data_px2[90], pcx_fpio_data_px2[91]}), 
        .out({pcx_fpio_data_px2_buf1[76], pcx_fpio_data_px2_buf1[77], 
        pcx_fpio_data_px2_buf1[78], pcx_fpio_data_px2_buf1[79], 
        pcx_fpio_data_px2_buf1[80], pcx_fpio_data_px2_buf1[81], 
        pcx_fpio_data_px2_buf1[82], pcx_fpio_data_px2_buf1[83], 
        pcx_fpio_data_px2_buf1[84], pcx_fpio_data_px2_buf1[85], 
        pcx_fpio_data_px2_buf1[86], pcx_fpio_data_px2_buf1[87], 
        pcx_fpio_data_px2_buf1[88], pcx_fpio_data_px2_buf1[89], 
        pcx_fpio_data_px2_buf1[90], pcx_fpio_data_px2_buf1[91]}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_3 ( .in({pcx_fpio_data_px2[3:0], 
        pcx_fpio_data_px2[64], pcx_fpio_data_px2[65], pcx_fpio_data_px2[66], 
        pcx_fpio_data_px2[67], pcx_fpio_data_px2[68], pcx_fpio_data_px2[69], 
        pcx_fpio_data_px2[70], pcx_fpio_data_px2[71], pcx_fpio_data_px2[72], 
        pcx_fpio_data_px2[73], pcx_fpio_data_px2[74], pcx_fpio_data_px2[75]}), 
        .out({pcx_fpio_data_px2_buf1[3:0], pcx_fpio_data_px2_buf1[64], 
        pcx_fpio_data_px2_buf1[65], pcx_fpio_data_px2_buf1[66], 
        pcx_fpio_data_px2_buf1[67], pcx_fpio_data_px2_buf1[68], 
        pcx_fpio_data_px2_buf1[69], pcx_fpio_data_px2_buf1[70], 
        pcx_fpio_data_px2_buf1[71], pcx_fpio_data_px2_buf1[72], 
        pcx_fpio_data_px2_buf1[73], pcx_fpio_data_px2_buf1[74], 
        pcx_fpio_data_px2_buf1[75]}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_4 ( .in(pcx_fpio_data_px2[19:4]), 
        .out(pcx_fpio_data_px2_buf1[19:4]) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_5 ( .in(pcx_fpio_data_px2[35:20]), 
        .out(pcx_fpio_data_px2_buf1[35:20]) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_6 ( .in({pcx_fpio_data_rdy_px2, 
        pcx_fpio_data_px2[50:36]}), .out({pcx_fpio_data_rdy_px2_buf1, 
        pcx_fpio_data_px2_buf1[50:36]}) );
  fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_7 ( .in({1'b0, 1'b0, 1'b0, 
        pcx_fpio_data_px2[63:51]}), .out({pcx_fpio_data_px2_buf1_unused, 
        pcx_fpio_data_px2_buf1[63:51]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_0 ( .in({fp_cpx_data_ca[142], 
        fp_cpx_data_ca[140], fp_cpx_data_ca[138], fp_cpx_data_ca[136], 
        fp_cpx_data_ca[134], fp_cpx_data_ca[132], fp_cpx_data_ca[130], 
        fp_cpx_data_ca[128], fp_cpx_req_cq[6], fp_cpx_req_cq[7], 
        fp_cpx_req_cq[3:2], fp_cpx_req_cq[5], fp_cpx_req_cq[1:0], 
        fp_cpx_req_cq[4]}), .out({fp_cpx_data_ca_buf1[142], 
        fp_cpx_data_ca_buf1[140], fp_cpx_data_ca_buf1[138], 
        fp_cpx_data_ca_buf1[136], fp_cpx_data_ca_buf1[134], 
        fp_cpx_data_ca_buf1[132], fp_cpx_data_ca_buf1[130], 
        fp_cpx_data_ca_buf1[128], fp_cpx_req_cq_buf1[6], fp_cpx_req_cq_buf1[7], 
        fp_cpx_req_cq_buf1[3:2], fp_cpx_req_cq_buf1[5], 
        fp_cpx_req_cq_buf1[1:0], fp_cpx_req_cq_buf1[4]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_1 ( .in({fp_cpx_data_ca[34], 
        fp_cpx_data_ca[36], fp_cpx_data_ca[38], fp_cpx_data_ca[40], 
        fp_cpx_data_ca[42], fp_cpx_data_ca[44], fp_cpx_data_ca[46], 
        fp_cpx_data_ca[48], fp_cpx_data_ca[50], fp_cpx_data_ca[52], 
        fp_cpx_data_ca[54], fp_cpx_data_ca[56], fp_cpx_data_ca[58], 
        fp_cpx_data_ca[60], fp_cpx_data_ca[62], fp_cpx_data_ca[144]}), .out({
        fp_cpx_data_ca_buf1[34], fp_cpx_data_ca_buf1[36], 
        fp_cpx_data_ca_buf1[38], fp_cpx_data_ca_buf1[40], 
        fp_cpx_data_ca_buf1[42], fp_cpx_data_ca_buf1[44], 
        fp_cpx_data_ca_buf1[46], fp_cpx_data_ca_buf1[48], 
        fp_cpx_data_ca_buf1[50], fp_cpx_data_ca_buf1[52], 
        fp_cpx_data_ca_buf1[54], fp_cpx_data_ca_buf1[56], 
        fp_cpx_data_ca_buf1[58], fp_cpx_data_ca_buf1[60], 
        fp_cpx_data_ca_buf1[62], fp_cpx_data_ca_buf1[144]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_2 ( .in({fp_cpx_data_ca[2], 
        fp_cpx_data_ca[4], fp_cpx_data_ca[6], fp_cpx_data_ca[8], 
        fp_cpx_data_ca[10], fp_cpx_data_ca[12], fp_cpx_data_ca[14], 
        fp_cpx_data_ca[16], fp_cpx_data_ca[18], fp_cpx_data_ca[20], 
        fp_cpx_data_ca[22], fp_cpx_data_ca[24], fp_cpx_data_ca[26], 
        fp_cpx_data_ca[28], fp_cpx_data_ca[30], fp_cpx_data_ca[32]}), .out({
        fp_cpx_data_ca_buf1[2], fp_cpx_data_ca_buf1[4], fp_cpx_data_ca_buf1[6], 
        fp_cpx_data_ca_buf1[8], fp_cpx_data_ca_buf1[10], 
        fp_cpx_data_ca_buf1[12], fp_cpx_data_ca_buf1[14], 
        fp_cpx_data_ca_buf1[16], fp_cpx_data_ca_buf1[18], 
        fp_cpx_data_ca_buf1[20], fp_cpx_data_ca_buf1[22], 
        fp_cpx_data_ca_buf1[24], fp_cpx_data_ca_buf1[26], 
        fp_cpx_data_ca_buf1[28], fp_cpx_data_ca_buf1[30], 
        fp_cpx_data_ca_buf1[32]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_3 ( .in({fp_cpx_data_ca[31], 
        fp_cpx_data_ca[27], fp_cpx_data_ca[23], fp_cpx_data_ca[25], 
        fp_cpx_data_ca[21], fp_cpx_data_ca[17], fp_cpx_data_ca[19], 
        fp_cpx_data_ca[15], fp_cpx_data_ca[11], fp_cpx_data_ca[13], 
        fp_cpx_data_ca[9], fp_cpx_data_ca[5], fp_cpx_data_ca[7], 
        fp_cpx_data_ca[3], fp_cpx_data_ca[0], fp_cpx_data_ca[1]}), .out({
        fp_cpx_data_ca_buf1[31], fp_cpx_data_ca_buf1[27], 
        fp_cpx_data_ca_buf1[23], fp_cpx_data_ca_buf1[25], 
        fp_cpx_data_ca_buf1[21], fp_cpx_data_ca_buf1[17], 
        fp_cpx_data_ca_buf1[19], fp_cpx_data_ca_buf1[15], 
        fp_cpx_data_ca_buf1[11], fp_cpx_data_ca_buf1[13], 
        fp_cpx_data_ca_buf1[9], fp_cpx_data_ca_buf1[5], fp_cpx_data_ca_buf1[7], 
        fp_cpx_data_ca_buf1[3], fp_cpx_data_ca_buf1[0], fp_cpx_data_ca_buf1[1]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_4 ( .in({fp_cpx_data_ca[59], 
        fp_cpx_data_ca[61], fp_cpx_data_ca[57], fp_cpx_data_ca[53], 
        fp_cpx_data_ca[55], fp_cpx_data_ca[51], fp_cpx_data_ca[47], 
        fp_cpx_data_ca[49], fp_cpx_data_ca[45], fp_cpx_data_ca[41], 
        fp_cpx_data_ca[43], fp_cpx_data_ca[39], fp_cpx_data_ca[35], 
        fp_cpx_data_ca[37], fp_cpx_data_ca[33], fp_cpx_data_ca[29]}), .out({
        fp_cpx_data_ca_buf1[59], fp_cpx_data_ca_buf1[61], 
        fp_cpx_data_ca_buf1[57], fp_cpx_data_ca_buf1[53], 
        fp_cpx_data_ca_buf1[55], fp_cpx_data_ca_buf1[51], 
        fp_cpx_data_ca_buf1[47], fp_cpx_data_ca_buf1[49], 
        fp_cpx_data_ca_buf1[45], fp_cpx_data_ca_buf1[41], 
        fp_cpx_data_ca_buf1[43], fp_cpx_data_ca_buf1[39], 
        fp_cpx_data_ca_buf1[35], fp_cpx_data_ca_buf1[37], 
        fp_cpx_data_ca_buf1[33], fp_cpx_data_ca_buf1[29]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_5 ( .in({fp_cpx_data_ca[113], 
        fp_cpx_data_ca[117], fp_cpx_data_ca[121], fp_cpx_data_ca[119], 
        fp_cpx_data_ca[123], fp_cpx_data_ca[127], fp_cpx_data_ca[125], 
        fp_cpx_data_ca[129], fp_cpx_data_ca[133], fp_cpx_data_ca[131], 
        fp_cpx_data_ca[135], fp_cpx_data_ca[139], fp_cpx_data_ca[137], 
        fp_cpx_data_ca[141], fp_cpx_data_ca[143], fp_cpx_data_ca[63]}), .out({
        fp_cpx_data_ca_buf1[113], fp_cpx_data_ca_buf1[117], 
        fp_cpx_data_ca_buf1[121], fp_cpx_data_ca_buf1[119], 
        fp_cpx_data_ca_buf1[123], fp_cpx_data_ca_buf1[127], 
        fp_cpx_data_ca_buf1[125], fp_cpx_data_ca_buf1[129], 
        fp_cpx_data_ca_buf1[133], fp_cpx_data_ca_buf1[131], 
        fp_cpx_data_ca_buf1[135], fp_cpx_data_ca_buf1[139], 
        fp_cpx_data_ca_buf1[137], fp_cpx_data_ca_buf1[141], 
        fp_cpx_data_ca_buf1[143], fp_cpx_data_ca_buf1[63]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_6 ( .in({fp_cpx_data_ca[85], 
        fp_cpx_data_ca[83], fp_cpx_data_ca[87], fp_cpx_data_ca[91], 
        fp_cpx_data_ca[89], fp_cpx_data_ca[93], fp_cpx_data_ca[97], 
        fp_cpx_data_ca[95], fp_cpx_data_ca[99], fp_cpx_data_ca[103], 
        fp_cpx_data_ca[101], fp_cpx_data_ca[105], fp_cpx_data_ca[109], 
        fp_cpx_data_ca[107], fp_cpx_data_ca[111], fp_cpx_data_ca[115]}), .out(
        {fp_cpx_data_ca_buf1[85], fp_cpx_data_ca_buf1[83], 
        fp_cpx_data_ca_buf1[87], fp_cpx_data_ca_buf1[91], 
        fp_cpx_data_ca_buf1[89], fp_cpx_data_ca_buf1[93], 
        fp_cpx_data_ca_buf1[97], fp_cpx_data_ca_buf1[95], 
        fp_cpx_data_ca_buf1[99], fp_cpx_data_ca_buf1[103], 
        fp_cpx_data_ca_buf1[101], fp_cpx_data_ca_buf1[105], 
        fp_cpx_data_ca_buf1[109], fp_cpx_data_ca_buf1[107], 
        fp_cpx_data_ca_buf1[111], fp_cpx_data_ca_buf1[115]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_7 ( .in({fp_cpx_data_ca[114], 
        fp_cpx_data_ca[116], fp_cpx_data_ca[118], fp_cpx_data_ca[120], 
        fp_cpx_data_ca[122], fp_cpx_data_ca[124], fp_cpx_data_ca[126], 
        fp_cpx_data_ca[65], fp_cpx_data_ca[67], fp_cpx_data_ca[69], 
        fp_cpx_data_ca[73], fp_cpx_data_ca[71], fp_cpx_data_ca[75], 
        fp_cpx_data_ca[79], fp_cpx_data_ca[77], fp_cpx_data_ca[81]}), .out({
        fp_cpx_data_ca_buf1[114], fp_cpx_data_ca_buf1[116], 
        fp_cpx_data_ca_buf1[118], fp_cpx_data_ca_buf1[120], 
        fp_cpx_data_ca_buf1[122], fp_cpx_data_ca_buf1[124], 
        fp_cpx_data_ca_buf1[126], fp_cpx_data_ca_buf1[65], 
        fp_cpx_data_ca_buf1[67], fp_cpx_data_ca_buf1[69], 
        fp_cpx_data_ca_buf1[73], fp_cpx_data_ca_buf1[71], 
        fp_cpx_data_ca_buf1[75], fp_cpx_data_ca_buf1[79], 
        fp_cpx_data_ca_buf1[77], fp_cpx_data_ca_buf1[81]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_8 ( .in({fp_cpx_data_ca[82], 
        fp_cpx_data_ca[84], fp_cpx_data_ca[86], fp_cpx_data_ca[88], 
        fp_cpx_data_ca[90], fp_cpx_data_ca[92], fp_cpx_data_ca[94], 
        fp_cpx_data_ca[96], fp_cpx_data_ca[98], fp_cpx_data_ca[100], 
        fp_cpx_data_ca[102], fp_cpx_data_ca[104], fp_cpx_data_ca[106], 
        fp_cpx_data_ca[108], fp_cpx_data_ca[110], fp_cpx_data_ca[112]}), .out(
        {fp_cpx_data_ca_buf1[82], fp_cpx_data_ca_buf1[84], 
        fp_cpx_data_ca_buf1[86], fp_cpx_data_ca_buf1[88], 
        fp_cpx_data_ca_buf1[90], fp_cpx_data_ca_buf1[92], 
        fp_cpx_data_ca_buf1[94], fp_cpx_data_ca_buf1[96], 
        fp_cpx_data_ca_buf1[98], fp_cpx_data_ca_buf1[100], 
        fp_cpx_data_ca_buf1[102], fp_cpx_data_ca_buf1[104], 
        fp_cpx_data_ca_buf1[106], fp_cpx_data_ca_buf1[108], 
        fp_cpx_data_ca_buf1[110], fp_cpx_data_ca_buf1[112]}) );
  fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_9 ( .in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, so_buf1, fp_cpx_data_ca[64], fp_cpx_data_ca[66], 
        fp_cpx_data_ca[68], fp_cpx_data_ca[70], fp_cpx_data_ca[72], 
        fp_cpx_data_ca[74], fp_cpx_data_ca[76], fp_cpx_data_ca[78], 
        fp_cpx_data_ca[80]}), .out({fp_cpx_buf1_9_unused, so, 
        fp_cpx_data_ca_buf1[64], fp_cpx_data_ca_buf1[66], 
        fp_cpx_data_ca_buf1[68], fp_cpx_data_ca_buf1[70], 
        fp_cpx_data_ca_buf1[72], fp_cpx_data_ca_buf1[74], 
        fp_cpx_data_ca_buf1[76], fp_cpx_data_ca_buf1[78], 
        fp_cpx_data_ca_buf1[80]}) );
  fpu_rptr_inq i_inq_sram_din_buf1 ( .in(inq_sram_din_unbuf), .out(
        inq_sram_din_buf1) );
endmodule


module fpu ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, arst_l, grst_l, gclk, 
        cluster_cken, fp_cpx_req_cq, fp_cpx_data_ca, ctu_tst_pre_grst_l, 
        global_shift_enable, ctu_tst_scan_disable, ctu_tst_scanmode, 
        ctu_tst_macrotest, ctu_tst_short_chain, si, so );
  input [123:0] pcx_fpio_data_px2;
  output [7:0] fp_cpx_req_cq;
  output [144:0] fp_cpx_data_ca;
  input pcx_fpio_data_rdy_px2, arst_l, grst_l, gclk, cluster_cken,
         ctu_tst_pre_grst_l, global_shift_enable, ctu_tst_scan_disable,
         ctu_tst_scanmode, ctu_tst_macrotest, ctu_tst_short_chain, si;
  output so;
  wire   pcx_fpio_data_rdy_px2_buf1, a1stg_step, m1stg_step, d1stg_step,
         add_pipe_active, mul_pipe_active, div_pipe_active, sehold,
         arst_l_in_buf3, fpu_grst_l_in_buf2, rclk, fadd_clken_l, fmul_clken_l,
         fdiv_clken_l, inq_add, inq_mul, inq_div, inq_in1_exp_neq_ffs,
         inq_in1_exp_eq_0, inq_in1_53_0_neq_0, inq_in1_50_0_neq_0,
         inq_in1_53_32_neq_0, inq_in2_exp_neq_ffs, inq_in2_exp_eq_0,
         inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0,
         inq_read_en, inq_we, se_in_buf3, manual_scan_0, scan_manual_1, se,
         si_buf1, scan_inq_sram_w, rst_tri_en, inq_in1_50_0_neq_0_add_buf1,
         inq_in1_53_32_neq_0_add_buf1, inq_in1_exp_eq_0_add_buf1,
         inq_in1_exp_neq_ffs_add_buf1, inq_in2_50_0_neq_0_add_buf1,
         inq_in2_53_32_neq_0_add_buf1, inq_in2_exp_eq_0_add_buf1,
         inq_in2_exp_neq_ffs_add_buf1, add_dest_rdy, arst_l_add_buf4,
         fpu_grst_l_add_buf3, a6stg_fadd_in, a6stg_fcmpop, a6stg_dbl_dst,
         a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, add_sign_out,
         se_add_exp_buf2, se_add_frac_buf2, scan_manual_2,
         inq_in1_50_0_neq_0_mul_buf1, inq_in1_53_32_neq_0_mul_buf1,
         inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_neq_ffs_mul_buf1,
         inq_in2_50_0_neq_0_mul_buf1, inq_in2_53_32_neq_0_mul_buf1,
         inq_in2_exp_eq_0_mul_buf1, inq_in2_exp_neq_ffs_mul_buf1, mul_dest_rdy,
         fmul_clken_l_buf1, arst_l_mul_buf2, fpu_grst_l_mul_buf1,
         m6stg_fmul_in, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out,
         se_mul_buf4, se_mul64_buf2, scan_manual_3,
         inq_in1_53_0_neq_0_div_buf1, inq_in1_50_0_neq_0_div_buf1,
         inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_div_buf1,
         inq_in1_exp_neq_ffs_div_buf1, inq_in2_53_0_neq_0_div_buf1,
         inq_in2_50_0_neq_0_div_buf1, inq_in2_53_32_neq_0_div_buf1,
         inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_div_buf1, div_dest_rdy,
         fdiv_clken_l_div_frac_buf1, fdiv_clken_l_div_exp_buf1,
         arst_l_div_buf2, fpu_grst_l, d8stg_fdiv_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, se_div_buf5, scan_manual_4, arst_l_out_buf3,
         se_out_buf2, scan_manual_5, ctu_tst_pre_grst_l_buf1,
         global_shift_enable_buf1, ctu_tst_scan_disable_buf1,
         ctu_tst_scanmode_buf1, ctu_tst_macrotest_buf1,
         ctu_tst_short_chain_buf1, scan_manual_6_buf1, so_unbuf,
         cluster_cken_buf1, arst_l_cluster_header_buf2, grst_l_buf1,
         se_cluster_header_buf2, scan_manual_6, inq_in1_53_0_neq_0_add_buf1,
         inq_in1_53_0_neq_0_mul_buf1, inq_in2_53_0_neq_0_add_buf1,
         inq_in2_53_0_neq_0_mul_buf1;
  wire   [123:0] pcx_fpio_data_px2_buf1;
  wire   [154:0] inq_dout;
  wire   [4:0] inq_id;
  wire   [1:0] inq_rnd_mode;
  wire   [1:0] inq_fcc;
  wire   [7:0] inq_op;
  wire   [63:0] inq_in1;
  wire   [63:0] inq_in2;
  wire   [4:0] fp_id_in;
  wire   [1:0] fp_rnd_mode_in;
  wire   [1:0] fp_fcc_in;
  wire   [7:0] fp_op_in;
  wire   [68:0] fp_src1_in;
  wire   [68:0] fp_src2_in;
  wire   [3:0] inq_rdaddr;
  wire   [3:0] inq_wraddr;
  wire   [4:0] inq_dout_unused;
  wire   [155:0] inq_sram_din_buf1;
  wire   [7:0] inq_op_add_buf1;
  wire   [1:0] inq_rnd_mode_add_buf1;
  wire   [4:0] inq_id_add_buf1;
  wire   [63:0] inq_in1_add_buf1;
  wire   [63:0] inq_in2_add_buf1;
  wire   [9:0] add_id_out_in;
  wire   [4:0] add_exc_out;
  wire   [10:0] add_exp_out;
  wire   [63:0] add_frac_out;
  wire   [1:0] add_cc_out;
  wire   [1:0] add_fcc_out;
  wire   [7:0] inq_op_mul_buf1;
  wire   [1:0] inq_rnd_mode_mul_buf1;
  wire   [4:0] inq_id_mul_buf1;
  wire   [63:0] inq_in1_mul_buf1;
  wire   [63:0] inq_in2_mul_buf1;
  wire   [9:0] m6stg_id_in;
  wire   [4:0] mul_exc_out;
  wire   [10:0] mul_exp_out;
  wire   [51:0] mul_frac_out;
  wire   [7:0] inq_op_div_buf1;
  wire   [1:0] inq_rnd_mode_div_buf1;
  wire   [4:0] inq_id_div_buf1;
  wire   [63:0] inq_in1_div_buf1;
  wire   [63:0] inq_in2_div_buf1;
  wire   [9:0] div_id_out_in;
  wire   [4:0] div_exc_out;
  wire   [10:0] div_exp_out;
  wire   [51:0] div_frac_out;
  wire   [7:0] fp_cpx_req_cq_unbuf;
  wire   [144:0] fp_cpx_data_ca_unbuf;

  fpu_in fpu_in ( .pcx_fpio_data_rdy_px2(pcx_fpio_data_rdy_px2_buf1), 
        .pcx_fpio_data_px2(pcx_fpio_data_px2_buf1), .a1stg_step(a1stg_step), 
        .m1stg_step(m1stg_step), .d1stg_step(d1stg_step), .add_pipe_active(
        add_pipe_active), .mul_pipe_active(mul_pipe_active), .div_pipe_active(
        div_pipe_active), .inq_dout(inq_dout), .sehold(sehold), .arst_l(
        arst_l_in_buf3), .grst_l(fpu_grst_l_in_buf2), .rclk(rclk), 
        .fadd_clken_l(fadd_clken_l), .fmul_clken_l(fmul_clken_l), 
        .fdiv_clken_l(fdiv_clken_l), .inq_add(inq_add), .inq_mul(inq_mul), 
        .inq_div(inq_div), .inq_id(inq_id), .inq_rnd_mode(inq_rnd_mode), 
        .inq_fcc(inq_fcc), .inq_op(inq_op), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in1_exp_eq_0(inq_in1_exp_eq_0), 
        .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1(inq_in1), .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), 
        .inq_in2_exp_eq_0(inq_in2_exp_eq_0), .inq_in2_53_0_neq_0(
        inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0), .inq_in2(inq_in2), 
        .fp_id_in(fp_id_in), .fp_rnd_mode_in(fp_rnd_mode_in), .fp_fcc_in(
        fp_fcc_in), .fp_op_in(fp_op_in), .fp_src1_in(fp_src1_in), .fp_src2_in(
        fp_src2_in), .inq_rdaddr(inq_rdaddr), .inq_wraddr(inq_wraddr), 
        .inq_read_en(inq_read_en), .inq_we(inq_we), .se(se_in_buf3), .si(
        manual_scan_0), .so(scan_manual_1) );
  bw_r_rf16x160 bw_r_rf16x160 ( .dout({inq_dout, inq_dout_unused}), .so_w(
        manual_scan_0), .so_r(scan_inq_sram_w), .din({inq_sram_din_buf1, 1'b0, 
        1'b0, 1'b0, 1'b0}), .rd_adr(inq_rdaddr), .wr_adr(inq_wraddr), 
        .read_en(inq_read_en), .wr_en(inq_we), .rst_tri_en(rst_tri_en), 
        .word_wen({1'b1, 1'b1, 1'b1, 1'b1}), .byte_wen({1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .rd_clk(rclk), .wr_clk(rclk), .se(se), 
        .si_r(si_buf1), .si_w(scan_inq_sram_w), .reset_l(arst_l_in_buf3), 
        .sehold(sehold) );
  fpu_add fpu_add ( .inq_op(inq_op_add_buf1), .inq_rnd_mode(
        inq_rnd_mode_add_buf1), .inq_id(inq_id_add_buf1), .inq_fcc(inq_fcc), 
        .inq_in1(inq_in1_add_buf1), .inq_in1_50_0_neq_0(
        inq_in1_50_0_neq_0_add_buf1), .inq_in1_53_32_neq_0(
        inq_in1_53_32_neq_0_add_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_add_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_add_buf1), .inq_in2(inq_in2_add_buf1), 
        .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0_add_buf1), 
        .inq_in2_53_32_neq_0(inq_in2_53_32_neq_0_add_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_add_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_add_buf1), .inq_add(inq_add), .add_dest_rdy(
        add_dest_rdy), .fadd_clken_l(fadd_clken_l), .arst_l(arst_l_add_buf4), 
        .grst_l(fpu_grst_l_add_buf3), .rclk(rclk), .add_pipe_active(
        add_pipe_active), .a1stg_step(a1stg_step), .a6stg_fadd_in(
        a6stg_fadd_in), .add_id_out_in(add_id_out_in), .a6stg_fcmpop(
        a6stg_fcmpop), .add_exc_out(add_exc_out), .a6stg_dbl_dst(a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), .a6stg_long_dst(a6stg_long_dst), 
        .a6stg_int_dst(a6stg_int_dst), .add_sign_out(add_sign_out), 
        .add_exp_out(add_exp_out), .add_frac_out(add_frac_out), .add_cc_out(
        add_cc_out), .add_fcc_out(add_fcc_out), .se_add_exp(se_add_exp_buf2), 
        .se_add_frac(se_add_frac_buf2), .si(scan_manual_1), .so(scan_manual_2)
         );
  fpu_mul fpu_mul ( .inq_op(inq_op_mul_buf1), .inq_rnd_mode(
        inq_rnd_mode_mul_buf1), .inq_id(inq_id_mul_buf1), .inq_in1(
        inq_in1_mul_buf1), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0_mul_buf1), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0_mul_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_mul_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_mul_buf1), .inq_in2(inq_in2_mul_buf1), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0_mul_buf1), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0_mul_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_mul_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_mul_buf1), .inq_mul(inq_mul), .mul_dest_rdy(
        mul_dest_rdy), .mul_dest_rdya(mul_dest_rdy), .fmul_clken_l(
        fmul_clken_l), .fmul_clken_l_buf1(fmul_clken_l_buf1), .arst_l(
        arst_l_mul_buf2), .grst_l(fpu_grst_l_mul_buf1), .rclk(rclk), 
        .mul_pipe_active(mul_pipe_active), .m1stg_step(m1stg_step), 
        .m6stg_fmul_in(m6stg_fmul_in), .m6stg_id_in(m6stg_id_in), 
        .mul_exc_out(mul_exc_out), .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), 
        .m6stg_fmuls(m6stg_fmuls), .mul_sign_out(mul_sign_out), .mul_exp_out(
        mul_exp_out), .mul_frac_out(mul_frac_out), .se_mul(se_mul_buf4), 
        .se_mul64(se_mul64_buf2), .si(scan_manual_2), .so(scan_manual_3) );
  fpu_div fpu_div ( .inq_op(inq_op_div_buf1), .inq_rnd_mode(
        inq_rnd_mode_div_buf1), .inq_id(inq_id_div_buf1), .inq_in1(
        inq_in1_div_buf1), .inq_in1_53_0_neq_0(inq_in1_53_0_neq_0_div_buf1), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0_div_buf1), 
        .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0_div_buf1), .inq_in1_exp_eq_0(
        inq_in1_exp_eq_0_div_buf1), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs_div_buf1), .inq_in2(inq_in2_div_buf1), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0_div_buf1), .inq_in2_50_0_neq_0(
        inq_in2_50_0_neq_0_div_buf1), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0_div_buf1), .inq_in2_exp_eq_0(
        inq_in2_exp_eq_0_div_buf1), .inq_in2_exp_neq_ffs(
        inq_in2_exp_neq_ffs_div_buf1), .inq_div(inq_div), .div_dest_rdy(
        div_dest_rdy), .fdiv_clken_l(fdiv_clken_l_div_frac_buf1), 
        .fdiv_clken_l_div_exp_buf1(fdiv_clken_l_div_exp_buf1), .arst_l(
        arst_l_div_buf2), .grst_l(fpu_grst_l), .rclk(rclk), .div_pipe_active(
        div_pipe_active), .d1stg_step(d1stg_step), .d8stg_fdiv_in(
        d8stg_fdiv_in), .div_id_out_in(div_id_out_in), .div_exc_out(
        div_exc_out), .d8stg_fdivd(d8stg_fdivd), .d8stg_fdivs(d8stg_fdivs), 
        .div_sign_out(div_sign_out), .div_exp_outa(div_exp_out), 
        .div_frac_outa(div_frac_out), .se(se_div_buf5), .si(scan_manual_3), 
        .so(scan_manual_4) );
  fpu_out fpu_out ( .d8stg_fdiv_in(d8stg_fdiv_in), .m6stg_fmul_in(
        m6stg_fmul_in), .a6stg_fadd_in(a6stg_fadd_in), .div_id_out_in(
        div_id_out_in), .m6stg_id_in(m6stg_id_in), .add_id_out_in(
        add_id_out_in), .div_exc_out(div_exc_out), .d8stg_fdivd(d8stg_fdivd), 
        .d8stg_fdivs(d8stg_fdivs), .div_sign_out(div_sign_out), .div_exp_out(
        div_exp_out), .div_frac_out(div_frac_out), .mul_exc_out(mul_exc_out), 
        .m6stg_fmul_dbl_dst(m6stg_fmul_dbl_dst), .m6stg_fmuls(m6stg_fmuls), 
        .mul_sign_out(mul_sign_out), .mul_exp_out(mul_exp_out), .mul_frac_out(
        mul_frac_out), .add_exc_out(add_exc_out), .a6stg_fcmpop(a6stg_fcmpop), 
        .add_cc_out(add_cc_out), .add_fcc_out(add_fcc_out), .a6stg_dbl_dst(
        a6stg_dbl_dst), .a6stg_sng_dst(a6stg_sng_dst), .a6stg_long_dst(
        a6stg_long_dst), .a6stg_int_dst(a6stg_int_dst), .add_sign_out(
        add_sign_out), .add_exp_out(add_exp_out), .add_frac_out(add_frac_out), 
        .arst_l(arst_l_out_buf3), .grst_l(fpu_grst_l_add_buf3), .rclk(rclk), 
        .fp_cpx_req_cq(fp_cpx_req_cq_unbuf), .add_dest_rdy(add_dest_rdy), 
        .mul_dest_rdy(mul_dest_rdy), .div_dest_rdy(div_dest_rdy), 
        .fp_cpx_data_ca(fp_cpx_data_ca_unbuf), .se(se_out_buf2), .si(
        scan_manual_4), .so(scan_manual_5) );
  test_stub_scan test_stub_scan ( .mem_write_disable(rst_tri_en), .sehold(
        sehold), .se(se), .so_0(so_unbuf), .ctu_tst_pre_grst_l(
        ctu_tst_pre_grst_l_buf1), .arst_l(arst_l_add_buf4), 
        .global_shift_enable(global_shift_enable_buf1), .ctu_tst_scan_disable(
        ctu_tst_scan_disable_buf1), .ctu_tst_scanmode(ctu_tst_scanmode_buf1), 
        .ctu_tst_macrotest(ctu_tst_macrotest_buf1), .ctu_tst_short_chain(
        ctu_tst_short_chain_buf1), .long_chain_so_0(scan_manual_6_buf1), 
        .short_chain_so_0(manual_scan_0), .long_chain_so_1(1'b0), 
        .short_chain_so_1(1'b0), .long_chain_so_2(1'b0), .short_chain_so_2(
        1'b0) );
  bw_clk_cl_fpu_cmp cluster_header ( .so(scan_manual_6), .cluster_grst_l(
        fpu_grst_l), .rclk(rclk), .si(scan_manual_5), .se(
        se_cluster_header_buf2), .adbginit_l(1'b1), .gdbginit_l(1'b1), 
        .arst_l(arst_l_cluster_header_buf2), .grst_l(grst_l_buf1), 
        .cluster_cken(cluster_cken_buf1), .gclk(gclk) );
  fpu_rptr_groups fpu_rptr_groups ( .inq_in1(inq_in1), .inq_in2(inq_in2), 
        .inq_id(inq_id), .inq_op(inq_op), .inq_rnd_mode(inq_rnd_mode), 
        .inq_in1_50_0_neq_0(inq_in1_50_0_neq_0), .inq_in1_53_0_neq_0(
        inq_in1_53_0_neq_0), .inq_in1_53_32_neq_0(inq_in1_53_32_neq_0), 
        .inq_in1_exp_eq_0(inq_in1_exp_eq_0), .inq_in1_exp_neq_ffs(
        inq_in1_exp_neq_ffs), .inq_in2_50_0_neq_0(inq_in2_50_0_neq_0), 
        .inq_in2_53_0_neq_0(inq_in2_53_0_neq_0), .inq_in2_53_32_neq_0(
        inq_in2_53_32_neq_0), .inq_in2_exp_eq_0(inq_in2_exp_eq_0), 
        .inq_in2_exp_neq_ffs(inq_in2_exp_neq_ffs), .ctu_tst_macrotest(
        ctu_tst_macrotest), .ctu_tst_pre_grst_l(ctu_tst_pre_grst_l), 
        .ctu_tst_scan_disable(ctu_tst_scan_disable), .ctu_tst_scanmode(
        ctu_tst_scanmode), .ctu_tst_short_chain(ctu_tst_short_chain), 
        .global_shift_enable(global_shift_enable), .grst_l(grst_l), 
        .cluster_cken(cluster_cken), .se(se), .arst_l(arst_l), .fpu_grst_l(
        fpu_grst_l), .fmul_clken_l(fmul_clken_l), .fdiv_clken_l(fdiv_clken_l), 
        .scan_manual_6(scan_manual_6), .si(si), .so_unbuf(so_unbuf), 
        .pcx_fpio_data_px2(pcx_fpio_data_px2), .pcx_fpio_data_rdy_px2(
        pcx_fpio_data_rdy_px2), .fp_cpx_req_cq(fp_cpx_req_cq_unbuf), 
        .fp_cpx_data_ca(fp_cpx_data_ca_unbuf), .inq_sram_din_unbuf({fp_id_in, 
        fp_rnd_mode_in, fp_fcc_in, fp_op_in, fp_src1_in, fp_src2_in, 1'b0}), 
        .inq_in1_add_buf1(inq_in1_add_buf1), .inq_in1_mul_buf1(
        inq_in1_mul_buf1), .inq_in1_div_buf1(inq_in1_div_buf1), 
        .inq_in2_add_buf1(inq_in2_add_buf1), .inq_in2_mul_buf1(
        inq_in2_mul_buf1), .inq_in2_div_buf1(inq_in2_div_buf1), 
        .inq_id_add_buf1(inq_id_add_buf1), .inq_id_mul_buf1(inq_id_mul_buf1), 
        .inq_id_div_buf1(inq_id_div_buf1), .inq_op_add_buf1(inq_op_add_buf1), 
        .inq_op_div_buf1(inq_op_div_buf1), .inq_op_mul_buf1(inq_op_mul_buf1), 
        .inq_rnd_mode_add_buf1(inq_rnd_mode_add_buf1), .inq_rnd_mode_div_buf1(
        inq_rnd_mode_div_buf1), .inq_rnd_mode_mul_buf1(inq_rnd_mode_mul_buf1), 
        .inq_in1_50_0_neq_0_add_buf1(inq_in1_50_0_neq_0_add_buf1), 
        .inq_in1_50_0_neq_0_mul_buf1(inq_in1_50_0_neq_0_mul_buf1), 
        .inq_in1_50_0_neq_0_div_buf1(inq_in1_50_0_neq_0_div_buf1), 
        .inq_in1_53_0_neq_0_add_buf1(inq_in1_53_0_neq_0_add_buf1), 
        .inq_in1_53_0_neq_0_mul_buf1(inq_in1_53_0_neq_0_mul_buf1), 
        .inq_in1_53_0_neq_0_div_buf1(inq_in1_53_0_neq_0_div_buf1), 
        .inq_in1_53_32_neq_0_add_buf1(inq_in1_53_32_neq_0_add_buf1), 
        .inq_in1_53_32_neq_0_mul_buf1(inq_in1_53_32_neq_0_mul_buf1), 
        .inq_in1_53_32_neq_0_div_buf1(inq_in1_53_32_neq_0_div_buf1), 
        .inq_in1_exp_eq_0_add_buf1(inq_in1_exp_eq_0_add_buf1), 
        .inq_in1_exp_eq_0_mul_buf1(inq_in1_exp_eq_0_mul_buf1), 
        .inq_in1_exp_eq_0_div_buf1(inq_in1_exp_eq_0_div_buf1), 
        .inq_in1_exp_neq_ffs_add_buf1(inq_in1_exp_neq_ffs_add_buf1), 
        .inq_in1_exp_neq_ffs_mul_buf1(inq_in1_exp_neq_ffs_mul_buf1), 
        .inq_in1_exp_neq_ffs_div_buf1(inq_in1_exp_neq_ffs_div_buf1), 
        .inq_in2_50_0_neq_0_add_buf1(inq_in2_50_0_neq_0_add_buf1), 
        .inq_in2_50_0_neq_0_mul_buf1(inq_in2_50_0_neq_0_mul_buf1), 
        .inq_in2_50_0_neq_0_div_buf1(inq_in2_50_0_neq_0_div_buf1), 
        .inq_in2_53_0_neq_0_add_buf1(inq_in2_53_0_neq_0_add_buf1), 
        .inq_in2_53_0_neq_0_mul_buf1(inq_in2_53_0_neq_0_mul_buf1), 
        .inq_in2_53_0_neq_0_div_buf1(inq_in2_53_0_neq_0_div_buf1), 
        .inq_in2_53_32_neq_0_add_buf1(inq_in2_53_32_neq_0_add_buf1), 
        .inq_in2_53_32_neq_0_mul_buf1(inq_in2_53_32_neq_0_mul_buf1), 
        .inq_in2_53_32_neq_0_div_buf1(inq_in2_53_32_neq_0_div_buf1), 
        .inq_in2_exp_eq_0_add_buf1(inq_in2_exp_eq_0_add_buf1), 
        .inq_in2_exp_eq_0_mul_buf1(inq_in2_exp_eq_0_mul_buf1), 
        .inq_in2_exp_eq_0_div_buf1(inq_in2_exp_eq_0_div_buf1), 
        .inq_in2_exp_neq_ffs_add_buf1(inq_in2_exp_neq_ffs_add_buf1), 
        .inq_in2_exp_neq_ffs_mul_buf1(inq_in2_exp_neq_ffs_mul_buf1), 
        .inq_in2_exp_neq_ffs_div_buf1(inq_in2_exp_neq_ffs_div_buf1), 
        .ctu_tst_macrotest_buf1(ctu_tst_macrotest_buf1), 
        .ctu_tst_pre_grst_l_buf1(ctu_tst_pre_grst_l_buf1), 
        .ctu_tst_scan_disable_buf1(ctu_tst_scan_disable_buf1), 
        .ctu_tst_scanmode_buf1(ctu_tst_scanmode_buf1), 
        .ctu_tst_short_chain_buf1(ctu_tst_short_chain_buf1), 
        .global_shift_enable_buf1(global_shift_enable_buf1), .grst_l_buf1(
        grst_l_buf1), .cluster_cken_buf1(cluster_cken_buf1), .se_add_exp_buf2(
        se_add_exp_buf2), .se_add_frac_buf2(se_add_frac_buf2), .se_out_buf2(
        se_out_buf2), .se_mul64_buf2(se_mul64_buf2), .se_cluster_header_buf2(
        se_cluster_header_buf2), .se_in_buf3(se_in_buf3), .se_mul_buf4(
        se_mul_buf4), .se_div_buf5(se_div_buf5), .arst_l_div_buf2(
        arst_l_div_buf2), .arst_l_mul_buf2(arst_l_mul_buf2), 
        .arst_l_cluster_header_buf2(arst_l_cluster_header_buf2), 
        .arst_l_in_buf3(arst_l_in_buf3), .arst_l_out_buf3(arst_l_out_buf3), 
        .arst_l_add_buf4(arst_l_add_buf4), .fpu_grst_l_mul_buf1(
        fpu_grst_l_mul_buf1), .fpu_grst_l_in_buf2(fpu_grst_l_in_buf2), 
        .fpu_grst_l_add_buf3(fpu_grst_l_add_buf3), .fmul_clken_l_buf1(
        fmul_clken_l_buf1), .fdiv_clken_l_div_exp_buf1(
        fdiv_clken_l_div_exp_buf1), .fdiv_clken_l_div_frac_buf1(
        fdiv_clken_l_div_frac_buf1), .scan_manual_6_buf1(scan_manual_6_buf1), 
        .si_buf1(si_buf1), .so(so), .pcx_fpio_data_px2_buf1(
        pcx_fpio_data_px2_buf1), .pcx_fpio_data_rdy_px2_buf1(
        pcx_fpio_data_rdy_px2_buf1), .fp_cpx_req_cq_buf1(fp_cpx_req_cq), 
        .fp_cpx_data_ca_buf1(fp_cpx_data_ca), .inq_sram_din_buf1(
        inq_sram_din_buf1) );
endmodule

